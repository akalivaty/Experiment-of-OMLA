//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n570, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT66), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(new_n467), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G137), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n468), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n478));
  OR2_X1    g053(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n473), .A2(new_n469), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n474), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n469), .B2(G112), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n468), .B(new_n492), .C1(new_n491), .C2(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n473), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n469), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n495), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n505), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n512), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n512), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n523), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(new_n511), .A2(new_n518), .A3(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(new_n517), .ZN(new_n532));
  INV_X1    g107(.A(new_n513), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n532), .A2(G51), .A3(G543), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n509), .A2(new_n510), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n508), .A2(G543), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n535), .A2(G63), .A3(G651), .A4(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n538), .B1(new_n534), .B2(new_n537), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n531), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT71), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n531), .B(new_n543), .C1(new_n539), .C2(new_n540), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(G168));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n519), .A2(new_n546), .B1(new_n521), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n512), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(G171));
  AND2_X1   g126(.A1(new_n511), .A2(new_n518), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G81), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n518), .A2(G43), .A3(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n505), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT69), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n557));
  OAI211_X1 g132(.A(G56), .B(new_n536), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT72), .B1(new_n560), .B2(G651), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  AOI211_X1 g137(.A(new_n562), .B(new_n512), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n553), .B(new_n555), .C1(new_n561), .C2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G860), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT73), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  XOR2_X1   g144(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n570));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G188));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n521), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n518), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(KEYINPUT75), .B(G65), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n511), .A2(new_n580), .B1(G78), .B2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G91), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n581), .A2(new_n512), .B1(new_n519), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n574), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n579), .A2(new_n583), .A3(new_n574), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(G299));
  INV_X1    g162(.A(G171), .ZN(G301));
  INV_X1    g163(.A(G168), .ZN(G286));
  INV_X1    g164(.A(new_n521), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G49), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n552), .A2(G87), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  INV_X1    g169(.A(G48), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n521), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n512), .ZN(new_n598));
  AOI211_X1 g173(.A(new_n596), .B(new_n598), .C1(G86), .C2(new_n552), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G305));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n519), .A2(new_n601), .B1(new_n521), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n512), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n603), .A2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n519), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n511), .A2(new_n518), .A3(KEYINPUT10), .A4(G92), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n590), .A2(G54), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(new_n512), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT77), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n607), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n607), .B1(new_n617), .B2(G868), .ZN(G321));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(G299), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(G168), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n620), .B2(G168), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n617), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(new_n564), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(G868), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n468), .A2(new_n480), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n483), .A2(G123), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n474), .A2(G135), .ZN(new_n636));
  NOR2_X1   g211(.A1(G99), .A2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(new_n469), .B2(G111), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n634), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT78), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2430), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT79), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n654), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n656), .B2(KEYINPUT80), .ZN(new_n657));
  AOI211_X1 g232(.A(new_n655), .B(new_n657), .C1(KEYINPUT80), .C2(new_n656), .ZN(G401));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XOR2_X1   g234(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT82), .Z(new_n665));
  INV_X1    g240(.A(new_n663), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n659), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n666), .B(new_n667), .C1(new_n661), .C2(new_n662), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n666), .A2(new_n662), .A3(new_n659), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n665), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n675), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n679), .A2(KEYINPUT20), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n683), .A2(new_n675), .A3(new_n678), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n682), .B(new_n684), .C1(KEYINPUT20), .C2(new_n679), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1986), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1981), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1991), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(G229));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G22), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G1971), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(G6), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n599), .B2(new_n692), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n692), .A2(G23), .ZN(new_n700));
  INV_X1    g275(.A(G288), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n692), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT86), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n695), .A2(new_n699), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT34), .Z(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G24), .ZN(new_n708));
  XOR2_X1   g283(.A(G290), .B(KEYINPUT85), .Z(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G16), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G1986), .Z(new_n711));
  AOI22_X1  g286(.A1(G119), .A2(new_n483), .B1(new_n474), .B2(G131), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n464), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n715), .B1(new_n714), .B2(new_n713), .C1(G107), .C2(new_n469), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G25), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT83), .B1(new_n719), .B2(G29), .ZN(new_n720));
  OR3_X1    g295(.A1(new_n719), .A2(KEYINPUT83), .A3(G29), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n722), .B(new_n723), .Z(new_n724));
  NAND3_X1  g299(.A1(new_n707), .A2(new_n711), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT36), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n617), .A2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT87), .B1(G4), .B2(G16), .ZN(new_n728));
  OR3_X1    g303(.A1(KEYINPUT87), .A2(G4), .A3(G16), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT88), .B(G1348), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n730), .B(new_n731), .Z(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G33), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT90), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n736), .A2(G2105), .B1(G139), .B2(new_n474), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n480), .A2(G103), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G2072), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G5), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G171), .B2(G16), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n741), .A2(new_n742), .B1(G1961), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT28), .ZN(new_n747));
  INV_X1    g322(.A(G26), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G29), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n483), .A2(G128), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n474), .A2(G140), .ZN(new_n752));
  NOR2_X1   g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n749), .B1(new_n756), .B2(new_n747), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G2067), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(G2067), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n743), .A2(new_n746), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n761), .A2(new_n733), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G160), .B2(new_n733), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(G2084), .ZN(new_n765));
  NOR2_X1   g340(.A1(G29), .A2(G32), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n483), .A2(G129), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT91), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT26), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n480), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n766), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT27), .B(G1996), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n733), .A2(G27), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G164), .B2(new_n733), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G2078), .Z(new_n779));
  INV_X1    g354(.A(G28), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(KEYINPUT30), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT30), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n781), .A2(new_n782), .A3(new_n733), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n639), .B2(new_n733), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n764), .B2(G2084), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n760), .A2(new_n765), .A3(new_n776), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT31), .B(G11), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT92), .ZN(new_n789));
  INV_X1    g364(.A(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT89), .B1(new_n790), .B2(G16), .ZN(new_n791));
  OR3_X1    g366(.A1(new_n790), .A2(KEYINPUT89), .A3(G16), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n628), .C2(new_n692), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1341), .Z(new_n794));
  INV_X1    g369(.A(G35), .ZN(new_n795));
  OAI21_X1  g370(.A(KEYINPUT93), .B1(new_n795), .B2(G29), .ZN(new_n796));
  OR3_X1    g371(.A1(new_n795), .A2(KEYINPUT93), .A3(G29), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n796), .B(new_n797), .C1(G162), .C2(new_n733), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT29), .B(G2090), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G1961), .ZN(new_n801));
  INV_X1    g376(.A(new_n745), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n787), .A2(new_n789), .A3(new_n794), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n692), .A2(G21), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G168), .B2(new_n692), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(G1966), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(G1966), .ZN(new_n808));
  NAND2_X1  g383(.A1(G299), .A2(G16), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n692), .A2(KEYINPUT23), .A3(G20), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT23), .ZN(new_n811));
  INV_X1    g386(.A(G20), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G16), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n809), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1956), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n804), .A2(new_n807), .A3(new_n808), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n726), .A2(new_n732), .A3(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  NAND2_X1  g393(.A1(new_n617), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n511), .A2(G67), .ZN(new_n821));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n512), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n511), .A2(new_n518), .A3(G93), .ZN(new_n824));
  AND2_X1   g399(.A1(KEYINPUT94), .A2(G55), .ZN(new_n825));
  NOR2_X1   g400(.A1(KEYINPUT94), .A2(G55), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n532), .A2(G543), .A3(new_n533), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT95), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT95), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n824), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n823), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n564), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n823), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n824), .A2(new_n831), .A3(new_n828), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n831), .B1(new_n824), .B2(new_n828), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n559), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n511), .B2(G56), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n562), .B1(new_n840), .B2(new_n512), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n560), .A2(KEYINPUT72), .A3(G651), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n554), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n838), .A2(new_n553), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n834), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n820), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  OR3_X1    g423(.A1(new_n847), .A2(KEYINPUT96), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT96), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n848), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n565), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n833), .A2(new_n565), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT97), .ZN(G145));
  XNOR2_X1  g431(.A(new_n772), .B(new_n755), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n495), .B2(new_n503), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n492), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n494), .B1(new_n860), .B2(new_n473), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n469), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n498), .A2(G2105), .B1(new_n501), .B2(new_n500), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(KEYINPUT98), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n857), .B(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n737), .A2(KEYINPUT99), .A3(new_n739), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G160), .B(G162), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n483), .A2(G130), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n474), .A2(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(new_n469), .B2(G118), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n632), .B(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n868), .A2(new_n869), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n870), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT99), .B1(new_n737), .B2(new_n739), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n717), .B(new_n639), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n876), .B1(new_n877), .B2(new_n870), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n878), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n878), .B2(new_n883), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g463(.A1(new_n833), .A2(new_n620), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n616), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n585), .B2(new_n586), .ZN(new_n892));
  INV_X1    g467(.A(new_n583), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n893), .A2(KEYINPUT76), .A3(new_n577), .A4(new_n578), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n584), .A3(new_n616), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n897), .A2(KEYINPUT100), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(KEYINPUT100), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n626), .B(new_n846), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n902), .A2(KEYINPUT101), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(new_n892), .B2(new_n895), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n894), .A2(new_n584), .A3(new_n616), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n616), .B1(new_n894), .B2(new_n584), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n901), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n902), .A2(KEYINPUT101), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT102), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n701), .B(G303), .ZN(new_n913));
  INV_X1    g488(.A(G290), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G303), .B(G288), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(G290), .ZN(new_n917));
  OAI21_X1  g492(.A(G305), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(G290), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n599), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT42), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n912), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n911), .A2(KEYINPUT102), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n890), .B1(new_n926), .B2(G868), .ZN(G295));
  AOI21_X1  g502(.A(new_n890), .B1(new_n926), .B2(G868), .ZN(G331));
  AND3_X1   g503(.A1(new_n542), .A2(new_n544), .A3(G301), .ZN(new_n929));
  AOI21_X1  g504(.A(G301), .B1(new_n542), .B2(new_n544), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n929), .A2(new_n845), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n534), .A2(new_n537), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT70), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n543), .B1(new_n935), .B2(new_n531), .ZN(new_n936));
  INV_X1    g511(.A(new_n544), .ZN(new_n937));
  OAI21_X1  g512(.A(G171), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n542), .A2(new_n544), .A3(G301), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n938), .A2(new_n939), .B1(new_n844), .B2(new_n834), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n931), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(new_n898), .B2(new_n899), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n907), .B1(new_n905), .B2(new_n906), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n845), .B1(new_n929), .B2(new_n930), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n938), .A2(new_n844), .A3(new_n834), .A4(new_n939), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n892), .A2(KEYINPUT41), .A3(new_n895), .ZN(new_n946));
  AND4_X1   g521(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n921), .B(new_n918), .C1(new_n942), .C2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n896), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT104), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n922), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n948), .A2(new_n954), .A3(new_n885), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n948), .A2(new_n954), .A3(KEYINPUT107), .A4(new_n885), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(KEYINPUT43), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n918), .A2(new_n960), .A3(new_n921), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n950), .A2(new_n961), .A3(new_n953), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n918), .A2(new_n960), .A3(new_n921), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n897), .B1(new_n931), .B2(new_n940), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n952), .B1(new_n964), .B2(new_n951), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n908), .A2(new_n904), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT104), .B1(new_n941), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n962), .A2(new_n968), .A3(new_n885), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n970), .ZN(new_n974));
  INV_X1    g549(.A(new_n970), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n948), .A2(new_n954), .A3(new_n885), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g554(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n974), .C2(new_n976), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n972), .B(KEYINPUT108), .C1(new_n979), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(G397));
  AOI21_X1  g560(.A(G1384), .B1(new_n859), .B2(new_n864), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n987));
  AND4_X1   g562(.A1(G40), .A2(new_n477), .A3(new_n479), .A4(new_n481), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1996), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(new_n773), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(KEYINPUT109), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n991), .A2(KEYINPUT109), .ZN(new_n993));
  INV_X1    g568(.A(new_n989), .ZN(new_n994));
  INV_X1    g569(.A(G2067), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n755), .B(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n772), .B2(G1996), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n992), .B(new_n993), .C1(new_n994), .C2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n717), .B(new_n723), .Z(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n989), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(G290), .B(G1986), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n994), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n495), .B2(new_n503), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n862), .B2(new_n863), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n988), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT121), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1005), .A2(new_n988), .A3(new_n1008), .A4(KEYINPUT121), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n731), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n988), .A2(new_n995), .A3(new_n1006), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n579), .A2(new_n583), .A3(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1017), .A2(KEYINPUT120), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(KEYINPUT120), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n579), .A2(KEYINPUT119), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n577), .B2(new_n578), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1020), .A2(new_n583), .A3(new_n1022), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1018), .A2(new_n1019), .B1(new_n1023), .B2(KEYINPUT57), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1004), .A2(KEYINPUT110), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT56), .B(G2072), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1025), .A2(new_n1030), .A3(new_n988), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1956), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1009), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1024), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1015), .A2(new_n891), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1024), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT60), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1015), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1013), .A2(KEYINPUT60), .A3(new_n1014), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n891), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT61), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1035), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1024), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1039), .A2(KEYINPUT61), .A3(new_n1035), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1013), .A2(KEYINPUT60), .A3(new_n616), .A4(new_n1014), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1043), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1025), .A2(new_n1030), .A3(new_n990), .A4(new_n988), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT58), .B(G1341), .Z(new_n1052));
  INV_X1    g627(.A(new_n988), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1053), .B2(new_n1004), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n564), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT59), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1036), .B(new_n1039), .C1(new_n1050), .C2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(G171), .B(KEYINPUT54), .Z(new_n1058));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G2078), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n865), .A2(new_n1003), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1053), .B1(new_n1061), .B2(new_n1026), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1060), .B1(new_n1062), .B2(KEYINPUT124), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT124), .B(new_n988), .C1(new_n986), .C2(KEYINPUT45), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1025), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1058), .B1(new_n1066), .B2(KEYINPUT125), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1011), .A2(new_n801), .A3(new_n1012), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1025), .A2(new_n1030), .A3(new_n988), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1059), .B1(new_n1069), .B2(G2078), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n1074));
  INV_X1    g649(.A(G8), .ZN(new_n1075));
  OR3_X1    g650(.A1(G168), .A2(KEYINPUT122), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT122), .B1(G168), .B2(new_n1075), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1004), .A2(new_n1026), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n988), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1966), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT117), .B(G2084), .Z(new_n1085));
  NAND4_X1  g660(.A1(new_n1005), .A2(new_n988), .A3(new_n1008), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1075), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1074), .B1(new_n1079), .B2(new_n1088), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1078), .A2(new_n1087), .A3(KEYINPUT51), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1078), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n1078), .B2(new_n1092), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1089), .A2(new_n1090), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1060), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1070), .B(new_n1068), .C1(new_n1082), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1058), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1073), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1057), .A2(new_n1099), .ZN(new_n1100));
  OR3_X1    g675(.A1(new_n1088), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1095), .A2(KEYINPUT62), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n1103));
  OAI221_X1 g678(.A(new_n1103), .B1(new_n1093), .B2(new_n1094), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1102), .A2(new_n1104), .A3(G171), .A4(new_n1097), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1009), .A2(G2090), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT111), .B(G1971), .Z(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1069), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n1075), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G303), .A2(G8), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1111), .B(KEYINPUT55), .Z(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT114), .B(G86), .Z(new_n1115));
  OAI22_X1  g690(.A1(new_n519), .A2(new_n1115), .B1(new_n521), .B2(new_n595), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1116), .B(KEYINPUT115), .Z(new_n1117));
  OAI21_X1  g692(.A(G1981), .B1(new_n1117), .B2(new_n598), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT113), .B(G1981), .Z(new_n1119));
  NAND2_X1  g694(.A1(new_n599), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT49), .ZN(new_n1122));
  OAI21_X1  g697(.A(G8), .B1(new_n1053), .B2(new_n1004), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G1976), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G288), .A2(new_n1126), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1123), .A2(KEYINPUT112), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n1129));
  NAND2_X1  g704(.A1(G288), .A2(new_n1126), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1123), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1128), .B(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1133), .A2(KEYINPUT116), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(KEYINPUT116), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1106), .A2(new_n1114), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1125), .A2(new_n1126), .A3(new_n701), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1123), .B1(new_n1139), .B2(new_n1120), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT118), .B1(new_n1133), .B2(new_n1113), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1114), .A2(new_n1142), .A3(new_n1125), .A4(new_n1132), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1088), .A2(G286), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .A4(new_n1135), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1140), .B1(new_n1145), .B2(KEYINPUT63), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1135), .B2(new_n1133), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1002), .B1(new_n1138), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n755), .A2(G2067), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n717), .A2(new_n723), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n998), .B2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n989), .A2(G1986), .A3(G290), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT127), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT48), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1151), .A2(new_n989), .B1(new_n1000), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n994), .A2(KEYINPUT46), .A3(new_n990), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT46), .B1(new_n994), .B2(new_n990), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n989), .B1(new_n773), .B2(new_n996), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT126), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT47), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1155), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1148), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g738(.A1(G229), .A2(new_n462), .ZN(new_n1165));
  NOR2_X1   g739(.A1(G401), .A2(G227), .ZN(new_n1166));
  NAND4_X1  g740(.A1(new_n887), .A2(new_n977), .A3(new_n1165), .A4(new_n1166), .ZN(G225));
  INV_X1    g741(.A(G225), .ZN(G308));
endmodule


