//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G227), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G953), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G143), .B(G146), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  OAI211_X1 g008(.A(KEYINPUT76), .B(KEYINPUT1), .C1(new_n194), .C2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT76), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n193), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n194), .A2(G146), .ZN(new_n204));
  AND4_X1   g018(.A1(new_n203), .A2(new_n198), .A3(new_n204), .A4(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT77), .B(new_n193), .C1(new_n196), .C2(new_n199), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G104), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n214), .A2(KEYINPUT74), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n216), .A2(new_n211), .A3(new_n215), .A4(new_n213), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n210), .A2(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n213), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n217), .A2(new_n220), .B1(G101), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n208), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(G101), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n218), .A2(new_n219), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n218), .A2(new_n219), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n192), .B1(G128), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(new_n205), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT11), .A3(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(G137), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G131), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT64), .B(G131), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n242), .A2(new_n236), .A3(new_n238), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT12), .B1(new_n233), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n246));
  INV_X1    g060(.A(new_n244), .ZN(new_n247));
  AOI211_X1 g061(.A(new_n246), .B(new_n247), .C1(new_n224), .C2(new_n232), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n198), .A2(new_n204), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT0), .B(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n192), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n217), .A2(new_n220), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n216), .A2(new_n211), .A3(new_n213), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G101), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n253), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n255), .A3(G101), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n256), .A2(KEYINPUT75), .A3(new_n255), .A4(G101), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT10), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n231), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n258), .A2(new_n263), .B1(new_n223), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n224), .A2(new_n264), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n244), .B(KEYINPUT78), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n191), .B1(new_n249), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n257), .B1(new_n226), .B2(new_n227), .ZN(new_n272));
  INV_X1    g086(.A(new_n253), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n263), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n265), .A2(new_n223), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT10), .B1(new_n208), .B2(new_n223), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT79), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT79), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n266), .A2(new_n267), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n280), .A3(new_n244), .ZN(new_n281));
  INV_X1    g095(.A(new_n191), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n269), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n271), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n187), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n282), .B1(new_n281), .B2(new_n269), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n269), .A2(new_n282), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n249), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n187), .B(new_n285), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT80), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n291), .A2(new_n292), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n287), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n296));
  INV_X1    g110(.A(G221), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n299), .B2(new_n285), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n295), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n266), .A2(new_n267), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n247), .B1(new_n303), .B2(KEYINPUT79), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n270), .B1(new_n304), .B2(new_n280), .ZN(new_n305));
  OAI22_X1  g119(.A1(new_n305), .A2(new_n282), .B1(new_n249), .B2(new_n289), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n306), .A2(KEYINPUT80), .A3(new_n187), .A4(new_n285), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n291), .A2(new_n292), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n286), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT81), .B1(new_n309), .B2(new_n300), .ZN(new_n310));
  XNOR2_X1  g124(.A(G125), .B(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G125), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n314), .A2(KEYINPUT16), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(G146), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(G146), .B1(new_n312), .B2(new_n315), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  INV_X1    g134(.A(G953), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G214), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n194), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n320), .A2(new_n321), .A3(G143), .A4(G214), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT64), .B(G131), .Z(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(KEYINPUT17), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT86), .B1(new_n325), .B2(new_n326), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n323), .A2(new_n330), .A3(new_n242), .A4(new_n324), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n319), .B(new_n327), .C1(new_n332), .C2(KEYINPUT17), .ZN(new_n333));
  INV_X1    g147(.A(new_n325), .ZN(new_n334));
  NAND3_X1  g148(.A1(KEYINPUT85), .A2(KEYINPUT18), .A3(G131), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n314), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G146), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n311), .A2(new_n197), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n334), .A2(new_n335), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n336), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n333), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G113), .B(G122), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n212), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n333), .A2(new_n347), .A3(new_n344), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT89), .B(G475), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT19), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n339), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n311), .A2(KEYINPUT19), .ZN(new_n356));
  AOI21_X1  g170(.A(G146), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT87), .B1(new_n317), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n355), .A2(new_n356), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n316), .B(new_n359), .C1(new_n360), .C2(G146), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n361), .A3(new_n332), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT88), .A3(new_n344), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n348), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT88), .B1(new_n362), .B2(new_n344), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n350), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G475), .A2(G902), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT20), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n372), .A3(new_n367), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n353), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n321), .A2(G952), .ZN(new_n375));
  INV_X1    g189(.A(G234), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(new_n320), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT21), .ZN(new_n379));
  OAI21_X1  g193(.A(G953), .B1(new_n379), .B2(G898), .ZN(new_n380));
  INV_X1    g194(.A(G898), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(KEYINPUT21), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n285), .B1(G234), .B2(G237), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G478), .ZN(new_n387));
  INV_X1    g201(.A(G217), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n298), .A2(new_n388), .A3(G953), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G116), .B(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT90), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n210), .ZN(new_n393));
  INV_X1    g207(.A(G116), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT14), .A3(G122), .ZN(new_n395));
  INV_X1    g209(.A(new_n391), .ZN(new_n396));
  OAI211_X1 g210(.A(G107), .B(new_n395), .C1(new_n396), .C2(KEYINPUT14), .ZN(new_n397));
  XNOR2_X1  g211(.A(G128), .B(G143), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n235), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n393), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT90), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n391), .B(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G107), .ZN(new_n404));
  INV_X1    g218(.A(G128), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G143), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT13), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n235), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n408), .A2(new_n398), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n398), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n404), .A2(new_n393), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n390), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n404), .A2(new_n393), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n409), .A2(new_n410), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n400), .B(new_n389), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  AOI211_X1 g230(.A(KEYINPUT15), .B(new_n387), .C1(new_n416), .C2(new_n285), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n285), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n387), .A2(KEYINPUT15), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n374), .A2(new_n386), .A3(new_n421), .ZN(new_n422));
  XOR2_X1   g236(.A(KEYINPUT2), .B(G113), .Z(new_n423));
  XNOR2_X1  g237(.A(G116), .B(G119), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT65), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n427), .A3(new_n424), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n423), .ZN(new_n430));
  INV_X1    g244(.A(new_n424), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n263), .A3(new_n272), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n424), .A2(KEYINPUT5), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n394), .A2(G119), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n435), .B(G113), .C1(KEYINPUT5), .C2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n223), .A2(new_n429), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G122), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(new_n440), .A3(new_n438), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n439), .A2(new_n445), .A3(new_n441), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n231), .A2(new_n337), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n253), .A2(G125), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n321), .A2(G224), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n449), .B(new_n450), .Z(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n440), .B(KEYINPUT8), .Z(new_n453));
  NAND2_X1  g267(.A1(new_n429), .A2(new_n437), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n228), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n455), .B2(new_n438), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n450), .A2(KEYINPUT7), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n448), .B2(KEYINPUT82), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n449), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n447), .B(new_n448), .C1(KEYINPUT82), .C2(new_n457), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n462), .B2(new_n443), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n452), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT83), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n466), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n452), .A2(new_n468), .A3(new_n463), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G214), .B1(G237), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n422), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n302), .A2(new_n310), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT91), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n388), .B1(G234), .B2(new_n285), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n405), .A2(G119), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n479), .B(new_n480), .C1(G119), .C2(new_n405), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT24), .B(G110), .ZN(new_n482));
  OAI22_X1  g296(.A1(new_n317), .A2(new_n318), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n405), .A2(G119), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT23), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n485), .A2(KEYINPUT72), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n486), .B2(new_n478), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT72), .B(KEYINPUT23), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n487), .B1(new_n478), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G110), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT73), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(KEYINPUT73), .A3(G110), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n483), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n481), .A2(new_n482), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n489), .B2(G110), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n316), .A3(new_n341), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT22), .B(G137), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n297), .A2(new_n376), .A3(G953), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n499), .B(new_n500), .Z(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n501), .ZN(new_n503));
  INV_X1    g317(.A(new_n498), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n503), .B1(new_n504), .B2(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT25), .B1(new_n507), .B2(new_n285), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n506), .A2(new_n509), .A3(G902), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n477), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n477), .A2(G902), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n426), .A2(new_n428), .B1(new_n431), .B2(new_n430), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n244), .A2(new_n273), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n235), .A2(G137), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n237), .A2(G134), .ZN(new_n519));
  OAI21_X1  g333(.A(G131), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n240), .B2(new_n326), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT67), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n229), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n193), .B1(new_n524), .B2(new_n405), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n206), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n243), .A2(KEYINPUT67), .A3(new_n520), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT28), .B1(new_n517), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n273), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT66), .B1(new_n244), .B2(new_n273), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n528), .B(new_n515), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n243), .B(new_n520), .C1(new_n230), .C2(new_n205), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n516), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n433), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n529), .B1(new_n536), .B2(KEYINPUT28), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G101), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n320), .A2(new_n321), .A3(G210), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n532), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n528), .B(KEYINPUT30), .C1(new_n530), .C2(new_n531), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT68), .B1(new_n534), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT66), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n516), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n273), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n554), .A2(KEYINPUT68), .A3(KEYINPUT30), .A4(new_n528), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n546), .B1(new_n556), .B2(new_n433), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT31), .B1(new_n557), .B2(new_n543), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n515), .B1(new_n550), .B2(new_n555), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT31), .ZN(new_n560));
  NOR4_X1   g374(.A1(new_n559), .A2(new_n560), .A3(new_n546), .A4(new_n542), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n545), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G472), .A2(G902), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT32), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT70), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT70), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n567), .B(KEYINPUT32), .C1(new_n562), .C2(new_n563), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(KEYINPUT32), .A3(new_n563), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT29), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n557), .A2(new_n571), .A3(new_n542), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n537), .A2(new_n571), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n543), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n433), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n532), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n529), .B1(new_n577), .B2(KEYINPUT28), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n571), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n572), .B(new_n285), .C1(new_n574), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n570), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n514), .B1(new_n569), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n302), .A2(new_n310), .A3(new_n584), .A4(new_n474), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n476), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  AND2_X1   g401(.A1(new_n302), .A2(new_n310), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n387), .A2(G902), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n412), .A2(new_n415), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n412), .B2(new_n415), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT92), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(KEYINPUT92), .B(new_n589), .C1(new_n591), .C2(new_n592), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT93), .B(G478), .Z(new_n598));
  NAND2_X1  g412(.A1(new_n418), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n374), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n469), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n468), .B1(new_n452), .B2(new_n463), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n472), .B(new_n386), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n556), .A2(new_n433), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n532), .A3(new_n543), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n560), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n557), .A2(KEYINPUT31), .A3(new_n543), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n544), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(G472), .B1(new_n610), .B2(G902), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n564), .ZN(new_n612));
  INV_X1    g426(.A(new_n514), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n588), .A2(new_n605), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  OAI22_X1  g431(.A1(new_n417), .A2(new_n420), .B1(new_n351), .B2(new_n352), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n367), .ZN(new_n620));
  INV_X1    g434(.A(new_n365), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n348), .A3(new_n363), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n620), .B1(new_n622), .B2(new_n350), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n369), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n371), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT94), .B1(new_n604), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n618), .B1(new_n371), .B2(new_n624), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n473), .B1(new_n467), .B2(new_n469), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .A4(new_n386), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n588), .A2(new_n614), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n210), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT95), .B(KEYINPUT35), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NAND2_X1  g450(.A1(new_n495), .A2(new_n498), .ZN(new_n637));
  OR3_X1    g451(.A1(new_n637), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n637), .B1(KEYINPUT36), .B2(new_n503), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n512), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n511), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n612), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT96), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n476), .A3(new_n585), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT97), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n645), .B(new_n647), .ZN(G12));
  NAND2_X1  g462(.A1(new_n564), .A2(new_n565), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n567), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT32), .B1(new_n562), .B2(new_n563), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT70), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n582), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n642), .A2(new_n629), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n321), .A2(G900), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n384), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT98), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(KEYINPUT98), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n657), .A2(new_n377), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n628), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n653), .A2(new_n302), .A3(new_n310), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XOR2_X1   g478(.A(new_n659), .B(KEYINPUT39), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n588), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n577), .A2(new_n542), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(KEYINPUT99), .Z(new_n670));
  INV_X1    g484(.A(new_n607), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n285), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G472), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n650), .A2(new_n652), .A3(new_n570), .A4(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n470), .B(KEYINPUT38), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n373), .B1(new_n623), .B2(new_n369), .ZN(new_n677));
  INV_X1    g491(.A(new_n353), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n421), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n676), .A2(new_n472), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n675), .A2(new_n642), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n667), .A2(new_n668), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NAND4_X1  g497(.A1(new_n600), .A2(new_n629), .A3(new_n642), .A4(new_n660), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n569), .B2(new_n582), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n588), .A2(KEYINPUT100), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n374), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n597), .A2(new_n599), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n688), .A3(new_n660), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n654), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n653), .A2(new_n302), .A3(new_n310), .A4(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  OAI21_X1  g509(.A(new_n285), .B1(new_n288), .B2(new_n290), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT101), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n699), .A3(G469), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n307), .A2(new_n308), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n301), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT102), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n698), .A2(new_n700), .B1(new_n308), .B2(new_n307), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n301), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n653), .A2(new_n613), .A3(new_n605), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT41), .B(G113), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NOR2_X1   g526(.A1(new_n703), .A2(KEYINPUT102), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n706), .B1(new_n705), .B2(new_n301), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n653), .A2(new_n613), .A3(new_n632), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT103), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n653), .A2(new_n613), .A3(new_n632), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n708), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  AND4_X1   g536(.A1(new_n301), .A2(new_n701), .A3(new_n702), .A4(new_n629), .ZN(new_n723));
  INV_X1    g537(.A(new_n642), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n422), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n653), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NAND2_X1  g541(.A1(new_n608), .A2(new_n609), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n578), .A2(new_n543), .ZN(new_n729));
  AOI211_X1 g543(.A(G472), .B(G902), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n611), .A2(KEYINPUT104), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n732), .B(G472), .C1(new_n610), .C2(G902), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n730), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n679), .A2(new_n629), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n385), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n613), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n708), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n738), .B(G122), .Z(G24));
  INV_X1    g553(.A(new_n689), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n723), .A2(new_n642), .A3(new_n740), .A4(new_n734), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n467), .A2(new_n301), .A3(new_n472), .A4(new_n469), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n295), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT105), .B1(new_n309), .B2(new_n744), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n583), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n564), .B2(new_n565), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n570), .A2(new_n581), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n651), .A2(new_n751), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n514), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n748), .A3(new_n740), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n749), .A2(new_n750), .B1(new_n757), .B2(KEYINPUT42), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  INV_X1    g573(.A(new_n661), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n583), .A2(new_n760), .A3(new_n748), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT107), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n583), .A2(new_n748), .A3(new_n763), .A4(new_n760), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  INV_X1    g580(.A(new_n284), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n767), .A2(KEYINPUT45), .ZN(new_n768));
  OAI21_X1  g582(.A(G469), .B1(new_n767), .B2(KEYINPUT45), .ZN(new_n769));
  OAI22_X1  g583(.A1(new_n768), .A2(new_n769), .B1(new_n187), .B2(new_n285), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n702), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n771), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n301), .B(new_n665), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n688), .A2(new_n374), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT43), .Z(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n642), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(new_n612), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(KEYINPUT109), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n471), .A2(new_n472), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n783), .B(new_n785), .C1(new_n782), .C2(new_n781), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT109), .B1(new_n781), .B2(new_n782), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n777), .B1(new_n788), .B2(KEYINPUT110), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(KEYINPUT110), .B2(new_n788), .ZN(new_n790));
  XNOR2_X1  g604(.A(KEYINPUT111), .B(G137), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G39));
  OAI21_X1  g606(.A(new_n301), .B1(new_n774), .B2(new_n776), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n653), .A2(new_n613), .A3(new_n689), .A4(new_n784), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n765), .A2(new_n758), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n726), .B1(new_n708), .B2(new_n709), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n738), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(new_n721), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n374), .A2(new_n421), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n374), .B2(new_n688), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n604), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n588), .A2(new_n614), .A3(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n645), .A2(new_n586), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n421), .A2(new_n678), .A3(new_n660), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n511), .B2(new_n641), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n472), .A3(new_n471), .A4(new_n625), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n569), .B2(new_n582), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n588), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n812), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n642), .A2(new_n625), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n784), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n653), .A2(new_n302), .A3(new_n310), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT113), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n734), .A2(new_n642), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n689), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n816), .A2(new_n821), .B1(new_n823), .B2(new_n748), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n802), .A2(new_n805), .A3(new_n810), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n691), .B(KEYINPUT100), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n309), .A2(new_n735), .A3(new_n300), .A4(new_n659), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n674), .A3(new_n724), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n741), .A2(new_n828), .A3(new_n663), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT114), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n741), .A2(new_n828), .A3(new_n663), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n694), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT52), .B1(new_n826), .B2(new_n829), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n831), .A2(new_n694), .A3(new_n832), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n832), .B1(new_n831), .B2(new_n694), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n804), .A2(new_n824), .A3(new_n721), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n765), .A2(new_n758), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n830), .A2(KEYINPUT52), .A3(new_n833), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n846), .A3(new_n847), .A4(new_n810), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n838), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n801), .B1(new_n839), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n848), .A2(new_n838), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n848), .A2(new_n854), .A3(new_n838), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n835), .A2(new_n856), .A3(KEYINPUT53), .A4(new_n836), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n645), .A2(new_n586), .A3(new_n809), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n844), .A2(new_n845), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n843), .A4(new_n836), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n853), .A2(new_n855), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n851), .B1(new_n801), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n779), .A2(new_n613), .A3(new_n378), .A4(new_n734), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n784), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n705), .A2(new_n300), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n866), .B1(new_n797), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT117), .B1(new_n795), .B2(new_n796), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n864), .A2(new_n472), .A3(new_n676), .A4(new_n703), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT50), .Z(new_n872));
  INV_X1    g686(.A(new_n705), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n873), .A2(new_n377), .A3(new_n744), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n779), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n822), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n613), .A3(new_n675), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n877), .A2(new_n687), .A3(new_n688), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n872), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n870), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n880), .A2(KEYINPUT51), .ZN(new_n881));
  INV_X1    g695(.A(new_n866), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n865), .B1(new_n797), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n879), .A2(KEYINPUT51), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n723), .ZN(new_n885));
  OAI221_X1 g699(.A(new_n375), .B1(new_n864), .B2(new_n885), .C1(new_n877), .C2(new_n601), .ZN(new_n886));
  INV_X1    g700(.A(new_n756), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n875), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT118), .Z(new_n889));
  INV_X1    g703(.A(KEYINPUT48), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n889), .A2(KEYINPUT119), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n886), .B(new_n891), .C1(new_n889), .C2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n863), .A2(new_n881), .A3(new_n884), .A4(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n873), .A2(KEYINPUT49), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT112), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n873), .A2(KEYINPUT49), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n613), .A2(new_n301), .A3(new_n472), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n674), .A2(new_n676), .A3(new_n778), .A4(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n895), .A2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n862), .A2(new_n285), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n466), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n444), .A2(new_n446), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n451), .ZN(new_n907));
  XOR2_X1   g721(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n904), .A2(new_n905), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n904), .B2(new_n905), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n321), .A2(G952), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G51));
  AND3_X1   g727(.A1(new_n848), .A2(new_n854), .A3(new_n838), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n854), .B1(new_n848), .B2(new_n838), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n860), .B(new_n856), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT54), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n857), .A2(new_n861), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n919), .B(new_n801), .C1(new_n914), .C2(new_n915), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n187), .A2(new_n285), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT57), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n306), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n768), .A2(new_n769), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n903), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n912), .B1(new_n925), .B2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n350), .A3(new_n622), .ZN(new_n930));
  INV_X1    g744(.A(new_n912), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .A4(new_n366), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G60));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT59), .Z(new_n935));
  AOI21_X1  g749(.A(KEYINPUT53), .B1(new_n835), .B2(new_n836), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT54), .B1(new_n936), .B2(new_n849), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n920), .B2(new_n937), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n591), .A2(new_n592), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT122), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n939), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(new_n935), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT121), .B1(new_n921), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n944));
  INV_X1    g758(.A(new_n942), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n944), .B(new_n945), .C1(new_n918), .C2(new_n920), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n940), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n941), .B1(new_n863), .B2(new_n935), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n931), .B1(new_n948), .B2(KEYINPUT122), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n862), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n912), .B1(new_n953), .B2(new_n640), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n507), .B2(new_n953), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT123), .B1(new_n953), .B2(new_n640), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI221_X1 g772(.A(new_n954), .B1(new_n507), .B2(new_n953), .C1(new_n956), .C2(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(G66));
  OAI22_X1  g774(.A1(new_n380), .A2(new_n382), .B1(G224), .B2(new_n321), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT124), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n805), .A2(new_n810), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n321), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n906), .B1(new_n381), .B2(G953), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(G69));
  AOI21_X1  g780(.A(new_n655), .B1(new_n189), .B2(G953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n790), .A2(new_n799), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n694), .A2(new_n663), .A3(new_n741), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n682), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n973));
  INV_X1    g787(.A(new_n583), .ZN(new_n974));
  NOR4_X1   g788(.A1(new_n666), .A2(new_n974), .A3(new_n784), .A4(new_n807), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT125), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n969), .A2(new_n972), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n556), .B(new_n360), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n321), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n655), .B(KEYINPUT126), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n802), .A2(new_n970), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n777), .A2(new_n735), .A3(new_n887), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT127), .Z(new_n985));
  OR3_X1    g799(.A1(new_n968), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n982), .B1(new_n986), .B2(new_n321), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n967), .B1(new_n980), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n967), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n986), .A2(new_n321), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n979), .B(new_n989), .C1(new_n990), .C2(new_n982), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n977), .B2(new_n963), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n557), .A2(new_n542), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n559), .A2(new_n546), .A3(new_n543), .ZN(new_n998));
  NOR4_X1   g812(.A1(new_n968), .A2(new_n985), .A3(new_n963), .A4(new_n983), .ZN(new_n999));
  INV_X1    g813(.A(new_n994), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n997), .A2(new_n931), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n936), .A2(new_n849), .ZN(new_n1003));
  NOR4_X1   g817(.A1(new_n1003), .A2(new_n998), .A3(new_n996), .A4(new_n1000), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1002), .A2(new_n1004), .ZN(G57));
endmodule


