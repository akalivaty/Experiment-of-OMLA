//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n210), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n215), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n212), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n215), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT64), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n223), .B(new_n227), .C1(KEYINPUT1), .C2(new_n222), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G13), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(G1), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n202), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n214), .A2(G33), .B1(G1), .B2(G13), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n249), .B1(G1), .B2(new_n210), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n248), .B1(new_n251), .B2(new_n202), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n210), .A2(G33), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n249), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT9), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G223), .A3(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G222), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n263), .B1(new_n264), .B2(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n213), .A2(G274), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT65), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT65), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G41), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G41), .A2(G45), .ZN(new_n282));
  OAI22_X1  g0082(.A1(new_n281), .A2(new_n209), .B1(new_n282), .B2(G1), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n270), .A2(KEYINPUT66), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n280), .B1(new_n288), .B2(G226), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n272), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G200), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n261), .B(new_n291), .C1(new_n292), .C2(new_n290), .ZN(new_n293));
  XOR2_X1   g0093(.A(new_n293), .B(KEYINPUT10), .Z(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(G169), .B2(new_n290), .ZN(new_n297));
  INV_X1    g0097(.A(new_n260), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G68), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n246), .A2(G20), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT12), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n253), .A2(KEYINPUT68), .A3(G50), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n304), .B1(new_n210), .B2(G68), .C1(new_n264), .C2(new_n255), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT68), .B1(new_n253), .B2(G50), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n258), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT11), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n303), .B1(new_n301), .B2(new_n250), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n307), .A2(new_n308), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n270), .A2(KEYINPUT66), .A3(new_n286), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT66), .B1(new_n270), .B2(new_n286), .ZN(new_n313));
  OAI21_X1  g0113(.A(G238), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n273), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n275), .A2(new_n277), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(G45), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(KEYINPUT67), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G33), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n320), .A2(new_n322), .A3(G232), .A4(G1698), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n320), .A2(new_n322), .A3(G226), .A4(new_n265), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n271), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n318), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT67), .B1(new_n314), .B2(new_n317), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT13), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT67), .ZN(new_n331));
  INV_X1    g0131(.A(G238), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n285), .B2(new_n287), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(new_n280), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(new_n318), .A4(new_n327), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n330), .A2(new_n292), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(G200), .B1(new_n330), .B2(new_n336), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n311), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT69), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT69), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n311), .C1(new_n337), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n256), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n250), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n247), .A2(new_n256), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G58), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n301), .ZN(new_n350));
  OAI21_X1  g0150(.A(G20), .B1(new_n350), .B2(new_n201), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n253), .A2(G159), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n262), .B2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n320), .A2(new_n322), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n353), .B1(new_n358), .B2(G68), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n249), .B1(new_n359), .B2(KEYINPUT16), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT73), .B1(new_n321), .B2(G33), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT73), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(new_n319), .A3(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n364), .A3(new_n322), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n354), .A2(G20), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n301), .B1(new_n367), .B2(new_n355), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n361), .B1(new_n368), .B2(new_n353), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n348), .B1(new_n360), .B2(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n320), .A2(new_n322), .A3(G223), .A4(new_n265), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n320), .A2(new_n322), .A3(G226), .A4(G1698), .ZN(new_n372));
  INV_X1    g0172(.A(G87), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(new_n372), .C1(new_n319), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n271), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n270), .A2(G232), .A3(new_n286), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n317), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n377), .A3(new_n295), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n317), .A2(new_n376), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n271), .B2(new_n374), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n378), .B1(new_n380), .B2(G169), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT18), .B1(new_n370), .B2(new_n381), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n262), .A2(new_n354), .A3(G20), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT7), .B1(new_n356), .B2(new_n210), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n353), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n369), .A2(new_n387), .A3(new_n258), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n375), .A2(new_n377), .A3(new_n292), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n380), .B2(G200), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n390), .A3(new_n347), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(new_n347), .ZN(new_n394));
  INV_X1    g0194(.A(new_n381), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n370), .A2(KEYINPUT17), .A3(new_n390), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n382), .A2(new_n393), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n251), .A2(G77), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(G77), .B2(new_n247), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT15), .B(G87), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n403), .A2(new_n255), .B1(new_n210), .B2(new_n264), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n253), .B2(new_n344), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(new_n249), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n262), .A2(G238), .A3(G1698), .ZN(new_n409));
  INV_X1    g0209(.A(G107), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n409), .B1(new_n410), .B2(new_n262), .C1(new_n266), .C2(new_n232), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n271), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n280), .B1(new_n288), .B2(G244), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n292), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  INV_X1    g0215(.A(G200), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n408), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(G169), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n412), .A2(G179), .A3(new_n413), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n407), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n300), .A2(new_n343), .A3(new_n400), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n330), .A2(G179), .A3(new_n336), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT71), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT71), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n330), .A2(new_n426), .A3(G179), .A4(new_n336), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n326), .A2(new_n271), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n280), .B1(new_n288), .B2(G238), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(KEYINPUT67), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n335), .B1(new_n431), .B2(new_n334), .ZN(new_n432));
  INV_X1    g0232(.A(new_n336), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT70), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT14), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n437));
  INV_X1    g0237(.A(G169), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n330), .B2(new_n336), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n428), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT72), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT72), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n428), .A2(new_n436), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n311), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n423), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G116), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n247), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n213), .A2(G33), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n249), .A2(new_n247), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n452), .B2(new_n448), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n319), .A2(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  AOI21_X1  g0255(.A(G20), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n210), .A2(new_n448), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n258), .B(KEYINPUT20), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT20), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n456), .A2(new_n457), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(new_n249), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n438), .B1(new_n453), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n262), .A2(G264), .A3(G1698), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n262), .A2(G257), .A3(new_n265), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n356), .A2(G303), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT79), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT79), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n464), .A2(new_n465), .A3(new_n469), .A4(new_n466), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n271), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n213), .B(G45), .C1(new_n472), .C2(G41), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n316), .B2(new_n472), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n271), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n475), .A2(G270), .B1(G274), .B2(new_n474), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n463), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n463), .A2(new_n477), .A3(KEYINPUT21), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n453), .A2(new_n462), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(G179), .A3(new_n471), .A4(new_n476), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT6), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n410), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G97), .A2(G107), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n410), .A2(KEYINPUT6), .A3(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n384), .B1(new_n365), .B2(new_n366), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(new_n410), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n258), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n247), .A2(new_n486), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n452), .B2(new_n486), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .A4(new_n265), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n320), .A2(new_n322), .A3(G244), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n455), .C1(new_n500), .C2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n262), .A2(G250), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n265), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n271), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT74), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n475), .A2(G257), .B1(G274), .B2(new_n474), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT74), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(new_n271), .C1(new_n501), .C2(new_n503), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n498), .B1(G200), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT75), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n504), .A2(new_n511), .A3(new_n506), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n504), .B2(new_n506), .ZN(new_n514));
  OAI21_X1  g0314(.A(G190), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n504), .A2(new_n506), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT75), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n438), .A3(new_n512), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n498), .C1(G179), .C2(new_n509), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n477), .A2(G190), .ZN(new_n521));
  AOI21_X1  g0321(.A(G200), .B1(new_n471), .B2(new_n476), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n462), .B(new_n453), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n484), .A2(new_n516), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n262), .A2(new_n210), .A3(G68), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT76), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G87), .A2(G97), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(new_n410), .B1(new_n325), .B2(new_n210), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n210), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n529), .A2(new_n530), .B1(new_n325), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n262), .A2(KEYINPUT76), .A3(new_n210), .A4(G68), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n527), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n258), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n403), .A2(G20), .A3(new_n246), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n452), .A2(G87), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n315), .A2(G45), .ZN(new_n539));
  OAI21_X1  g0339(.A(G250), .B1(new_n279), .B2(G1), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n271), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n262), .A2(G244), .A3(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G116), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n266), .C2(new_n332), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n544), .B2(new_n271), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G200), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT78), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n538), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n545), .A2(new_n416), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT78), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n546), .A2(new_n292), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n403), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n452), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n535), .A2(new_n536), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT77), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n545), .A2(G179), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n438), .B2(new_n545), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n246), .A2(G20), .A3(new_n410), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT25), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n567), .A2(KEYINPUT25), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n451), .C2(new_n410), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n543), .A2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n210), .B2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n410), .A2(KEYINPUT23), .A3(G20), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n262), .A2(new_n210), .A3(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n262), .A2(new_n580), .A3(new_n210), .A4(G87), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n577), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g0382(.A(KEYINPUT80), .B(KEYINPUT24), .Z(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n258), .B1(new_n582), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n571), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT81), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n262), .A2(G257), .A3(G1698), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G294), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n502), .C2(G1698), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n271), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n475), .A2(G264), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n474), .A2(G274), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n596), .A2(new_n438), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(G179), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n571), .B(KEYINPUT81), .C1(new_n585), .C2(new_n586), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n589), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n586), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n570), .B1(new_n602), .B2(new_n584), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n596), .A2(new_n416), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(G190), .B2(new_n596), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n556), .A2(new_n566), .A3(new_n601), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n524), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n447), .A2(new_n608), .ZN(G372));
  NAND2_X1  g0409(.A1(new_n443), .A2(new_n445), .ZN(new_n610));
  INV_X1    g0410(.A(new_n311), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n339), .ZN(new_n613));
  INV_X1    g0413(.A(new_n421), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n612), .B(KEYINPUT83), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n446), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n615), .A2(new_n393), .A3(new_n398), .A4(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n382), .A2(new_n397), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n294), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n299), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n554), .A2(new_n550), .A3(new_n551), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n603), .A2(new_n597), .A3(new_n598), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n516), .B(new_n606), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  AOI211_X1 g0427(.A(KEYINPUT26), .B(new_n624), .C1(new_n627), .C2(new_n520), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n565), .B(KEYINPUT82), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n559), .ZN(new_n630));
  INV_X1    g0430(.A(new_n565), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n562), .B2(new_n561), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n554), .B1(new_n549), .B2(new_n552), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n520), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n447), .B1(new_n628), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n623), .A2(new_n637), .ZN(G369));
  INV_X1    g0438(.A(new_n246), .ZN(new_n639));
  OR3_X1    g0439(.A1(new_n639), .A2(KEYINPUT27), .A3(G20), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT27), .B1(new_n639), .B2(G20), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g0443(.A(KEYINPUT84), .B(G343), .Z(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n589), .A2(new_n600), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n601), .A2(new_n647), .A3(new_n606), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n601), .B2(new_n645), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(KEYINPUT85), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(KEYINPUT85), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n523), .A2(new_n481), .A3(new_n480), .A4(new_n483), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n482), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n625), .A2(new_n654), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G330), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n484), .A2(new_n646), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n650), .B2(new_n651), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n626), .A2(new_n645), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(G399));
  NAND2_X1  g0466(.A1(new_n224), .A2(new_n278), .ZN(new_n667));
  NOR4_X1   g0467(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G1), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n207), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n645), .B1(new_n628), .B2(new_n636), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n627), .A2(new_n520), .ZN(new_n674));
  INV_X1    g0474(.A(new_n624), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n635), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n630), .ZN(new_n677));
  OR3_X1    g0477(.A1(new_n520), .A2(new_n632), .A3(new_n633), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(KEYINPUT26), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n646), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT88), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT29), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n673), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n624), .B1(new_n603), .B2(new_n605), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n685), .A2(new_n516), .A3(new_n520), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n484), .A2(new_n601), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n677), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n634), .A2(KEYINPUT26), .B1(new_n520), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n646), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(KEYINPUT29), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n545), .B(KEYINPUT86), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n596), .A2(new_n295), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n695), .A2(new_n509), .A3(new_n696), .A4(new_n477), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n518), .A2(new_n512), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n593), .A2(new_n594), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n477), .A2(new_n700), .A3(new_n564), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n699), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n698), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n694), .B1(new_n706), .B2(new_n645), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT87), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n703), .A2(new_n705), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n645), .B1(new_n710), .B2(new_n697), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n608), .A2(new_n645), .B1(new_n711), .B2(KEYINPUT31), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n708), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n693), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n671), .B1(new_n718), .B2(G1), .ZN(G364));
  NOR2_X1   g0519(.A1(new_n245), .A2(G20), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G45), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n667), .A2(G1), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n657), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n724), .B2(new_n659), .ZN(new_n725));
  INV_X1    g0525(.A(new_n722), .ZN(new_n726));
  OR3_X1    g0526(.A1(KEYINPUT89), .A2(G13), .A3(G33), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT89), .B1(G13), .B2(G33), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n723), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n210), .A2(new_n292), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n416), .A2(G179), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT90), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(KEYINPUT90), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G87), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n210), .B1(new_n742), .B2(G190), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G97), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n295), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n734), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n210), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n735), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n750), .A2(new_n349), .B1(new_n752), .B2(new_n410), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n295), .A2(new_n416), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n751), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n749), .A2(new_n751), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n301), .B1(new_n756), .B2(new_n264), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n734), .A2(new_n754), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n262), .B1(new_n758), .B2(new_n202), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n753), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n751), .A2(new_n742), .ZN(new_n761));
  INV_X1    g0561(.A(G159), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT32), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n741), .A2(new_n748), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n761), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n262), .B1(new_n766), .B2(G329), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n767), .B1(new_n768), .B2(new_n752), .C1(new_n769), .C2(new_n756), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(G303), .B2(new_n740), .ZN(new_n771));
  INV_X1    g0571(.A(new_n758), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n747), .A2(G294), .B1(G326), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT92), .ZN(new_n774));
  XOR2_X1   g0574(.A(KEYINPUT33), .B(G317), .Z(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n755), .B1(new_n750), .B2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT93), .Z(new_n778));
  NAND3_X1  g0578(.A1(new_n771), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n773), .A2(KEYINPUT92), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n765), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n209), .B1(G20), .B2(new_n438), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n224), .A2(G355), .A3(new_n262), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n208), .A2(G45), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n240), .B2(G45), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n224), .A2(new_n356), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n784), .B1(G116), .B2(new_n224), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n731), .A2(new_n782), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n726), .B1(new_n733), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n725), .A2(new_n792), .ZN(G396));
  NAND2_X1  g0593(.A1(new_n740), .A2(G107), .ZN(new_n794));
  INV_X1    g0594(.A(G303), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n758), .A2(new_n795), .B1(new_n752), .B2(new_n373), .ZN(new_n796));
  INV_X1    g0596(.A(new_n750), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n262), .B(new_n796), .C1(G294), .C2(new_n797), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n755), .A2(new_n768), .B1(new_n761), .B2(new_n769), .ZN(new_n799));
  INV_X1    g0599(.A(new_n756), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(G116), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n794), .A2(new_n798), .A3(new_n748), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n758), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G143), .ZN(new_n805));
  INV_X1    g0605(.A(G150), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n805), .A2(new_n750), .B1(new_n755), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n804), .B(new_n807), .C1(G159), .C2(new_n800), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n349), .B2(new_n746), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n262), .B1(new_n752), .B2(new_n301), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G132), .B2(new_n766), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n812), .B1(new_n202), .B2(new_n739), .C1(new_n808), .C2(KEYINPUT34), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n802), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n782), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n729), .A2(new_n782), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT94), .Z(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n722), .B1(new_n818), .B2(new_n264), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n418), .B1(new_n408), .B2(new_n646), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n421), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n421), .A2(new_n645), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n815), .B(new_n819), .C1(new_n824), .C2(new_n730), .ZN(new_n825));
  INV_X1    g0625(.A(new_n824), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n673), .A2(new_n682), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n680), .A2(new_n824), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n716), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n722), .B1(new_n829), .B2(new_n716), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n825), .B1(new_n831), .B2(new_n832), .ZN(G384));
  OAI211_X1 g0633(.A(G116), .B(new_n211), .C1(new_n491), .C2(KEYINPUT35), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(KEYINPUT35), .B2(new_n491), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT36), .ZN(new_n836));
  OR3_X1    g0636(.A1(new_n207), .A2(new_n264), .A3(new_n350), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n202), .A2(G68), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n213), .B(G13), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT95), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n443), .A2(new_n445), .A3(new_n343), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n311), .A2(new_n645), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n843), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n339), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n610), .B2(new_n611), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n841), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n842), .A2(new_n843), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n849), .B(KEYINPUT95), .C1(new_n446), .C2(new_n846), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n826), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT101), .B1(new_n712), .B2(new_n707), .ZN(new_n852));
  INV_X1    g0652(.A(new_n524), .ZN(new_n853));
  INV_X1    g0653(.A(new_n607), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(new_n854), .A3(new_n645), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n711), .A2(KEYINPUT31), .ZN(new_n856));
  AND4_X1   g0656(.A1(KEYINPUT101), .A2(new_n855), .A3(new_n856), .A4(new_n707), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT102), .Z(new_n860));
  NOR2_X1   g0660(.A1(new_n370), .A2(new_n642), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n399), .A2(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n388), .A2(new_n347), .B1(new_n381), .B2(new_n642), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n864), .A2(KEYINPUT97), .A3(KEYINPUT37), .A4(new_n391), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n391), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n863), .B2(KEYINPUT97), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n862), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT98), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n864), .A2(new_n873), .A3(new_n391), .ZN(new_n874));
  INV_X1    g0674(.A(new_n391), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n361), .A2(KEYINPUT96), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n359), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n301), .B1(new_n355), .B2(new_n357), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT96), .B(new_n361), .C1(new_n878), .C2(new_n353), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n258), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n381), .B1(new_n880), .B2(new_n347), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n642), .B1(new_n880), .B2(new_n347), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n875), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n874), .B1(new_n883), .B2(new_n873), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n399), .A2(new_n882), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n872), .A2(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n399), .A2(new_n861), .B1(new_n866), .B2(new_n867), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n888), .B2(new_n865), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n889), .A2(new_n870), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n891), .A2(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n885), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n871), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n886), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n851), .A2(new_n895), .A3(new_n858), .ZN(new_n896));
  XOR2_X1   g0696(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n897));
  AOI22_X1  g0697(.A1(new_n860), .A2(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n858), .A2(new_n447), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n898), .B(new_n899), .Z(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n658), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n872), .A2(new_n886), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n889), .A2(new_n870), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT99), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(KEYINPUT99), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n612), .A2(new_n646), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n620), .A2(new_n643), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n848), .A2(new_n850), .B1(new_n828), .B2(new_n822), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n916), .B2(new_n895), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n684), .A2(new_n447), .A3(new_n692), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n623), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  OAI22_X1  g0721(.A1(new_n901), .A2(new_n921), .B1(new_n213), .B2(new_n720), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n901), .A2(new_n921), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n840), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT103), .ZN(G367));
  NOR2_X1   g0725(.A1(new_n538), .A2(new_n645), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n630), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n677), .A2(new_n624), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n926), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n498), .A2(new_n646), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n516), .A2(new_n520), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n520), .B2(new_n645), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n663), .B(new_n935), .C1(new_n650), .C2(new_n651), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(KEYINPUT104), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(KEYINPUT104), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n934), .A2(new_n601), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n646), .B1(new_n940), .B2(new_n520), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n936), .B2(KEYINPUT42), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n932), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n943), .A2(new_n932), .A3(new_n944), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n661), .A2(new_n935), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n667), .B(KEYINPUT41), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n935), .B1(new_n664), .B2(new_n665), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT44), .Z(new_n954));
  NAND3_X1  g0754(.A1(new_n664), .A2(new_n665), .A3(new_n935), .ZN(new_n955));
  XOR2_X1   g0755(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n662), .B1(new_n958), .B2(KEYINPUT106), .ZN(new_n959));
  INV_X1    g0759(.A(new_n958), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT106), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n961), .A3(new_n661), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n652), .B1(new_n484), .B2(new_n646), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(new_n664), .C1(KEYINPUT107), .C2(new_n659), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n659), .A2(KEYINPUT107), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(new_n717), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n959), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n952), .B1(new_n968), .B2(new_n718), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n721), .A2(G1), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n951), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n789), .B1(new_n224), .B2(new_n403), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n236), .A2(new_n787), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n726), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n740), .A2(G58), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n758), .A2(new_n805), .B1(new_n755), .B2(new_n762), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n356), .B(new_n976), .C1(G50), .C2(new_n800), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n747), .A2(G68), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n752), .A2(new_n264), .B1(new_n761), .B2(new_n803), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G150), .B2(new_n797), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n975), .A2(new_n977), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n739), .A2(new_n448), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT46), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n750), .A2(new_n795), .B1(new_n756), .B2(new_n768), .ZN(new_n984));
  INV_X1    g0784(.A(new_n752), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n984), .B1(G97), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(G294), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n758), .A2(new_n769), .B1(new_n755), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n262), .B(new_n988), .C1(G317), .C2(new_n766), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n983), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n982), .A2(KEYINPUT46), .B1(new_n410), .B2(new_n746), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT47), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n994), .A2(new_n782), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n993), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n974), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n930), .B2(new_n732), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n971), .A2(new_n998), .ZN(G387));
  INV_X1    g0799(.A(new_n789), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n224), .A2(new_n262), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n1001), .A2(new_n668), .B1(G107), .B2(new_n224), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n233), .A2(G45), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n279), .B1(new_n301), .B2(new_n264), .C1(new_n668), .C2(KEYINPUT108), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(KEYINPUT108), .B2(new_n668), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n256), .A2(G50), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT50), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n787), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1002), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n755), .A2(new_n256), .B1(new_n756), .B2(new_n301), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT109), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n740), .A2(G77), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n747), .A2(new_n557), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n262), .B1(new_n752), .B2(new_n486), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n758), .A2(new_n762), .B1(new_n750), .B2(new_n202), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G150), .C2(new_n766), .ZN(new_n1017));
  AND4_X1   g0817(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n747), .A2(G283), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G322), .A2(new_n772), .B1(new_n800), .B2(G303), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n769), .B2(new_n755), .C1(new_n1021), .C2(new_n750), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1019), .B1(new_n987), .B2(new_n739), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT110), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1029));
  INV_X1    g0829(.A(G326), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n356), .B1(new_n761), .B2(new_n1030), .C1(new_n448), .C2(new_n752), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1028), .B2(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1018), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n782), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n726), .B1(new_n1000), .B2(new_n1009), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n652), .B2(new_n731), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n966), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n970), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1037), .A2(new_n718), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n667), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n966), .B2(new_n717), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1038), .B1(new_n1039), .B2(new_n1041), .ZN(G393));
  XNOR2_X1  g0842(.A(new_n958), .B(new_n661), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(new_n967), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1044), .A2(new_n667), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n968), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(new_n970), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n935), .A2(new_n732), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT111), .Z(new_n1049));
  OAI21_X1  g0849(.A(new_n789), .B1(new_n486), .B2(new_n224), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n243), .A2(new_n787), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n726), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n356), .B1(new_n752), .B2(new_n410), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n755), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G303), .A2(new_n1054), .B1(new_n800), .B2(G294), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n776), .B2(new_n761), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1053), .B(new_n1056), .C1(G116), .C2(new_n747), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT52), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n758), .A2(new_n1021), .B1(new_n750), .B2(new_n769), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n740), .A2(G283), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1057), .B(new_n1060), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n755), .A2(new_n202), .B1(new_n756), .B2(new_n256), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n356), .B(new_n1062), .C1(G87), .C2(new_n985), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n758), .A2(new_n806), .B1(new_n750), .B2(new_n762), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT51), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(new_n264), .C2(new_n746), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n739), .A2(new_n301), .B1(new_n805), .B2(new_n761), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT112), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1061), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1052), .B1(new_n1069), .B2(new_n782), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1049), .A2(new_n1070), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1046), .A2(new_n1047), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G390));
  AND3_X1   g0873(.A1(new_n905), .A2(KEYINPUT99), .A3(new_n906), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT99), .B1(new_n905), .B2(new_n906), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n916), .A2(new_n913), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n851), .A2(new_n715), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n821), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n823), .B1(new_n691), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n850), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n846), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n612), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT95), .B1(new_n1083), .B2(new_n849), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1080), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n913), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n891), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT113), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1079), .B1(new_n848), .B2(new_n850), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT113), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1090), .A2(new_n1091), .A3(new_n1087), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1076), .B(new_n1077), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n826), .A2(new_n658), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n852), .B2(new_n857), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1085), .A2(KEYINPUT113), .A3(new_n1088), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1091), .B1(new_n1090), .B2(new_n1087), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n828), .A2(new_n822), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1086), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1100), .A2(new_n1101), .B1(new_n1104), .B2(new_n911), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1099), .B1(new_n1105), .B2(KEYINPUT114), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1076), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT114), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1094), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n970), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n722), .B1(new_n818), .B2(new_n256), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n741), .A2(new_n356), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT118), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n746), .A2(new_n264), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n752), .A2(new_n301), .B1(new_n761), .B2(new_n987), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n758), .A2(new_n768), .B1(new_n750), .B2(new_n448), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n755), .A2(new_n410), .B1(new_n756), .B2(new_n486), .ZN(new_n1118));
  NOR4_X1   g0918(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G137), .A2(new_n1054), .B1(new_n766), .B2(G125), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT54), .B(G143), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n756), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n356), .B1(new_n985), .B2(G50), .ZN(new_n1123));
  INV_X1    g0923(.A(G128), .ZN(new_n1124));
  INV_X1    g0924(.A(G132), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1123), .B1(new_n1124), .B2(new_n758), .C1(new_n1125), .C2(new_n750), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1122), .B(new_n1126), .C1(G159), .C2(new_n747), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n739), .A2(new_n806), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1114), .A2(new_n1119), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1112), .B1(new_n1034), .B2(new_n1130), .C1(new_n912), .C2(new_n730), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n621), .A2(new_n622), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n299), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n858), .A2(G330), .A3(new_n447), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n919), .A4(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1097), .A2(new_n848), .A3(new_n850), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT115), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT115), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1097), .A2(new_n1138), .A3(new_n848), .A4(new_n850), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1137), .A2(new_n1079), .A3(new_n1077), .A4(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n714), .A2(G330), .A3(new_n824), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1141), .A2(new_n848), .A3(new_n850), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1102), .B1(new_n1098), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1135), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(KEYINPUT114), .B(new_n1076), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1098), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT114), .B1(new_n1147), .B2(new_n1076), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1093), .B(new_n1144), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT116), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1109), .A2(new_n1145), .A3(new_n1098), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1152), .A2(KEYINPUT116), .A3(new_n1093), .A4(new_n1144), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(KEYINPUT117), .A3(new_n1040), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1110), .B2(new_n1144), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT117), .B1(new_n1154), .B2(new_n1040), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1111), .B(new_n1131), .C1(new_n1156), .C2(new_n1157), .ZN(G378));
  NAND2_X1  g0958(.A1(new_n898), .A2(G330), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n298), .A2(new_n642), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n300), .B(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n914), .B2(new_n917), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n914), .A2(new_n917), .A3(new_n1163), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1159), .B(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1163), .A2(new_n729), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n729), .A2(G50), .A3(new_n782), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G125), .A2(new_n772), .B1(new_n797), .B2(G128), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G132), .A2(new_n1054), .B1(new_n800), .B2(G137), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n806), .B2(new_n746), .C1(new_n739), .C2(new_n1121), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n319), .B(new_n274), .C1(new_n752), .C2(new_n762), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G124), .B2(new_n766), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n772), .A2(G116), .B1(new_n766), .B2(G283), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n403), .B2(new_n756), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n278), .B(new_n356), .C1(new_n752), .C2(new_n349), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n486), .A2(new_n755), .B1(new_n750), .B2(new_n410), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n978), .C1(new_n264), .C2(new_n739), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT58), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n316), .C2(new_n262), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1180), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n722), .B(new_n1171), .C1(new_n1191), .C2(new_n782), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1169), .A2(new_n970), .B1(new_n1170), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT119), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1135), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1154), .B2(new_n1196), .ZN(new_n1197));
  AOI211_X1 g0997(.A(KEYINPUT119), .B(new_n1135), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1169), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT57), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT57), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1169), .B(new_n1201), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1194), .B1(new_n1203), .B2(new_n1040), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(G375));
  INV_X1    g1005(.A(new_n1144), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n952), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1140), .A2(new_n1143), .A3(new_n1135), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1095), .A2(new_n729), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n726), .B1(new_n817), .B2(G68), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n750), .A2(new_n803), .B1(new_n756), .B2(new_n806), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n758), .A2(new_n1125), .B1(new_n761), .B2(new_n1124), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n262), .B1(new_n752), .B2(new_n349), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n755), .A2(new_n1121), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n202), .B2(new_n746), .C1(new_n762), .C2(new_n739), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G116), .A2(new_n1054), .B1(new_n766), .B2(G303), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n410), .B2(new_n756), .C1(new_n987), .C2(new_n758), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n262), .B(new_n1220), .C1(G77), .C2(new_n985), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n486), .B2(new_n739), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1014), .B1(new_n768), .B2(new_n750), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT120), .Z(new_n1224));
  OAI21_X1  g1024(.A(new_n1218), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1212), .B1(new_n1225), .B2(new_n782), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1210), .A2(new_n970), .B1(new_n1211), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1209), .A2(new_n1227), .ZN(G381));
  AOI21_X1  g1028(.A(new_n667), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1229), .A2(G378), .A3(new_n1194), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1072), .A2(new_n971), .A3(new_n998), .ZN(new_n1231));
  OR2_X1    g1031(.A1(G393), .A2(G396), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1231), .A2(G384), .A3(G381), .A4(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(G407));
  INV_X1    g1034(.A(G378), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1204), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(G213), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n644), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT121), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1208), .B(KEYINPUT60), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT122), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1144), .A2(new_n667), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1227), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1245), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1243), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT122), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1252), .A2(G384), .A3(new_n1227), .A4(new_n1247), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT123), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT123), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1250), .A2(new_n1256), .A3(new_n1253), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1229), .A2(new_n1235), .A3(new_n1194), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT116), .B1(new_n1110), .B2(new_n1144), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1196), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT119), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1154), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n1207), .A3(new_n1169), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G378), .B1(new_n1267), .B2(new_n1193), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1239), .B(new_n1259), .C1(new_n1260), .C2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT62), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1201), .B1(new_n1266), .B2(new_n1169), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1202), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1040), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(G378), .A3(new_n1193), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1268), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1239), .A4(new_n1259), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT124), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1250), .A2(new_n1256), .A3(new_n1253), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1256), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1238), .A2(G2897), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1281), .A2(new_n1282), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1254), .A2(new_n1284), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1280), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(KEYINPUT124), .B(new_n1286), .C1(new_n1258), .C2(new_n1284), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1268), .B1(new_n1204), .B2(G378), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1291), .B2(new_n1238), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1270), .A2(new_n1271), .A3(new_n1279), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G390), .A2(G387), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(KEYINPUT125), .A3(new_n1231), .ZN(new_n1295));
  XOR2_X1   g1095(.A(G393), .B(G396), .Z(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1296), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1294), .A2(KEYINPUT125), .A3(new_n1231), .A4(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1293), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1297), .A2(new_n1271), .A3(new_n1299), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1303), .B(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1239), .A4(new_n1259), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1239), .B1(new_n1260), .B2(new_n1268), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1308), .B2(new_n1290), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1269), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1305), .B(new_n1306), .C1(new_n1309), .C2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1302), .A2(new_n1311), .ZN(G405));
  AOI21_X1  g1112(.A(new_n1235), .B1(new_n1274), .B2(new_n1193), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1250), .B(new_n1253), .C1(new_n1313), .C2(new_n1230), .ZN(new_n1314));
  OAI21_X1  g1114(.A(G378), .B1(new_n1229), .B2(new_n1194), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1236), .A2(new_n1258), .A3(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(new_n1316), .A3(new_n1300), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1300), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1318), .B2(KEYINPUT127), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT127), .ZN(new_n1320));
  AOI211_X1 g1120(.A(new_n1320), .B(new_n1300), .C1(new_n1314), .C2(new_n1316), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1319), .A2(new_n1321), .ZN(G402));
endmodule


