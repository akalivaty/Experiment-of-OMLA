

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777;

  OR2_X1 U378 ( .A1(n688), .A2(G902), .ZN(n468) );
  AND2_X2 U379 ( .A1(n426), .A2(n423), .ZN(n422) );
  AND2_X2 U380 ( .A1(n395), .A2(n394), .ZN(n396) );
  AND2_X4 U381 ( .A1(n388), .A2(n653), .ZN(n676) );
  AND2_X2 U382 ( .A1(n532), .A2(n721), .ZN(n552) );
  XNOR2_X2 U383 ( .A(n458), .B(G134), .ZN(n512) );
  XNOR2_X2 U384 ( .A(n585), .B(n446), .ZN(n670) );
  INV_X4 U385 ( .A(G953), .ZN(n483) );
  AND2_X1 U386 ( .A1(n555), .A2(n661), .ZN(n556) );
  NOR2_X1 U387 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U388 ( .A(n415), .B(KEYINPUT40), .ZN(n776) );
  NAND2_X1 U389 ( .A1(n422), .A2(n418), .ZN(n619) );
  AND2_X1 U390 ( .A1(n536), .A2(n725), .ZN(n401) );
  XNOR2_X1 U391 ( .A(n595), .B(n526), .ZN(n617) );
  XNOR2_X1 U392 ( .A(KEYINPUT15), .B(G902), .ZN(n650) );
  AND2_X1 U393 ( .A1(n532), .A2(n721), .ZN(n358) );
  XNOR2_X2 U394 ( .A(n525), .B(n524), .ZN(n532) );
  XNOR2_X1 U395 ( .A(n384), .B(n439), .ZN(n471) );
  XNOR2_X2 U396 ( .A(n764), .B(G146), .ZN(n382) );
  XNOR2_X2 U397 ( .A(n512), .B(n459), .ZN(n764) );
  XNOR2_X1 U398 ( .A(n630), .B(n436), .ZN(n410) );
  XNOR2_X1 U399 ( .A(n469), .B(G137), .ZN(n404) );
  NAND2_X1 U400 ( .A1(n410), .A2(KEYINPUT48), .ZN(n408) );
  NAND2_X1 U401 ( .A1(n405), .A2(n409), .ZN(n370) );
  NOR2_X1 U402 ( .A1(n631), .A2(KEYINPUT48), .ZN(n405) );
  INV_X1 U403 ( .A(n410), .ZN(n409) );
  NAND2_X1 U404 ( .A1(n407), .A2(n645), .ZN(n406) );
  XNOR2_X1 U405 ( .A(KEYINPUT4), .B(G131), .ZN(n459) );
  NOR2_X1 U406 ( .A1(n420), .A2(KEYINPUT83), .ZN(n419) );
  NOR2_X1 U407 ( .A1(n433), .A2(n425), .ZN(n424) );
  INV_X1 U408 ( .A(KEYINPUT83), .ZN(n425) );
  OR2_X1 U409 ( .A1(n670), .A2(n430), .ZN(n429) );
  NAND2_X1 U410 ( .A1(n650), .A2(n431), .ZN(n430) );
  INV_X1 U411 ( .A(n449), .ZN(n431) );
  INV_X1 U412 ( .A(G902), .ZN(n515) );
  OR2_X1 U413 ( .A1(n655), .A2(G902), .ZN(n400) );
  XNOR2_X1 U414 ( .A(G116), .B(G113), .ZN(n439) );
  XNOR2_X1 U415 ( .A(n440), .B(G119), .ZN(n384) );
  XNOR2_X1 U416 ( .A(G119), .B(KEYINPUT24), .ZN(n486) );
  XNOR2_X1 U417 ( .A(KEYINPUT87), .B(KEYINPUT23), .ZN(n485) );
  XNOR2_X1 U418 ( .A(G128), .B(G110), .ZN(n487) );
  XNOR2_X1 U419 ( .A(n374), .B(n371), .ZN(n664) );
  XNOR2_X1 U420 ( .A(n502), .B(n360), .ZN(n374) );
  XNOR2_X1 U421 ( .A(n373), .B(n372), .ZN(n371) );
  XNOR2_X1 U422 ( .A(G140), .B(G137), .ZN(n482) );
  XNOR2_X1 U423 ( .A(n416), .B(n435), .ZN(n633) );
  NOR2_X1 U424 ( .A1(n627), .A2(n628), .ZN(n416) );
  NAND2_X1 U425 ( .A1(n390), .A2(n389), .ZN(n388) );
  NOR2_X1 U426 ( .A1(n483), .A2(G952), .ZN(n691) );
  NAND2_X1 U427 ( .A1(n379), .A2(n569), .ZN(n378) );
  NAND2_X1 U428 ( .A1(n377), .A2(n375), .ZN(n631) );
  NAND2_X1 U429 ( .A1(n376), .A2(KEYINPUT47), .ZN(n375) );
  AND2_X1 U430 ( .A1(n363), .A2(n378), .ZN(n377) );
  NAND2_X1 U431 ( .A1(n613), .A2(n614), .ZN(n376) );
  INV_X1 U432 ( .A(G237), .ZN(n448) );
  NAND2_X1 U433 ( .A1(n393), .A2(n359), .ZN(n397) );
  XNOR2_X1 U434 ( .A(n501), .B(n498), .ZN(n373) );
  XOR2_X1 U435 ( .A(G140), .B(G104), .Z(n498) );
  XNOR2_X1 U436 ( .A(n499), .B(n497), .ZN(n372) );
  XNOR2_X1 U437 ( .A(G143), .B(G131), .ZN(n497) );
  XOR2_X1 U438 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n499) );
  NOR2_X1 U439 ( .A1(n406), .A2(n369), .ZN(n387) );
  NAND2_X1 U440 ( .A1(n370), .A2(n362), .ZN(n369) );
  NAND2_X1 U441 ( .A1(n447), .A2(n449), .ZN(n432) );
  XNOR2_X1 U442 ( .A(n563), .B(KEYINPUT1), .ZN(n536) );
  XNOR2_X1 U443 ( .A(n471), .B(n403), .ZN(n402) );
  XNOR2_X1 U444 ( .A(n404), .B(n470), .ZN(n403) );
  NOR2_X1 U445 ( .A1(n406), .A2(n368), .ZN(n770) );
  NAND2_X1 U446 ( .A1(n370), .A2(n408), .ZN(n368) );
  XNOR2_X1 U447 ( .A(G122), .B(KEYINPUT9), .ZN(n505) );
  XOR2_X1 U448 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n506) );
  XNOR2_X1 U449 ( .A(G116), .B(G107), .ZN(n508) );
  NAND2_X1 U450 ( .A1(n718), .A2(KEYINPUT77), .ZN(n389) );
  XNOR2_X1 U451 ( .A(G146), .B(G125), .ZN(n481) );
  XNOR2_X1 U452 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n443) );
  NAND2_X1 U453 ( .A1(n646), .A2(n770), .ZN(n718) );
  XNOR2_X1 U454 ( .A(n700), .B(n380), .ZN(n632) );
  INV_X1 U455 ( .A(KEYINPUT99), .ZN(n380) );
  NAND2_X1 U456 ( .A1(n421), .A2(n419), .ZN(n418) );
  NAND2_X1 U457 ( .A1(n428), .A2(KEYINPUT83), .ZN(n426) );
  AND2_X1 U458 ( .A1(n412), .A2(n411), .ZN(n626) );
  INV_X1 U459 ( .A(n601), .ZN(n411) );
  XNOR2_X1 U460 ( .A(n414), .B(n413), .ZN(n412) );
  INV_X1 U461 ( .A(KEYINPUT30), .ZN(n413) );
  XNOR2_X1 U462 ( .A(n503), .B(n504), .ZN(n559) );
  XNOR2_X1 U463 ( .A(n517), .B(n516), .ZN(n560) );
  BUF_X1 U464 ( .A(n536), .Z(n726) );
  XNOR2_X1 U465 ( .A(n462), .B(n438), .ZN(n385) );
  XNOR2_X1 U466 ( .A(KEYINPUT16), .B(G122), .ZN(n438) );
  XNOR2_X1 U467 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U468 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U469 ( .A(n382), .B(n464), .ZN(n688) );
  OR2_X1 U470 ( .A1(n633), .A2(n706), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n381), .B(KEYINPUT98), .ZN(n700) );
  OR2_X1 U472 ( .A1(n559), .A2(n560), .ZN(n381) );
  XNOR2_X1 U473 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U474 ( .A1(n676), .A2(G478), .ZN(n683) );
  AND2_X1 U475 ( .A1(n571), .A2(n361), .ZN(n359) );
  XOR2_X1 U476 ( .A(G113), .B(G122), .Z(n360) );
  XNOR2_X1 U477 ( .A(n562), .B(KEYINPUT100), .ZN(n742) );
  AND2_X1 U478 ( .A1(n570), .A2(n392), .ZN(n361) );
  AND2_X1 U479 ( .A1(n408), .A2(n417), .ZN(n362) );
  AND2_X1 U480 ( .A1(n622), .A2(n715), .ZN(n363) );
  AND2_X1 U481 ( .A1(n432), .A2(n737), .ZN(n364) );
  XNOR2_X1 U482 ( .A(n385), .B(n471), .ZN(n585) );
  AND2_X1 U483 ( .A1(n447), .A2(n647), .ZN(n365) );
  AND2_X1 U484 ( .A1(n557), .A2(KEYINPUT81), .ZN(n366) );
  NAND2_X1 U485 ( .A1(n650), .A2(n649), .ZN(n367) );
  NOR2_X2 U486 ( .A1(n658), .A2(n691), .ZN(n660) );
  NOR2_X2 U487 ( .A1(n667), .A2(n691), .ZN(n669) );
  NOR2_X2 U488 ( .A1(n674), .A2(n691), .ZN(n675) );
  OR2_X1 U489 ( .A1(n611), .A2(n612), .ZN(n379) );
  XNOR2_X1 U490 ( .A(n402), .B(n382), .ZN(n655) );
  XNOR2_X2 U491 ( .A(n383), .B(KEYINPUT45), .ZN(n646) );
  NAND2_X1 U492 ( .A1(n398), .A2(n578), .ZN(n383) );
  XNOR2_X2 U493 ( .A(n437), .B(G104), .ZN(n462) );
  NAND2_X1 U494 ( .A1(n386), .A2(n365), .ZN(n391) );
  NAND2_X1 U495 ( .A1(n646), .A2(n387), .ZN(n386) );
  NAND2_X1 U496 ( .A1(n391), .A2(n367), .ZN(n390) );
  NAND2_X1 U497 ( .A1(n571), .A2(n570), .ZN(n399) );
  INV_X1 U498 ( .A(KEYINPUT81), .ZN(n392) );
  NAND2_X1 U499 ( .A1(n558), .A2(n557), .ZN(n393) );
  NAND2_X1 U500 ( .A1(n399), .A2(KEYINPUT81), .ZN(n394) );
  NAND2_X1 U501 ( .A1(n558), .A2(n366), .ZN(n395) );
  NAND2_X1 U502 ( .A1(n397), .A2(n396), .ZN(n398) );
  INV_X1 U503 ( .A(n726), .ZN(n533) );
  NAND2_X1 U504 ( .A1(n401), .A2(n617), .ZN(n537) );
  XNOR2_X2 U505 ( .A(n400), .B(G472), .ZN(n595) );
  XNOR2_X2 U506 ( .A(n537), .B(KEYINPUT33), .ZN(n755) );
  NAND2_X1 U507 ( .A1(n631), .A2(KEYINPUT48), .ZN(n407) );
  NAND2_X1 U508 ( .A1(n595), .A2(n737), .ZN(n414) );
  INV_X1 U509 ( .A(KEYINPUT77), .ZN(n417) );
  INV_X1 U510 ( .A(n433), .ZN(n420) );
  INV_X1 U511 ( .A(n428), .ZN(n421) );
  INV_X1 U512 ( .A(n424), .ZN(n423) );
  NAND2_X1 U513 ( .A1(n427), .A2(n433), .ZN(n596) );
  AND2_X1 U514 ( .A1(n429), .A2(n432), .ZN(n427) );
  NAND2_X1 U515 ( .A1(n429), .A2(n364), .ZN(n428) );
  NAND2_X1 U516 ( .A1(n670), .A2(n449), .ZN(n433) );
  AND2_X1 U517 ( .A1(n572), .A2(n573), .ZN(n434) );
  XNOR2_X1 U518 ( .A(KEYINPUT70), .B(KEYINPUT39), .ZN(n435) );
  XOR2_X1 U519 ( .A(n629), .B(KEYINPUT64), .Z(n436) );
  XNOR2_X1 U520 ( .A(n619), .B(KEYINPUT19), .ZN(n609) );
  BUF_X1 U521 ( .A(n609), .Z(n705) );
  INV_X1 U522 ( .A(n681), .ZN(n682) );
  XNOR2_X1 U523 ( .A(G116), .B(KEYINPUT115), .ZN(n520) );
  XNOR2_X2 U524 ( .A(G110), .B(G107), .ZN(n437) );
  XNOR2_X2 U525 ( .A(G101), .B(KEYINPUT3), .ZN(n440) );
  XNOR2_X2 U526 ( .A(G128), .B(G143), .ZN(n458) );
  NAND2_X1 U527 ( .A1(n483), .A2(G224), .ZN(n441) );
  XNOR2_X1 U528 ( .A(n441), .B(KEYINPUT4), .ZN(n442) );
  XNOR2_X1 U529 ( .A(n458), .B(n442), .ZN(n445) );
  XNOR2_X1 U530 ( .A(n481), .B(n443), .ZN(n444) );
  XNOR2_X1 U531 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U532 ( .A(n650), .ZN(n447) );
  NAND2_X1 U533 ( .A1(n515), .A2(n448), .ZN(n450) );
  NAND2_X1 U534 ( .A1(n450), .A2(G210), .ZN(n449) );
  NAND2_X1 U535 ( .A1(n450), .A2(G214), .ZN(n737) );
  XNOR2_X1 U536 ( .A(G898), .B(KEYINPUT86), .ZN(n581) );
  NOR2_X1 U537 ( .A1(n483), .A2(n581), .ZN(n586) );
  NAND2_X1 U538 ( .A1(n586), .A2(G902), .ZN(n451) );
  NAND2_X1 U539 ( .A1(n483), .A2(G952), .ZN(n591) );
  NAND2_X1 U540 ( .A1(n451), .A2(n591), .ZN(n453) );
  NAND2_X1 U541 ( .A1(G237), .A2(G234), .ZN(n452) );
  XNOR2_X1 U542 ( .A(n452), .B(KEYINPUT14), .ZN(n719) );
  NAND2_X1 U543 ( .A1(n453), .A2(n719), .ZN(n454) );
  OR2_X2 U544 ( .A1(n609), .A2(n454), .ZN(n456) );
  INV_X1 U545 ( .A(KEYINPUT0), .ZN(n455) );
  XNOR2_X2 U546 ( .A(n456), .B(n455), .ZN(n538) );
  BUF_X1 U547 ( .A(n538), .Z(n457) );
  NAND2_X1 U548 ( .A1(n483), .A2(G227), .ZN(n460) );
  XNOR2_X1 U549 ( .A(n460), .B(G101), .ZN(n461) );
  XNOR2_X1 U550 ( .A(n461), .B(n482), .ZN(n463) );
  XOR2_X1 U551 ( .A(n463), .B(n462), .Z(n464) );
  XNOR2_X1 U552 ( .A(KEYINPUT67), .B(G469), .ZN(n466) );
  INV_X1 U553 ( .A(KEYINPUT66), .ZN(n465) );
  XNOR2_X1 U554 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X2 U555 ( .A(n468), .B(n467), .ZN(n563) );
  XOR2_X1 U556 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n470) );
  NOR2_X1 U557 ( .A1(G953), .A2(G237), .ZN(n500) );
  NAND2_X1 U558 ( .A1(G210), .A2(n500), .ZN(n469) );
  NAND2_X1 U559 ( .A1(n650), .A2(G234), .ZN(n472) );
  XNOR2_X1 U560 ( .A(n472), .B(KEYINPUT88), .ZN(n473) );
  XNOR2_X1 U561 ( .A(n473), .B(KEYINPUT20), .ZN(n476) );
  NAND2_X1 U562 ( .A1(n476), .A2(G221), .ZN(n475) );
  XNOR2_X1 U563 ( .A(KEYINPUT90), .B(KEYINPUT21), .ZN(n474) );
  XNOR2_X1 U564 ( .A(n475), .B(n474), .ZN(n720) );
  XNOR2_X1 U565 ( .A(n720), .B(KEYINPUT91), .ZN(n521) );
  NAND2_X1 U566 ( .A1(n476), .A2(G217), .ZN(n480) );
  XNOR2_X1 U567 ( .A(KEYINPUT73), .B(KEYINPUT89), .ZN(n478) );
  XNOR2_X1 U568 ( .A(KEYINPUT25), .B(KEYINPUT72), .ZN(n477) );
  XNOR2_X1 U569 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U570 ( .A(n480), .B(n479), .ZN(n494) );
  XNOR2_X1 U571 ( .A(n481), .B(KEYINPUT10), .ZN(n502) );
  XNOR2_X1 U572 ( .A(n502), .B(n482), .ZN(n763) );
  AND2_X1 U573 ( .A1(G234), .A2(n483), .ZN(n484) );
  XNOR2_X1 U574 ( .A(KEYINPUT8), .B(n484), .ZN(n510) );
  NAND2_X1 U575 ( .A1(n510), .A2(G221), .ZN(n491) );
  XNOR2_X1 U576 ( .A(n486), .B(n485), .ZN(n489) );
  XNOR2_X1 U577 ( .A(n487), .B(KEYINPUT68), .ZN(n488) );
  XNOR2_X1 U578 ( .A(n763), .B(n492), .ZN(n677) );
  AND2_X1 U579 ( .A1(n677), .A2(n515), .ZN(n493) );
  XNOR2_X1 U580 ( .A(n494), .B(n493), .ZN(n602) );
  AND2_X1 U581 ( .A1(n521), .A2(n602), .ZN(n725) );
  AND2_X1 U582 ( .A1(n595), .A2(n725), .ZN(n495) );
  AND2_X1 U583 ( .A1(n726), .A2(n495), .ZN(n731) );
  NAND2_X1 U584 ( .A1(n457), .A2(n731), .ZN(n496) );
  XNOR2_X1 U585 ( .A(n496), .B(KEYINPUT31), .ZN(n712) );
  XNOR2_X1 U586 ( .A(KEYINPUT13), .B(G475), .ZN(n504) );
  NAND2_X1 U587 ( .A1(G214), .A2(n500), .ZN(n501) );
  NOR2_X1 U588 ( .A1(G902), .A2(n664), .ZN(n503) );
  XNOR2_X1 U589 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U590 ( .A(n507), .B(KEYINPUT7), .Z(n509) );
  XNOR2_X1 U591 ( .A(n509), .B(n508), .ZN(n514) );
  NAND2_X1 U592 ( .A1(n510), .A2(G217), .ZN(n511) );
  XNOR2_X1 U593 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U594 ( .A(n514), .B(n513), .ZN(n681) );
  NAND2_X1 U595 ( .A1(n681), .A2(n515), .ZN(n517) );
  XOR2_X1 U596 ( .A(KEYINPUT96), .B(G478), .Z(n516) );
  INV_X1 U597 ( .A(n700), .ZN(n518) );
  NAND2_X1 U598 ( .A1(n712), .A2(n518), .ZN(n519) );
  XOR2_X1 U599 ( .A(n520), .B(n519), .Z(G18) );
  INV_X1 U600 ( .A(n559), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n560), .A2(n541), .ZN(n741) );
  INV_X1 U602 ( .A(n521), .ZN(n522) );
  NOR2_X1 U603 ( .A1(n741), .A2(n522), .ZN(n523) );
  NAND2_X1 U604 ( .A1(n538), .A2(n523), .ZN(n525) );
  XNOR2_X1 U605 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n524) );
  INV_X1 U606 ( .A(KEYINPUT6), .ZN(n526) );
  INV_X1 U607 ( .A(n617), .ZN(n527) );
  NAND2_X1 U608 ( .A1(n532), .A2(n527), .ZN(n528) );
  XNOR2_X1 U609 ( .A(n528), .B(KEYINPUT80), .ZN(n530) );
  INV_X1 U610 ( .A(n602), .ZN(n721) );
  OR2_X1 U611 ( .A1(n726), .A2(n721), .ZN(n529) );
  OR2_X1 U612 ( .A1(n530), .A2(n529), .ZN(n571) );
  XOR2_X1 U613 ( .A(G101), .B(KEYINPUT109), .Z(n531) );
  XNOR2_X1 U614 ( .A(n571), .B(n531), .ZN(G3) );
  NOR2_X1 U615 ( .A1(n617), .A2(n533), .ZN(n534) );
  NAND2_X1 U616 ( .A1(n358), .A2(n534), .ZN(n535) );
  XNOR2_X1 U617 ( .A(n535), .B(KEYINPUT32), .ZN(n574) );
  XNOR2_X1 U618 ( .A(n574), .B(G119), .ZN(G21) );
  NAND2_X1 U619 ( .A1(n538), .A2(n755), .ZN(n540) );
  INV_X1 U620 ( .A(KEYINPUT34), .ZN(n539) );
  XNOR2_X1 U621 ( .A(n540), .B(n539), .ZN(n543) );
  OR2_X1 U622 ( .A1(n560), .A2(n541), .ZN(n597) );
  INV_X1 U623 ( .A(n597), .ZN(n542) );
  NAND2_X1 U624 ( .A1(n543), .A2(n542), .ZN(n546) );
  INV_X1 U625 ( .A(KEYINPUT74), .ZN(n544) );
  XNOR2_X1 U626 ( .A(n544), .B(KEYINPUT35), .ZN(n545) );
  XNOR2_X2 U627 ( .A(n546), .B(n545), .ZN(n572) );
  INV_X1 U628 ( .A(n572), .ZN(n548) );
  INV_X1 U629 ( .A(KEYINPUT44), .ZN(n573) );
  NOR2_X1 U630 ( .A1(n573), .A2(KEYINPUT82), .ZN(n547) );
  NAND2_X1 U631 ( .A1(n548), .A2(n547), .ZN(n550) );
  NAND2_X1 U632 ( .A1(n572), .A2(KEYINPUT82), .ZN(n549) );
  NAND2_X1 U633 ( .A1(n550), .A2(n549), .ZN(n555) );
  INV_X1 U634 ( .A(n595), .ZN(n724) );
  AND2_X1 U635 ( .A1(n533), .A2(n724), .ZN(n551) );
  NAND2_X1 U636 ( .A1(n552), .A2(n551), .ZN(n554) );
  INV_X1 U637 ( .A(KEYINPUT101), .ZN(n553) );
  XNOR2_X2 U638 ( .A(n554), .B(n553), .ZN(n661) );
  NAND2_X1 U639 ( .A1(n556), .A2(n574), .ZN(n558) );
  NAND2_X1 U640 ( .A1(n573), .A2(KEYINPUT82), .ZN(n557) );
  NAND2_X1 U641 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U642 ( .A(n561), .B(KEYINPUT97), .ZN(n711) );
  INV_X1 U643 ( .A(n711), .ZN(n706) );
  AND2_X1 U644 ( .A1(n632), .A2(n706), .ZN(n562) );
  INV_X1 U645 ( .A(n742), .ZN(n569) );
  NAND2_X1 U646 ( .A1(n563), .A2(n725), .ZN(n565) );
  INV_X1 U647 ( .A(KEYINPUT92), .ZN(n564) );
  XNOR2_X1 U648 ( .A(n565), .B(n564), .ZN(n599) );
  AND2_X1 U649 ( .A1(n599), .A2(n724), .ZN(n566) );
  NAND2_X1 U650 ( .A1(n457), .A2(n566), .ZN(n695) );
  INV_X1 U651 ( .A(n695), .ZN(n567) );
  OR2_X1 U652 ( .A1(n712), .A2(n567), .ZN(n568) );
  NAND2_X1 U653 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U654 ( .A1(n661), .A2(n434), .ZN(n576) );
  INV_X1 U655 ( .A(n574), .ZN(n575) );
  XNOR2_X1 U656 ( .A(n577), .B(KEYINPUT69), .ZN(n578) );
  NAND2_X1 U657 ( .A1(n646), .A2(n483), .ZN(n584) );
  NAND2_X1 U658 ( .A1(G224), .A2(G953), .ZN(n579) );
  XNOR2_X1 U659 ( .A(n579), .B(KEYINPUT124), .ZN(n580) );
  XNOR2_X1 U660 ( .A(KEYINPUT61), .B(n580), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n589) );
  NOR2_X1 U663 ( .A1(n585), .A2(n586), .ZN(n587) );
  XOR2_X1 U664 ( .A(KEYINPUT125), .B(n587), .Z(n588) );
  XNOR2_X1 U665 ( .A(n589), .B(n588), .ZN(G69) );
  NOR2_X1 U666 ( .A1(G900), .A2(n483), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n590), .A2(G902), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n593), .A2(n719), .ZN(n594) );
  XOR2_X1 U670 ( .A(KEYINPUT75), .B(n594), .Z(n601) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n626), .A2(n598), .ZN(n600) );
  INV_X1 U673 ( .A(n599), .ZN(n628) );
  NOR2_X1 U674 ( .A1(n600), .A2(n628), .ZN(n616) );
  XOR2_X1 U675 ( .A(G143), .B(n616), .Z(G45) );
  INV_X1 U676 ( .A(KEYINPUT76), .ZN(n612) );
  XOR2_X1 U677 ( .A(KEYINPUT104), .B(KEYINPUT28), .Z(n605) );
  OR2_X1 U678 ( .A1(n720), .A2(n601), .ZN(n603) );
  OR2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n638) );
  OR2_X1 U680 ( .A1(n724), .A2(n638), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n605), .B(n604), .ZN(n607) );
  XOR2_X1 U682 ( .A(KEYINPUT103), .B(n563), .Z(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n608), .B(KEYINPUT105), .ZN(n708) );
  INV_X1 U685 ( .A(n705), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n708), .A2(n610), .ZN(n701) );
  NOR2_X1 U687 ( .A1(n701), .A2(KEYINPUT47), .ZN(n611) );
  INV_X1 U688 ( .A(n701), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n742), .A2(KEYINPUT76), .ZN(n613) );
  NOR2_X1 U690 ( .A1(KEYINPUT47), .A2(KEYINPUT76), .ZN(n615) );
  NOR2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n711), .A2(n617), .ZN(n635) );
  NOR2_X1 U693 ( .A1(n638), .A2(n635), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U695 ( .A(n620), .B(KEYINPUT36), .Z(n621) );
  NAND2_X1 U696 ( .A1(n621), .A2(n726), .ZN(n715) );
  XNOR2_X1 U697 ( .A(n596), .B(KEYINPUT38), .ZN(n738) );
  NAND2_X1 U698 ( .A1(n738), .A2(n737), .ZN(n743) );
  NOR2_X1 U699 ( .A1(n743), .A2(n741), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT41), .B(KEYINPUT106), .Z(n623) );
  XNOR2_X1 U701 ( .A(n624), .B(n623), .ZN(n756) );
  NAND2_X1 U702 ( .A1(n756), .A2(n708), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT42), .ZN(n777) );
  NAND2_X1 U704 ( .A1(n626), .A2(n738), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n777), .A2(n776), .ZN(n630) );
  XNOR2_X1 U706 ( .A(KEYINPUT46), .B(KEYINPUT79), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U708 ( .A(KEYINPUT107), .B(n634), .ZN(n774) );
  INV_X1 U709 ( .A(n635), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n737), .A2(n636), .ZN(n637) );
  NOR2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U712 ( .A1(n533), .A2(n639), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n640), .B(KEYINPUT43), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n641), .A2(n596), .ZN(n643) );
  INV_X1 U715 ( .A(KEYINPUT102), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n643), .B(n642), .ZN(n775) );
  INV_X1 U717 ( .A(n775), .ZN(n644) );
  AND2_X1 U718 ( .A1(n774), .A2(n644), .ZN(n645) );
  NAND2_X1 U719 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n647) );
  INV_X1 U720 ( .A(KEYINPUT2), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n651), .A2(KEYINPUT78), .ZN(n648) );
  NOR2_X1 U722 ( .A1(KEYINPUT77), .A2(n648), .ZN(n649) );
  NOR2_X1 U723 ( .A1(n718), .A2(n651), .ZN(n652) );
  INV_X1 U724 ( .A(n652), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n676), .A2(G472), .ZN(n657) );
  XNOR2_X1 U726 ( .A(KEYINPUT108), .B(KEYINPUT62), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U729 ( .A(KEYINPUT84), .B(KEYINPUT63), .Z(n659) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(G57) );
  XNOR2_X1 U731 ( .A(n661), .B(G110), .ZN(G12) );
  NAND2_X1 U732 ( .A1(n676), .A2(G475), .ZN(n666) );
  XNOR2_X1 U733 ( .A(KEYINPUT85), .B(KEYINPUT122), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n662), .B(KEYINPUT59), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U737 ( .A(KEYINPUT65), .B(KEYINPUT60), .Z(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(G60) );
  NAND2_X1 U739 ( .A1(n676), .A2(G210), .ZN(n673) );
  XOR2_X1 U740 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n671) );
  XNOR2_X1 U741 ( .A(n670), .B(n671), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n675), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U744 ( .A(n572), .B(G122), .ZN(G24) );
  NAND2_X1 U745 ( .A1(n676), .A2(G217), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT123), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n680), .A2(n691), .ZN(G66) );
  NOR2_X1 U749 ( .A1(n684), .A2(n691), .ZN(G63) );
  NAND2_X1 U750 ( .A1(n676), .A2(G469), .ZN(n690) );
  XOR2_X1 U751 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n686) );
  XNOR2_X1 U752 ( .A(KEYINPUT121), .B(KEYINPUT120), .ZN(n685) );
  XOR2_X1 U753 ( .A(n686), .B(n685), .Z(n687) );
  XNOR2_X1 U754 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U755 ( .A(n690), .B(n689), .ZN(n692) );
  NOR2_X1 U756 ( .A1(n692), .A2(n691), .ZN(G54) );
  NOR2_X1 U757 ( .A1(n706), .A2(n695), .ZN(n693) );
  XOR2_X1 U758 ( .A(KEYINPUT110), .B(n693), .Z(n694) );
  XNOR2_X1 U759 ( .A(G104), .B(n694), .ZN(G6) );
  NOR2_X1 U760 ( .A1(n695), .A2(n700), .ZN(n699) );
  XOR2_X1 U761 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n697) );
  XNOR2_X1 U762 ( .A(G107), .B(KEYINPUT26), .ZN(n696) );
  XNOR2_X1 U763 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U764 ( .A(n699), .B(n698), .ZN(G9) );
  NOR2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n703) );
  XNOR2_X1 U766 ( .A(KEYINPUT112), .B(KEYINPUT29), .ZN(n702) );
  XNOR2_X1 U767 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U768 ( .A(G128), .B(n704), .ZN(G30) );
  XOR2_X1 U769 ( .A(G146), .B(KEYINPUT113), .Z(n710) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U772 ( .A(n710), .B(n709), .ZN(G48) );
  NAND2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U774 ( .A(n713), .B(G113), .ZN(n714) );
  XNOR2_X1 U775 ( .A(KEYINPUT114), .B(n714), .ZN(G15) );
  XOR2_X1 U776 ( .A(KEYINPUT116), .B(n715), .Z(n716) );
  XNOR2_X1 U777 ( .A(n716), .B(KEYINPUT37), .ZN(n717) );
  XNOR2_X1 U778 ( .A(G125), .B(n717), .ZN(G27) );
  XNOR2_X1 U779 ( .A(n718), .B(KEYINPUT2), .ZN(n760) );
  INV_X1 U780 ( .A(n719), .ZN(n753) );
  INV_X1 U781 ( .A(n756), .ZN(n736) );
  NAND2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U783 ( .A(KEYINPUT49), .B(n722), .Z(n723) );
  NAND2_X1 U784 ( .A1(n724), .A2(n723), .ZN(n729) );
  NOR2_X1 U785 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U786 ( .A(n727), .B(KEYINPUT50), .ZN(n728) );
  NOR2_X1 U787 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U788 ( .A(n730), .B(KEYINPUT117), .ZN(n733) );
  INV_X1 U789 ( .A(n731), .ZN(n732) );
  NAND2_X1 U790 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U791 ( .A(KEYINPUT51), .B(n734), .ZN(n735) );
  NOR2_X1 U792 ( .A1(n736), .A2(n735), .ZN(n750) );
  NOR2_X1 U793 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U794 ( .A(n739), .B(KEYINPUT118), .ZN(n740) );
  NOR2_X1 U795 ( .A1(n741), .A2(n740), .ZN(n745) );
  NOR2_X1 U796 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U797 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U798 ( .A(KEYINPUT119), .B(n746), .Z(n748) );
  INV_X1 U799 ( .A(n755), .ZN(n747) );
  NOR2_X1 U800 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U801 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U802 ( .A(n751), .B(KEYINPUT52), .ZN(n752) );
  NOR2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U804 ( .A1(G952), .A2(n754), .ZN(n758) );
  NAND2_X1 U805 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U807 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U808 ( .A1(n483), .A2(n761), .ZN(n762) );
  XOR2_X1 U809 ( .A(KEYINPUT53), .B(n762), .Z(G75) );
  XNOR2_X1 U810 ( .A(n764), .B(n763), .ZN(n769) );
  XOR2_X1 U811 ( .A(G227), .B(n769), .Z(n765) );
  XNOR2_X1 U812 ( .A(n765), .B(KEYINPUT126), .ZN(n766) );
  NAND2_X1 U813 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U814 ( .A1(G953), .A2(n767), .ZN(n768) );
  XOR2_X1 U815 ( .A(KEYINPUT127), .B(n768), .Z(n773) );
  XNOR2_X1 U816 ( .A(n770), .B(n769), .ZN(n771) );
  NAND2_X1 U817 ( .A1(n771), .A2(n483), .ZN(n772) );
  NAND2_X1 U818 ( .A1(n773), .A2(n772), .ZN(G72) );
  XNOR2_X1 U819 ( .A(G134), .B(n774), .ZN(G36) );
  XOR2_X1 U820 ( .A(G140), .B(n775), .Z(G42) );
  XNOR2_X1 U821 ( .A(G131), .B(n776), .ZN(G33) );
  XNOR2_X1 U822 ( .A(G137), .B(n777), .ZN(G39) );
endmodule

