//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT67), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n209), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n218), .A2(G50), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n209), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n226), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n225), .B1(new_n231), .B2(KEYINPUT0), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n217), .B(new_n232), .C1(KEYINPUT0), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G116), .Z(new_n246));
  INV_X1    g0046(.A(G107), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G97), .ZN(new_n248));
  INV_X1    g0048(.A(G97), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G107), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n245), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G222), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n260), .B(new_n261), .C1(new_n202), .C2(new_n258), .ZN(new_n262));
  INV_X1    g0062(.A(new_n222), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(KEYINPUT69), .A2(G33), .A3(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n263), .A3(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n275), .A2(new_n269), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n271), .B1(new_n276), .B2(G226), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n267), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n222), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT70), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT70), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n283), .A3(new_n222), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n223), .A2(G1), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n223), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n223), .A2(new_n254), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n223), .B1(new_n201), .B2(new_n203), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n285), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n268), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G50), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n288), .A2(new_n295), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n279), .A2(G200), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(G190), .B2(new_n278), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n278), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n301), .C1(G169), .C2(new_n278), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n280), .A2(new_n283), .A3(new_n222), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n283), .B1(new_n280), .B2(new_n222), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n255), .A2(new_n257), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT7), .B1(new_n316), .B2(new_n223), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT7), .ZN(new_n318));
  AOI211_X1 g0118(.A(new_n318), .B(G20), .C1(new_n255), .C2(new_n257), .ZN(new_n319));
  OAI21_X1  g0119(.A(G68), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G58), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(G20), .B1(new_n323), .B2(new_n203), .ZN(new_n324));
  INV_X1    g0124(.A(new_n292), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G159), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT16), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n315), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT7), .A2(G20), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n254), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT75), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n256), .B2(G33), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n256), .A2(G33), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT76), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT75), .B1(new_n254), .B2(KEYINPUT3), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n255), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT76), .A3(new_n334), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n333), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(G20), .B1(new_n342), .B2(new_n334), .ZN(new_n345));
  OAI21_X1  g0145(.A(G68), .B1(new_n345), .B2(new_n318), .ZN(new_n346));
  OAI211_X1 g0146(.A(KEYINPUT16), .B(new_n328), .C1(new_n344), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n331), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n286), .A2(G13), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n289), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n287), .B2(new_n289), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(G226), .A2(G1698), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n334), .B(new_n353), .C1(new_n336), .C2(new_n337), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT77), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G87), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n342), .A2(G223), .A3(new_n259), .A4(new_n334), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n342), .A2(KEYINPUT77), .A3(new_n334), .A4(new_n353), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n356), .A2(new_n357), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n266), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n275), .A2(new_n269), .ZN(new_n362));
  INV_X1    g0162(.A(G232), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n362), .A2(new_n363), .B1(new_n270), .B2(new_n269), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(G179), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n364), .B1(new_n360), .B2(new_n266), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n352), .A2(new_n369), .A3(KEYINPUT18), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n352), .A2(new_n369), .A3(KEYINPUT78), .A4(KEYINPUT18), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n352), .A2(new_n369), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT18), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n368), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G200), .B2(new_n368), .ZN(new_n380));
  INV_X1    g0180(.A(new_n351), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n331), .B2(new_n347), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT17), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT17), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n380), .A2(new_n385), .A3(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n377), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT71), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n315), .B2(new_n349), .ZN(new_n391));
  NOR4_X1   g0191(.A1(new_n313), .A2(new_n298), .A3(new_n314), .A4(KEYINPUT71), .ZN(new_n392));
  OAI211_X1 g0192(.A(G68), .B(new_n296), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT73), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n223), .A2(G33), .A3(G77), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n322), .A2(G20), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n292), .A2(new_n299), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n394), .A3(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n285), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT11), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n298), .A2(new_n322), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT12), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n393), .A2(new_n404), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n271), .B1(new_n276), .B2(G238), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n316), .A2(new_n363), .A3(new_n259), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n255), .A2(new_n257), .A3(G226), .A4(new_n259), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G97), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n266), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT13), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n409), .A2(new_n417), .A3(new_n414), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(G179), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n367), .B1(new_n416), .B2(new_n418), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT14), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n409), .A2(new_n417), .A3(new_n414), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n417), .B1(new_n409), .B2(new_n414), .ZN(new_n424));
  OAI21_X1  g0224(.A(G169), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(KEYINPUT14), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n408), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT74), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n423), .A2(new_n424), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n408), .B1(G190), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(G200), .B1(new_n423), .B2(new_n424), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND4_X1   g0232(.A1(new_n393), .A2(new_n404), .A3(new_n406), .A4(new_n407), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n416), .A2(G190), .A3(new_n418), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(KEYINPUT74), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n427), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT72), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n247), .B2(new_n258), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n316), .A2(new_n363), .A3(G1698), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n266), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n271), .B1(new_n276), .B2(G244), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n439), .B1(new_n445), .B2(G179), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n443), .A2(KEYINPUT72), .A3(new_n308), .A4(new_n444), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n289), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(new_n325), .B1(G20), .B2(G77), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT15), .B(G87), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n290), .B2(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(new_n285), .B1(new_n202), .B2(new_n298), .ZN(new_n453));
  OAI211_X1 g0253(.A(G77), .B(new_n296), .C1(new_n391), .C2(new_n392), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n445), .A2(new_n367), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n454), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n445), .A2(G200), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n459), .C1(new_n378), .C2(new_n445), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n312), .A2(new_n389), .A3(new_n438), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT79), .ZN(new_n463));
  INV_X1    g0263(.A(G41), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(KEYINPUT79), .B2(G41), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(new_n275), .A3(G257), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n465), .A2(new_n467), .A3(new_n469), .A4(G274), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT80), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n471), .A2(KEYINPUT80), .A3(new_n472), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT4), .A2(G244), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n255), .A2(new_n257), .A3(new_n475), .A4(new_n259), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n255), .A2(new_n257), .A3(G250), .A4(G1698), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n342), .A2(G244), .A3(new_n259), .A4(new_n334), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n473), .A2(new_n474), .B1(new_n482), .B2(new_n265), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G200), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n471), .A2(new_n472), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(G190), .B(new_n486), .C1(new_n482), .C2(new_n265), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT81), .ZN(new_n488));
  OAI21_X1  g0288(.A(G107), .B1(new_n317), .B2(new_n319), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n247), .A2(KEYINPUT6), .A3(G97), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n251), .B2(KEYINPUT6), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G20), .B1(G77), .B2(new_n325), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n315), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n268), .A2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n282), .A2(new_n284), .A3(new_n349), .A4(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n249), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n349), .A2(G97), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n481), .A2(new_n480), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n266), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(G190), .A4(new_n486), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n484), .A2(new_n488), .A3(new_n498), .A4(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n496), .ZN(new_n506));
  INV_X1    g0306(.A(new_n497), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n489), .A2(new_n492), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n315), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n502), .B(new_n308), .C1(new_n473), .C2(new_n474), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n265), .B1(new_n499), .B2(new_n500), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n367), .B1(new_n511), .B2(new_n485), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n469), .A2(new_n226), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n275), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n469), .A2(G274), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n342), .A2(G238), .A3(new_n259), .A4(new_n334), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n342), .A2(G244), .A3(G1698), .A4(new_n334), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G116), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n518), .B1(new_n522), .B2(new_n266), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G190), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n342), .A2(new_n223), .A3(G68), .A4(new_n334), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT19), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n526), .A2(new_n223), .A3(G33), .A4(G97), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  INV_X1    g0328(.A(G87), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n529), .B1(new_n412), .B2(new_n223), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n285), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n298), .A2(new_n451), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n315), .A2(G87), .A3(new_n349), .A4(new_n494), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G200), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n524), .B(new_n536), .C1(new_n537), .C2(new_n523), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n315), .B1(new_n525), .B2(new_n531), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n495), .A2(new_n451), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  INV_X1    g0341(.A(new_n534), .ZN(new_n542));
  NOR4_X1   g0342(.A1(new_n539), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n532), .B2(new_n285), .ZN(new_n544));
  INV_X1    g0344(.A(new_n540), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT82), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n523), .A2(new_n308), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G169), .B2(new_n523), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n538), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT83), .B1(new_n514), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G116), .ZN(new_n552));
  AOI221_X4 g0352(.A(KEYINPUT84), .B1(new_n552), .B2(G20), .C1(new_n280), .C2(new_n222), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT84), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(G20), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n554), .B1(new_n281), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(G20), .B1(G33), .B2(G283), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n254), .A2(G97), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n553), .A2(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI221_X1 g0364(.A(KEYINPUT20), .B1(new_n560), .B2(new_n561), .C1(new_n553), .C2(new_n556), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n552), .B1(new_n268), .B2(G33), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n391), .B2(new_n392), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n298), .A2(new_n552), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n229), .A2(new_n259), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n230), .A2(G1698), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n342), .A2(new_n334), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n316), .A2(G303), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n265), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n470), .A2(new_n275), .ZN(new_n576));
  INV_X1    g0376(.A(G270), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n472), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n367), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n570), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(G190), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n564), .A2(new_n565), .B1(new_n552), .B2(new_n298), .ZN(new_n585));
  OAI21_X1  g0385(.A(G200), .B1(new_n575), .B2(new_n578), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n568), .A4(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(KEYINPUT21), .B(G169), .C1(new_n575), .C2(new_n578), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n573), .A2(new_n574), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n266), .ZN(new_n590));
  INV_X1    g0390(.A(new_n472), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n470), .A2(new_n275), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(G270), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n593), .A3(G179), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT86), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(new_n570), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n595), .B2(new_n570), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n583), .B(new_n587), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n544), .A2(new_n545), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n541), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n544), .A2(KEYINPUT82), .A3(new_n545), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n523), .A2(G169), .ZN(new_n605));
  AOI211_X1 g0405(.A(G179), .B(new_n518), .C1(new_n522), .C2(new_n266), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n522), .A2(new_n266), .ZN(new_n609));
  INV_X1    g0409(.A(new_n518), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n611), .B2(G200), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n604), .A2(new_n607), .B1(new_n612), .B2(new_n524), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n513), .A4(new_n505), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G250), .A2(G1698), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n229), .B2(G1698), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n342), .A2(new_n617), .A3(new_n334), .ZN(new_n618));
  INV_X1    g0418(.A(G294), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n254), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n265), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n470), .A2(new_n275), .A3(G264), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n308), .A3(new_n472), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n254), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n255), .B2(new_n341), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n620), .B1(new_n628), .B2(new_n617), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n472), .B(new_n623), .C1(new_n629), .C2(new_n265), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n367), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT87), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT22), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n529), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n342), .A2(new_n223), .A3(new_n334), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n223), .A2(G87), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n316), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n521), .A2(G20), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT23), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n223), .B2(G107), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n247), .A2(KEYINPUT23), .A3(G20), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n636), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT24), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n315), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n636), .A2(KEYINPUT24), .A3(new_n638), .A4(new_n643), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n495), .A2(new_n247), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT25), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n349), .B2(G107), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n298), .A2(KEYINPUT25), .A3(new_n247), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n632), .A2(new_n633), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n626), .A2(new_n631), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n649), .A2(new_n653), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n646), .B2(new_n647), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT87), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n622), .A2(new_n591), .A3(new_n624), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT88), .B1(new_n660), .B2(G200), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n378), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT88), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n630), .A2(new_n663), .A3(new_n537), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n655), .A2(new_n659), .B1(new_n658), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n551), .A2(new_n600), .A3(new_n615), .A4(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n462), .A2(new_n667), .ZN(G372));
  NAND3_X1  g0468(.A1(new_n430), .A2(new_n428), .A3(new_n431), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n435), .A2(KEYINPUT74), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n456), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n673), .A2(new_n427), .B1(new_n384), .B2(new_n386), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n368), .A2(new_n367), .ZN(new_n675));
  AOI211_X1 g0475(.A(new_n308), .B(new_n364), .C1(new_n360), .C2(new_n266), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT91), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n677), .A2(new_n678), .A3(new_n382), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT91), .B1(new_n352), .B2(new_n369), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n375), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n678), .B1(new_n677), .B2(new_n382), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n352), .A2(new_n369), .A3(KEYINPUT91), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(KEYINPUT18), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n307), .B1(new_n674), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n310), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n611), .A2(new_n367), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n689), .B(new_n548), .C1(new_n543), .C2(new_n546), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n513), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n613), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n691), .B1(new_n693), .B2(KEYINPUT26), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT26), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT89), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n690), .A2(new_n696), .A3(new_n538), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n690), .B2(new_n538), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n695), .B(new_n692), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n505), .A2(new_n513), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n664), .A2(new_n662), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n663), .B1(new_n630), .B2(new_n537), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n658), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n701), .B(new_n704), .C1(new_n697), .C2(new_n698), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n656), .A2(new_n658), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n595), .A2(new_n570), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n583), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n705), .A2(KEYINPUT90), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n550), .A2(KEYINPUT89), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n690), .A2(new_n696), .A3(new_n538), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT90), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(new_n701), .A4(new_n704), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n700), .B1(new_n711), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n688), .B1(new_n462), .B2(new_n717), .ZN(G369));
  NOR2_X1   g0518(.A1(new_n297), .A2(G20), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n268), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G213), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g0523(.A(KEYINPUT92), .B(G343), .Z(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n707), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT93), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n654), .A2(new_n726), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n666), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n706), .A2(new_n726), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n728), .B1(new_n666), .B2(new_n729), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n583), .B1(new_n597), .B2(new_n598), .ZN(new_n735));
  INV_X1    g0535(.A(new_n726), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT94), .Z(new_n738));
  AOI21_X1  g0538(.A(new_n727), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n736), .B1(new_n585), .B2(new_n568), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n709), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n599), .B2(new_n740), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n739), .A2(new_n745), .ZN(G399));
  INV_X1    g0546(.A(KEYINPUT95), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(new_n228), .B2(G41), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n227), .A2(KEYINPUT95), .A3(new_n464), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n528), .A2(new_n529), .A3(new_n552), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n751), .A2(new_n268), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n221), .B2(new_n751), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  AND2_X1   g0555(.A1(new_n694), .A2(new_n699), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n710), .A2(new_n707), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n704), .A2(new_n513), .A3(new_n505), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n712), .B2(new_n713), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n757), .B1(new_n759), .B2(new_n715), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n705), .A2(KEYINPUT90), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n756), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT29), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n762), .A2(new_n763), .A3(new_n736), .ZN(new_n764));
  OAI211_X1 g0564(.A(KEYINPUT26), .B(new_n692), .C1(new_n697), .C2(new_n698), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT97), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT97), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n714), .A2(new_n767), .A3(KEYINPUT26), .A4(new_n692), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n693), .A2(new_n695), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n633), .B1(new_n632), .B2(new_n654), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n656), .A2(new_n658), .A3(KEYINPUT87), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(new_n735), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n691), .B1(new_n774), .B2(new_n759), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n726), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n764), .B1(new_n763), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(G179), .B1(new_n590), .B2(new_n593), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n483), .A2(new_n779), .A3(new_n611), .A4(new_n630), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n511), .A2(new_n485), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n575), .A2(new_n578), .A3(new_n308), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n782), .A2(new_n523), .A3(new_n625), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n781), .B1(new_n785), .B2(KEYINPUT30), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT30), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n784), .A2(KEYINPUT96), .A3(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(KEYINPUT31), .B(new_n736), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT31), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n785), .A2(KEYINPUT30), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(new_n788), .A3(new_n780), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(new_n792), .B2(new_n726), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n667), .A2(new_n726), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G330), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n778), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n755), .B1(new_n797), .B2(G1), .ZN(G364));
  AOI21_X1  g0598(.A(new_n268), .B1(new_n719), .B2(G45), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n751), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n744), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G330), .B2(new_n742), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n222), .B1(G20), .B2(new_n367), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n223), .A2(G190), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT99), .Z(new_n807));
  NOR3_X1   g0607(.A1(new_n807), .A2(G179), .A3(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G159), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT32), .Z(new_n810));
  NOR2_X1   g0610(.A1(new_n223), .A2(new_n378), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n308), .A2(new_n537), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n308), .A2(G200), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n813), .A2(new_n299), .B1(new_n815), .B2(new_n321), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n806), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(G77), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT98), .Z(new_n820));
  NOR2_X1   g0620(.A1(G179), .A2(G200), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n223), .B1(new_n821), .B2(G190), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n249), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n537), .A2(G179), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n811), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n812), .A2(new_n806), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n258), .B1(new_n825), .B2(new_n529), .C1(new_n322), .C2(new_n826), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n807), .A2(G179), .A3(new_n537), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n823), .B(new_n827), .C1(new_n828), .C2(G107), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n810), .A2(new_n820), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n808), .A2(G329), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n316), .B1(new_n822), .B2(new_n619), .C1(new_n832), .C2(new_n817), .ZN(new_n833));
  INV_X1    g0633(.A(G303), .ZN(new_n834));
  INV_X1    g0634(.A(G322), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n834), .A2(new_n825), .B1(new_n815), .B2(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(KEYINPUT33), .B(G317), .Z(new_n837));
  INV_X1    g0637(.A(G326), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n826), .A2(new_n837), .B1(new_n813), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n833), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n828), .ZN(new_n841));
  INV_X1    g0641(.A(G283), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n831), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n805), .B1(new_n830), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n228), .A2(new_n316), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G355), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(G116), .B2(new_n227), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n220), .A2(G45), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n245), .B2(G45), .ZN(new_n849));
  INV_X1    g0649(.A(new_n343), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT76), .B1(new_n342), .B2(new_n334), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n228), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n847), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(G13), .A2(G33), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(G20), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n804), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n801), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n844), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n857), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n742), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n803), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G396));
  INV_X1    g0665(.A(new_n801), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n804), .A2(new_n855), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(new_n202), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n825), .ZN(new_n869));
  INV_X1    g0669(.A(new_n815), .ZN(new_n870));
  AOI22_X1  g0670(.A1(G107), .A2(new_n869), .B1(new_n870), .B2(G294), .ZN(new_n871));
  AOI22_X1  g0671(.A1(G87), .A2(new_n828), .B1(new_n808), .B2(G311), .ZN(new_n872));
  INV_X1    g0672(.A(new_n813), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G303), .A2(new_n873), .B1(new_n818), .B2(G116), .ZN(new_n874));
  INV_X1    g0674(.A(new_n826), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n258), .B(new_n823), .C1(G283), .C2(new_n875), .ZN(new_n876));
  AND4_X1   g0676(.A1(new_n871), .A2(new_n872), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n828), .A2(G68), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n808), .A2(G132), .ZN(new_n879));
  INV_X1    g0679(.A(new_n822), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(G58), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n869), .A2(G50), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n878), .A2(new_n879), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n852), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT100), .ZN(new_n886));
  AOI22_X1  g0686(.A1(G143), .A2(new_n870), .B1(new_n875), .B2(G150), .ZN(new_n887));
  AOI22_X1  g0687(.A1(G137), .A2(new_n873), .B1(new_n818), .B2(G159), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT34), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n877), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n460), .B1(new_n458), .B2(new_n736), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n456), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n672), .A2(new_n736), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI221_X1 g0696(.A(new_n868), .B1(new_n805), .B2(new_n891), .C1(new_n896), .C2(new_n856), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n717), .B2(new_n726), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n762), .A2(new_n736), .A3(new_n896), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(KEYINPUT101), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT101), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n895), .C1(new_n717), .C2(new_n726), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(new_n795), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n795), .B1(new_n900), .B2(new_n902), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n866), .B(new_n903), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI211_X1 g0706(.A(KEYINPUT102), .B(new_n795), .C1(new_n900), .C2(new_n902), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n897), .B1(new_n906), .B2(new_n907), .ZN(G384));
  OAI211_X1 g0708(.A(G116), .B(new_n224), .C1(new_n491), .C2(KEYINPUT35), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(KEYINPUT35), .B2(new_n491), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT36), .ZN(new_n911));
  OR3_X1    g0711(.A1(new_n220), .A2(new_n202), .A3(new_n323), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n201), .A2(G68), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n268), .B(G13), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  INV_X1    g0716(.A(new_n723), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT104), .B1(new_n352), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT104), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n382), .A2(new_n919), .A3(new_n723), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT37), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n383), .A2(new_n374), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n332), .B1(new_n850), .B2(new_n851), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n338), .A2(new_n223), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n322), .B1(new_n927), .B2(KEYINPUT7), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n327), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n925), .B(new_n285), .C1(new_n929), .C2(KEYINPUT16), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n347), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n328), .B1(new_n344), .B2(new_n346), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n330), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n925), .B1(new_n933), .B2(new_n285), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n351), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n917), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n369), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n937), .A3(new_n383), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n924), .B1(new_n938), .B2(KEYINPUT37), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n936), .B1(new_n377), .B2(new_n387), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n916), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n936), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n388), .A2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n935), .A2(new_n917), .B1(new_n382), .B2(new_n380), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n922), .B1(new_n944), .B2(new_n937), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n943), .B(KEYINPUT38), .C1(new_n945), .C2(new_n924), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n408), .A2(new_n726), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n437), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n671), .A2(new_n427), .A3(new_n948), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n895), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n794), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT106), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT40), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n794), .A2(new_n952), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n947), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n921), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n679), .A2(new_n680), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT105), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n380), .A2(new_n962), .A3(new_n382), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n383), .A2(KEYINPUT105), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n960), .A2(new_n961), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n924), .B1(new_n965), .B2(KEYINPUT37), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n681), .A2(new_n387), .A3(new_n684), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(new_n921), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n916), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n958), .B1(new_n969), .B2(new_n946), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n959), .B1(new_n970), .B2(new_n956), .ZN(new_n971));
  INV_X1    g0771(.A(new_n462), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n972), .A3(new_n794), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n947), .A2(new_n955), .A3(new_n958), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n964), .A2(new_n682), .A3(new_n683), .A4(new_n963), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT37), .B1(new_n975), .B2(new_n921), .ZN(new_n976));
  INV_X1    g0776(.A(new_n924), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n976), .A2(new_n977), .B1(new_n967), .B2(new_n921), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n946), .B1(KEYINPUT38), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n958), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n956), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(G330), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n462), .A2(new_n795), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n973), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n687), .B1(new_n777), .B2(new_n972), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n899), .A2(new_n894), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n950), .A2(new_n951), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(new_n947), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n685), .A2(new_n723), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n427), .A2(new_n726), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n947), .A2(KEYINPUT39), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT39), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n969), .A2(new_n996), .A3(new_n946), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n994), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n987), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n268), .B2(new_n719), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n987), .A2(new_n999), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n915), .B1(new_n1001), .B2(new_n1002), .ZN(G367));
  NOR2_X1   g0803(.A1(new_n536), .A2(new_n736), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n712), .B2(new_n713), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n691), .B2(new_n1004), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1006), .A2(new_n857), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(KEYINPUT108), .B(G137), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G77), .A2(new_n828), .B1(new_n808), .B2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G150), .A2(new_n870), .B1(new_n875), .B2(G159), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G143), .A2(new_n873), .B1(new_n869), .B2(G58), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n258), .B1(new_n817), .B2(new_n201), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G68), .B2(new_n880), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n828), .A2(G97), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n808), .A2(G317), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G294), .A2(new_n875), .B1(new_n818), .B2(G283), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G311), .A2(new_n873), .B1(new_n870), .B2(G303), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n869), .A2(G116), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT46), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1020), .A2(new_n1021), .B1(new_n880), .B2(G107), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n884), .B(new_n1022), .C1(new_n1021), .C2(new_n1020), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1014), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT47), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n805), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n853), .A2(new_n241), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1028), .B(new_n858), .C1(new_n227), .C2(new_n451), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n801), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1007), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n739), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n513), .A2(new_n736), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT107), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n701), .B1(new_n498), .B2(new_n736), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1033), .A2(KEYINPUT44), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT44), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n739), .B2(new_n1037), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n734), .A2(new_n738), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n727), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n1044), .A3(new_n1037), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT45), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n739), .A2(KEYINPUT45), .A3(new_n1037), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n745), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n732), .A2(new_n733), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n743), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n745), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(new_n738), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n795), .A3(new_n778), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1042), .A2(new_n1049), .A3(new_n745), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1051), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n797), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n750), .B(KEYINPUT41), .Z(new_n1061));
  AOI21_X1  g0861(.A(new_n800), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT43), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1006), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n734), .A2(new_n738), .A3(new_n1037), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(KEYINPUT42), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n655), .A2(new_n659), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n513), .B1(new_n1038), .B2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1065), .A2(KEYINPUT42), .B1(new_n1068), .B2(new_n736), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1064), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1006), .A2(new_n1063), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n745), .A2(new_n1038), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1072), .A2(new_n1075), .A3(new_n1073), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1032), .B1(new_n1062), .B2(new_n1079), .ZN(G387));
  INV_X1    g0880(.A(KEYINPUT112), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n797), .B2(new_n1055), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1055), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(KEYINPUT112), .A3(new_n796), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1082), .A2(new_n1084), .A3(new_n751), .A4(new_n1056), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n238), .A2(G45), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1086), .A2(new_n853), .B1(new_n752), .B2(new_n845), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT50), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n449), .B2(new_n299), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n289), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n468), .B1(new_n322), .B2(new_n202), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n752), .A4(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1087), .A2(new_n1092), .B1(G107), .B2(new_n227), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n866), .B1(new_n1093), .B2(new_n858), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT109), .B(G150), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n808), .A2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G50), .A2(new_n870), .B1(new_n869), .B2(G77), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n875), .A2(new_n449), .B1(new_n818), .B2(G68), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1015), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n822), .A2(new_n451), .ZN(new_n1100));
  INV_X1    g0900(.A(G159), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n813), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT110), .ZN(new_n1103));
  NOR4_X1   g0903(.A1(new_n1099), .A2(new_n884), .A3(new_n1100), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n813), .A2(new_n835), .B1(new_n826), .B2(new_n832), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT111), .ZN(new_n1106));
  INV_X1    g0906(.A(G317), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1106), .B1(new_n834), .B2(new_n817), .C1(new_n1107), .C2(new_n815), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT48), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n869), .A2(G294), .B1(new_n880), .B2(G283), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1111), .A2(KEYINPUT49), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n808), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n552), .A2(new_n841), .B1(new_n1113), .B2(new_n838), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1112), .A2(new_n852), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1111), .A2(KEYINPUT49), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1104), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1094), .B1(new_n1117), .B2(new_n805), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1052), .B2(new_n857), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n800), .B2(new_n1055), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1085), .A2(new_n1120), .ZN(G393));
  NAND3_X1  g0921(.A1(new_n1051), .A2(new_n800), .A3(new_n1058), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G150), .A2(new_n873), .B1(new_n870), .B2(G159), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(KEYINPUT51), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G87), .B2(new_n828), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n808), .A2(G143), .B1(new_n1123), .B2(KEYINPUT51), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n822), .A2(new_n202), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n322), .A2(new_n825), .B1(new_n826), .B2(new_n201), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n449), .C2(new_n818), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1125), .A2(new_n852), .A3(new_n1126), .A4(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G107), .A2(new_n828), .B1(new_n808), .B2(G322), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n316), .B1(new_n826), .B2(new_n834), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n825), .A2(new_n842), .B1(new_n817), .B2(new_n619), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(G116), .C2(new_n880), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n813), .A2(new_n1107), .B1(new_n815), .B2(new_n832), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT52), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n805), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n853), .A2(new_n252), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n859), .B1(new_n228), .B2(G97), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n866), .B(new_n1138), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1037), .B2(new_n862), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1059), .A2(new_n751), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1057), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1122), .B(new_n1142), .C1(new_n1143), .C2(new_n1144), .ZN(G390));
  INV_X1    g0945(.A(KEYINPUT115), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n993), .B1(new_n969), .B2(new_n946), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n894), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n776), .B2(new_n893), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n989), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n993), .B1(new_n988), .B2(new_n989), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n995), .A2(new_n997), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(G330), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n792), .A2(new_n726), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT31), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n792), .A2(new_n790), .A3(new_n726), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n704), .B1(new_n771), .B2(new_n772), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(new_n599), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1161), .A2(new_n551), .A3(new_n615), .A4(new_n736), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1155), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n952), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1154), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1151), .B(new_n1164), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n794), .A2(G330), .A3(new_n896), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1169), .A2(new_n1150), .B1(new_n1163), .B2(new_n952), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT114), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1149), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1150), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1164), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT114), .B1(new_n1174), .B2(new_n988), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1170), .A2(new_n1149), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1172), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n770), .A2(new_n775), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n763), .B1(new_n1178), .B2(new_n736), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n705), .A2(KEYINPUT90), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n716), .A3(new_n757), .ZN(new_n1181));
  AOI211_X1 g0981(.A(KEYINPUT29), .B(new_n726), .C1(new_n1181), .C2(new_n756), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n972), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n984), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n688), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT113), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT113), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n986), .A2(new_n1187), .A3(new_n1184), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1177), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n751), .B1(new_n1168), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n986), .B2(new_n1184), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n773), .A2(new_n735), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n690), .B1(new_n705), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n765), .A2(KEYINPUT97), .B1(new_n695), .B2(new_n693), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n1194), .B2(new_n768), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT29), .B1(new_n1195), .B2(new_n726), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n462), .B1(new_n1196), .B2(new_n764), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1197), .A2(KEYINPUT113), .A3(new_n687), .A4(new_n984), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1191), .A2(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1199), .A2(new_n1177), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1146), .B1(new_n1190), .B2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1199), .A2(new_n1166), .A3(new_n1167), .A4(new_n1177), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1168), .A2(new_n1189), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1202), .A2(new_n1203), .A3(KEYINPUT115), .A4(new_n751), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n995), .A2(new_n997), .A3(new_n855), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n826), .A2(new_n247), .B1(new_n817), .B2(new_n249), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n808), .A2(G294), .B1(KEYINPUT118), .B2(new_n1207), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n813), .A2(new_n842), .B1(new_n815), .B2(new_n552), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n316), .B1(new_n825), .B2(new_n529), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1127), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1207), .A2(KEYINPUT118), .ZN(new_n1212));
  AND4_X1   g1012(.A1(new_n878), .A2(new_n1208), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n841), .A2(new_n201), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n869), .A2(new_n1095), .ZN(new_n1215));
  XOR2_X1   g1015(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1216));
  XNOR2_X1  g1016(.A(new_n1215), .B(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n316), .B1(new_n870), .B2(G132), .ZN(new_n1218));
  INV_X1    g1018(.A(G128), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1217), .B(new_n1218), .C1(new_n1219), .C2(new_n813), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1214), .B(new_n1220), .C1(G125), .C2(new_n808), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n875), .A2(new_n1008), .ZN(new_n1222));
  XOR2_X1   g1022(.A(KEYINPUT54), .B(G143), .Z(new_n1223));
  NAND2_X1  g1023(.A1(new_n818), .A2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(new_n1101), .C2(new_n822), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT116), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1213), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(new_n805), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n866), .B(new_n1228), .C1(new_n289), .C2(new_n867), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1206), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1168), .B2(new_n799), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1205), .A2(new_n1232), .ZN(G378));
  OAI21_X1  g1033(.A(new_n1199), .B1(new_n1168), .B2(new_n1189), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n998), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n991), .A3(new_n990), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n311), .A2(new_n301), .A3(new_n917), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n301), .A2(new_n917), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n307), .A2(new_n310), .A3(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n939), .A2(new_n916), .A3(new_n940), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n976), .A2(new_n977), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n967), .A2(new_n921), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT38), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT40), .B1(new_n1248), .B2(new_n958), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1155), .B(new_n1243), .C1(new_n1249), .C2(new_n959), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1243), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n971), .B2(G330), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1236), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n982), .A2(new_n1243), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n971), .A2(G330), .A3(new_n1251), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n999), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1234), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT57), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT119), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT119), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n999), .ZN(new_n1264));
  OAI211_X1 g1064(.A(KEYINPUT57), .B(new_n1234), .C1(new_n1261), .C2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1260), .A2(new_n1265), .A3(new_n751), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1257), .A2(new_n800), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n866), .B1(new_n201), .B2(new_n867), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n825), .A2(new_n202), .B1(new_n817), .B2(new_n451), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G97), .A2(new_n875), .B1(new_n870), .B2(G107), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n552), .B2(new_n813), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1269), .B(new_n1271), .C1(G68), .C2(new_n880), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G58), .A2(new_n828), .B1(new_n808), .B2(G283), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n464), .A3(new_n884), .A4(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT58), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n873), .A2(G125), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(G128), .A2(new_n870), .B1(new_n875), .B2(G132), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n869), .A2(new_n1223), .B1(new_n818), .B2(G137), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n880), .A2(G150), .ZN(new_n1280));
  AND4_X1   g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT59), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n828), .A2(G159), .ZN(new_n1285));
  AOI211_X1 g1085(.A(G33), .B(G41), .C1(new_n808), .C2(G124), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(G50), .B1(new_n254), .B2(new_n464), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n852), .B2(G41), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1290));
  AND4_X1   g1090(.A1(new_n1276), .A2(new_n1287), .A3(new_n1289), .A4(new_n1290), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1268), .B1(new_n805), .B2(new_n1291), .C1(new_n1251), .C2(new_n856), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1267), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1266), .A2(new_n1293), .ZN(G375));
  AND3_X1   g1094(.A1(new_n1170), .A2(new_n1149), .A3(new_n1171), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1170), .A2(new_n1149), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n726), .B1(new_n1181), .B2(new_n756), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1148), .B1(new_n1297), .B2(new_n896), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1171), .B1(new_n1170), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1295), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1191), .B2(new_n1198), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n1061), .A3(new_n1189), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n866), .B1(new_n322), .B2(new_n867), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n321), .A2(new_n841), .B1(new_n1113), .B2(new_n1219), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n870), .A2(new_n1008), .ZN(new_n1305));
  OAI221_X1 g1105(.A(new_n1305), .B1(new_n291), .B2(new_n817), .C1(new_n1101), .C2(new_n825), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(G132), .A2(new_n873), .B1(new_n875), .B2(new_n1223), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n299), .B2(new_n822), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1304), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1309));
  OAI22_X1  g1109(.A1(new_n813), .A2(new_n619), .B1(new_n815), .B2(new_n842), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n825), .A2(new_n249), .B1(new_n817), .B2(new_n247), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n316), .B1(new_n826), .B2(new_n552), .ZN(new_n1312));
  NOR4_X1   g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .A4(new_n1100), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(G77), .A2(new_n828), .B1(new_n808), .B2(G303), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1309), .A2(new_n852), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1303), .B1(new_n805), .B2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(new_n1150), .B2(new_n855), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1177), .B2(new_n800), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1302), .A2(new_n1318), .ZN(G381));
  NOR2_X1   g1119(.A1(new_n1190), .A2(new_n1200), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1320), .A2(new_n1231), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1266), .A2(new_n1293), .A3(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1085), .A2(new_n864), .A3(new_n1120), .ZN(new_n1323));
  OR3_X1    g1123(.A1(G390), .A2(G384), .A3(new_n1323), .ZN(new_n1324));
  OR4_X1    g1124(.A1(G387), .A2(new_n1322), .A3(G381), .A4(new_n1324), .ZN(G407));
  OAI211_X1 g1125(.A(G407), .B(G213), .C1(new_n724), .C2(new_n1322), .ZN(G409));
  NAND2_X1  g1126(.A1(G393), .A2(G396), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1323), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT123), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1328), .B(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT124), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1122), .A2(new_n1142), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1042), .A2(new_n1049), .A3(new_n745), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1333), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1334), .A2(new_n750), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1144), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1332), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1061), .B1(new_n1334), .B2(new_n796), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1079), .B1(new_n1338), .B2(new_n799), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1331), .B(new_n1337), .C1(new_n1339), .C2(new_n1031), .ZN(new_n1340));
  OAI211_X1 g1140(.A(G390), .B(new_n1032), .C1(new_n1062), .C2(new_n1079), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1331), .B1(G387), .B2(new_n1337), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1330), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(G387), .A2(new_n1337), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1345), .A2(new_n1341), .A3(new_n1328), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n725), .A2(G213), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(G378), .A2(new_n1266), .A3(new_n1293), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n800), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1061), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1351), .B(new_n1292), .C1(new_n1352), .C2(new_n1258), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1321), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1349), .B1(new_n1350), .B2(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n750), .B1(new_n1199), .B2(new_n1177), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT60), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1301), .A2(new_n1357), .ZN(new_n1358));
  OAI211_X1 g1158(.A(new_n1300), .B(KEYINPUT60), .C1(new_n1191), .C2(new_n1198), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1356), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT120), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1361), .B(new_n897), .C1(new_n906), .C2(new_n907), .ZN(new_n1362));
  AND2_X1   g1162(.A1(new_n1362), .A2(new_n1318), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1360), .A2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(G384), .A2(KEYINPUT120), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1364), .A2(new_n1366), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1360), .A2(new_n1365), .A3(new_n1363), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(KEYINPUT63), .B1(new_n1355), .B2(new_n1369), .ZN(new_n1370));
  NOR3_X1   g1170(.A1(new_n1347), .A2(new_n1370), .A3(KEYINPUT61), .ZN(new_n1371));
  OR2_X1    g1171(.A1(new_n1355), .A2(KEYINPUT121), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1355), .A2(KEYINPUT121), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1349), .A2(G2897), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1374), .A2(KEYINPUT122), .ZN(new_n1375));
  OR2_X1    g1175(.A1(new_n1374), .A2(KEYINPUT122), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1360), .A2(new_n1365), .A3(new_n1363), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1365), .B1(new_n1360), .B2(new_n1363), .ZN(new_n1378));
  OAI211_X1 g1178(.A(new_n1375), .B(new_n1376), .C1(new_n1377), .C2(new_n1378), .ZN(new_n1379));
  NAND4_X1  g1179(.A1(new_n1367), .A2(KEYINPUT122), .A3(new_n1374), .A4(new_n1368), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1372), .A2(new_n1373), .A3(new_n1381), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1355), .A2(KEYINPUT63), .A3(new_n1369), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1371), .A2(new_n1382), .A3(new_n1383), .ZN(new_n1384));
  XNOR2_X1  g1184(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1385));
  AND2_X1   g1185(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1385), .B1(new_n1355), .B2(new_n1386), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1350), .A2(new_n1354), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1388), .A2(new_n1348), .A3(new_n1369), .ZN(new_n1389));
  INV_X1    g1189(.A(KEYINPUT62), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1389), .A2(new_n1390), .ZN(new_n1391));
  NAND3_X1  g1191(.A1(new_n1355), .A2(KEYINPUT62), .A3(new_n1369), .ZN(new_n1392));
  AOI21_X1  g1192(.A(new_n1387), .B1(new_n1391), .B2(new_n1392), .ZN(new_n1393));
  OAI21_X1  g1193(.A(new_n1347), .B1(new_n1393), .B2(KEYINPUT126), .ZN(new_n1394));
  INV_X1    g1194(.A(new_n1385), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1388), .A2(new_n1348), .ZN(new_n1396));
  AOI21_X1  g1196(.A(new_n1395), .B1(new_n1396), .B2(new_n1381), .ZN(new_n1397));
  INV_X1    g1197(.A(new_n1392), .ZN(new_n1398));
  AOI21_X1  g1198(.A(KEYINPUT62), .B1(new_n1355), .B2(new_n1369), .ZN(new_n1399));
  OAI211_X1 g1199(.A(new_n1397), .B(KEYINPUT126), .C1(new_n1398), .C2(new_n1399), .ZN(new_n1400));
  INV_X1    g1200(.A(new_n1400), .ZN(new_n1401));
  OAI21_X1  g1201(.A(new_n1384), .B1(new_n1394), .B2(new_n1401), .ZN(G405));
  INV_X1    g1202(.A(new_n1347), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(G375), .A2(new_n1321), .ZN(new_n1404));
  NAND2_X1  g1204(.A1(new_n1404), .A2(new_n1350), .ZN(new_n1405));
  OR2_X1    g1205(.A1(new_n1405), .A2(KEYINPUT127), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1406), .A2(new_n1369), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(new_n1405), .A2(KEYINPUT127), .ZN(new_n1408));
  AND2_X1   g1208(.A1(new_n1406), .A2(new_n1408), .ZN(new_n1409));
  OAI211_X1 g1209(.A(new_n1403), .B(new_n1407), .C1(new_n1409), .C2(new_n1369), .ZN(new_n1410));
  INV_X1    g1210(.A(new_n1407), .ZN(new_n1411));
  AOI21_X1  g1211(.A(new_n1369), .B1(new_n1406), .B2(new_n1408), .ZN(new_n1412));
  OAI21_X1  g1212(.A(new_n1347), .B1(new_n1411), .B2(new_n1412), .ZN(new_n1413));
  NAND2_X1  g1213(.A1(new_n1410), .A2(new_n1413), .ZN(G402));
endmodule


