

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U550 ( .A1(n710), .A2(n709), .ZN(n765) );
  BUF_X1 U551 ( .A(n602), .Z(n603) );
  BUF_X1 U552 ( .A(n604), .Z(n605) );
  XNOR2_X1 U553 ( .A(n723), .B(n722), .ZN(n755) );
  XOR2_X1 U554 ( .A(KEYINPUT17), .B(n518), .Z(n604) );
  XNOR2_X1 U555 ( .A(n515), .B(KEYINPUT64), .ZN(n516) );
  INV_X1 U556 ( .A(KEYINPUT23), .ZN(n515) );
  NOR2_X1 U557 ( .A1(n799), .A2(n798), .ZN(n513) );
  INV_X1 U558 ( .A(KEYINPUT26), .ZN(n730) );
  XNOR2_X1 U559 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n724) );
  XNOR2_X1 U560 ( .A(n725), .B(n724), .ZN(n727) );
  XNOR2_X1 U561 ( .A(n716), .B(KEYINPUT30), .ZN(n717) );
  XNOR2_X1 U562 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U563 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n722) );
  INV_X1 U564 ( .A(KEYINPUT100), .ZN(n756) );
  XNOR2_X1 U565 ( .A(n756), .B(KEYINPUT99), .ZN(n757) );
  XNOR2_X1 U566 ( .A(n773), .B(KEYINPUT32), .ZN(n774) );
  XNOR2_X1 U567 ( .A(n779), .B(n778), .ZN(n792) );
  OR2_X1 U568 ( .A1(n795), .A2(KEYINPUT33), .ZN(n802) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XNOR2_X1 U570 ( .A(n517), .B(n516), .ZN(n520) );
  INV_X1 U571 ( .A(G2105), .ZN(n514) );
  AND2_X1 U572 ( .A1(n514), .A2(G2104), .ZN(n602) );
  NAND2_X1 U573 ( .A1(G101), .A2(n602), .ZN(n517) );
  NAND2_X1 U574 ( .A1(G137), .A2(n604), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n520), .A2(n519), .ZN(n525) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n871) );
  NAND2_X1 U577 ( .A1(G113), .A2(n871), .ZN(n523) );
  INV_X1 U578 ( .A(G2105), .ZN(n521) );
  NOR2_X4 U579 ( .A1(G2104), .A2(n521), .ZN(n872) );
  NAND2_X1 U580 ( .A1(G125), .A2(n872), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X2 U582 ( .A1(n525), .A2(n524), .ZN(G160) );
  INV_X1 U583 ( .A(G651), .ZN(n532) );
  NOR2_X1 U584 ( .A1(G543), .A2(n532), .ZN(n526) );
  XOR2_X2 U585 ( .A(KEYINPUT1), .B(n526), .Z(n642) );
  NAND2_X1 U586 ( .A1(n642), .A2(G65), .ZN(n527) );
  XNOR2_X1 U587 ( .A(n527), .B(KEYINPUT68), .ZN(n530) );
  XNOR2_X1 U588 ( .A(G543), .B(KEYINPUT0), .ZN(n528) );
  XNOR2_X1 U589 ( .A(n528), .B(KEYINPUT65), .ZN(n627) );
  NOR2_X2 U590 ( .A1(G651), .A2(n627), .ZN(n649) );
  NAND2_X1 U591 ( .A1(G53), .A2(n649), .ZN(n529) );
  NAND2_X1 U592 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n531), .B(KEYINPUT69), .ZN(n537) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U595 ( .A1(G91), .A2(n643), .ZN(n534) );
  NOR2_X1 U596 ( .A1(n627), .A2(n532), .ZN(n639) );
  NAND2_X1 U597 ( .A1(G78), .A2(n639), .ZN(n533) );
  NAND2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(KEYINPUT67), .B(n535), .ZN(n536) );
  NAND2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X2 U601 ( .A(n538), .B(KEYINPUT70), .ZN(G299) );
  NAND2_X1 U602 ( .A1(G102), .A2(n602), .ZN(n540) );
  NAND2_X1 U603 ( .A1(G138), .A2(n604), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U605 ( .A1(G114), .A2(n871), .ZN(n542) );
  NAND2_X1 U606 ( .A1(G126), .A2(n872), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT85), .B(n543), .Z(n544) );
  NOR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(G164) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U611 ( .A1(G88), .A2(n643), .ZN(n547) );
  NAND2_X1 U612 ( .A1(G75), .A2(n639), .ZN(n546) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U614 ( .A1(G62), .A2(n642), .ZN(n549) );
  NAND2_X1 U615 ( .A1(G50), .A2(n649), .ZN(n548) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(G166) );
  NAND2_X1 U618 ( .A1(n643), .A2(G89), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G76), .A2(n639), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(KEYINPUT5), .ZN(n561) );
  XNOR2_X1 U623 ( .A(KEYINPUT73), .B(KEYINPUT6), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G63), .A2(n642), .ZN(n557) );
  NAND2_X1 U625 ( .A1(G51), .A2(n649), .ZN(n556) );
  NAND2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT7), .B(n562), .ZN(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n563), .B(KEYINPUT10), .ZN(n564) );
  XNOR2_X1 U633 ( .A(KEYINPUT72), .B(n564), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n826) );
  NAND2_X1 U635 ( .A1(n826), .A2(G567), .ZN(n565) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U637 ( .A1(G56), .A2(n642), .ZN(n566) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n566), .Z(n572) );
  NAND2_X1 U639 ( .A1(n643), .A2(G81), .ZN(n567) );
  XNOR2_X1 U640 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U641 ( .A1(G68), .A2(n639), .ZN(n568) );
  NAND2_X1 U642 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U643 ( .A(KEYINPUT13), .B(n570), .Z(n571) );
  NOR2_X1 U644 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n649), .A2(G43), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n1007) );
  INV_X1 U647 ( .A(G860), .ZN(n594) );
  OR2_X1 U648 ( .A1(n1007), .A2(n594), .ZN(G153) );
  NAND2_X1 U649 ( .A1(G52), .A2(n649), .ZN(n575) );
  XOR2_X1 U650 ( .A(KEYINPUT66), .B(n575), .Z(n580) );
  NAND2_X1 U651 ( .A1(G90), .A2(n643), .ZN(n577) );
  NAND2_X1 U652 ( .A1(G77), .A2(n639), .ZN(n576) );
  NAND2_X1 U653 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U654 ( .A(KEYINPUT9), .B(n578), .Z(n579) );
  NOR2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n642), .A2(G64), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n582), .A2(n581), .ZN(G301) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G66), .A2(n642), .ZN(n584) );
  NAND2_X1 U660 ( .A1(G92), .A2(n643), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U662 ( .A1(G79), .A2(n639), .ZN(n586) );
  NAND2_X1 U663 ( .A1(G54), .A2(n649), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U665 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U666 ( .A(KEYINPUT15), .B(n589), .Z(n1008) );
  OR2_X1 U667 ( .A1(n1008), .A2(G868), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(G284) );
  NOR2_X1 U669 ( .A1(G299), .A2(G868), .ZN(n593) );
  INV_X1 U670 ( .A(G868), .ZN(n659) );
  NOR2_X1 U671 ( .A1(G286), .A2(n659), .ZN(n592) );
  NOR2_X1 U672 ( .A1(n593), .A2(n592), .ZN(G297) );
  NAND2_X1 U673 ( .A1(n594), .A2(G559), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n595), .A2(n1008), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U676 ( .A1(n1008), .A2(G868), .ZN(n597) );
  NOR2_X1 U677 ( .A1(G559), .A2(n597), .ZN(n598) );
  XNOR2_X1 U678 ( .A(n598), .B(KEYINPUT74), .ZN(n600) );
  NOR2_X1 U679 ( .A1(n1007), .A2(G868), .ZN(n599) );
  NOR2_X1 U680 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G123), .A2(n872), .ZN(n601) );
  XNOR2_X1 U682 ( .A(n601), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G99), .A2(n603), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G135), .A2(n605), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G111), .A2(n871), .ZN(n608) );
  XNOR2_X1 U687 ( .A(KEYINPUT75), .B(n608), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U690 ( .A(KEYINPUT76), .B(n613), .ZN(n914) );
  XOR2_X1 U691 ( .A(n914), .B(G2096), .Z(n615) );
  XNOR2_X1 U692 ( .A(G2100), .B(KEYINPUT77), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G559), .A2(n1008), .ZN(n616) );
  XOR2_X1 U695 ( .A(n1007), .B(n616), .Z(n657) );
  XOR2_X1 U696 ( .A(n657), .B(KEYINPUT78), .Z(n617) );
  NOR2_X1 U697 ( .A1(G860), .A2(n617), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G67), .A2(n642), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G80), .A2(n639), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U701 ( .A1(G93), .A2(n643), .ZN(n620) );
  XNOR2_X1 U702 ( .A(KEYINPUT79), .B(n620), .ZN(n621) );
  NOR2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n649), .A2(G55), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n660) );
  XOR2_X1 U706 ( .A(n625), .B(n660), .Z(G145) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n626), .B(KEYINPUT80), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G49), .A2(n649), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G87), .A2(n627), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U712 ( .A1(n642), .A2(n630), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(G288) );
  AND2_X1 U714 ( .A1(n642), .A2(G60), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G85), .A2(n643), .ZN(n634) );
  NAND2_X1 U716 ( .A1(G72), .A2(n639), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n649), .A2(G47), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(G290) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n641) );
  NAND2_X1 U722 ( .A1(G73), .A2(n639), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n641), .B(n640), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G61), .A2(n642), .ZN(n645) );
  NAND2_X1 U725 ( .A1(G86), .A2(n643), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U727 ( .A(KEYINPUT81), .B(n646), .Z(n647) );
  NOR2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n649), .A2(G48), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(G305) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(G288), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n652), .B(n660), .ZN(n653) );
  XNOR2_X1 U733 ( .A(G299), .B(n653), .ZN(n655) );
  XNOR2_X1 U734 ( .A(G290), .B(G166), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(G305), .ZN(n892) );
  XOR2_X1 U737 ( .A(n892), .B(n657), .Z(n658) );
  NOR2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n662) );
  NOR2_X1 U739 ( .A1(G868), .A2(n660), .ZN(n661) );
  NOR2_X1 U740 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XNOR2_X1 U742 ( .A(n663), .B(KEYINPUT83), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n664), .B(KEYINPUT20), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U748 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  NAND2_X1 U749 ( .A1(G132), .A2(G82), .ZN(n668) );
  XNOR2_X1 U750 ( .A(n668), .B(KEYINPUT84), .ZN(n669) );
  XNOR2_X1 U751 ( .A(n669), .B(KEYINPUT22), .ZN(n670) );
  NOR2_X1 U752 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U753 ( .A1(G96), .A2(n671), .ZN(n831) );
  NAND2_X1 U754 ( .A1(n831), .A2(G2106), .ZN(n675) );
  NAND2_X1 U755 ( .A1(G108), .A2(G120), .ZN(n672) );
  NOR2_X1 U756 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U757 ( .A1(G69), .A2(n673), .ZN(n830) );
  NAND2_X1 U758 ( .A1(G567), .A2(n830), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n675), .A2(n674), .ZN(n832) );
  NAND2_X1 U760 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U761 ( .A1(n832), .A2(n676), .ZN(n829) );
  NAND2_X1 U762 ( .A1(n829), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  NAND2_X1 U764 ( .A1(n872), .A2(G119), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G95), .A2(n603), .ZN(n677) );
  XOR2_X1 U766 ( .A(KEYINPUT89), .B(n677), .Z(n678) );
  NAND2_X1 U767 ( .A1(n679), .A2(n678), .ZN(n683) );
  NAND2_X1 U768 ( .A1(G131), .A2(n605), .ZN(n681) );
  NAND2_X1 U769 ( .A1(G107), .A2(n871), .ZN(n680) );
  NAND2_X1 U770 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U771 ( .A1(n683), .A2(n682), .ZN(n881) );
  INV_X1 U772 ( .A(G1991), .ZN(n966) );
  NOR2_X1 U773 ( .A1(n881), .A2(n966), .ZN(n694) );
  NAND2_X1 U774 ( .A1(G105), .A2(n603), .ZN(n684) );
  XNOR2_X1 U775 ( .A(n684), .B(KEYINPUT38), .ZN(n689) );
  NAND2_X1 U776 ( .A1(G117), .A2(n871), .ZN(n686) );
  NAND2_X1 U777 ( .A1(G129), .A2(n872), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U779 ( .A(KEYINPUT90), .B(n687), .Z(n688) );
  NAND2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U781 ( .A1(G141), .A2(n605), .ZN(n690) );
  XNOR2_X1 U782 ( .A(KEYINPUT91), .B(n690), .ZN(n691) );
  NOR2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n885) );
  INV_X1 U784 ( .A(G1996), .ZN(n968) );
  NOR2_X1 U785 ( .A1(n885), .A2(n968), .ZN(n693) );
  OR2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n912) );
  NAND2_X1 U787 ( .A1(G40), .A2(G160), .ZN(n695) );
  XNOR2_X1 U788 ( .A(n695), .B(KEYINPUT86), .ZN(n708) );
  NOR2_X1 U789 ( .A1(G164), .A2(G1384), .ZN(n709) );
  NOR2_X1 U790 ( .A1(n708), .A2(n709), .ZN(n821) );
  AND2_X1 U791 ( .A1(n912), .A2(n821), .ZN(n812) );
  XOR2_X1 U792 ( .A(KEYINPUT92), .B(n812), .Z(n707) );
  XNOR2_X1 U793 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  NAND2_X1 U794 ( .A1(G104), .A2(n603), .ZN(n697) );
  NAND2_X1 U795 ( .A1(G140), .A2(n605), .ZN(n696) );
  NAND2_X1 U796 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U797 ( .A(n698), .B(KEYINPUT34), .ZN(n699) );
  XNOR2_X1 U798 ( .A(n699), .B(KEYINPUT87), .ZN(n705) );
  XNOR2_X1 U799 ( .A(KEYINPUT35), .B(KEYINPUT88), .ZN(n703) );
  NAND2_X1 U800 ( .A1(G116), .A2(n871), .ZN(n701) );
  NAND2_X1 U801 ( .A1(G128), .A2(n872), .ZN(n700) );
  NAND2_X1 U802 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U803 ( .A(n703), .B(n702), .ZN(n704) );
  NAND2_X1 U804 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U805 ( .A(KEYINPUT36), .B(n706), .Z(n886) );
  NOR2_X1 U806 ( .A1(n818), .A2(n886), .ZN(n913) );
  NAND2_X1 U807 ( .A1(n821), .A2(n913), .ZN(n816) );
  NAND2_X1 U808 ( .A1(n707), .A2(n816), .ZN(n807) );
  INV_X1 U809 ( .A(n708), .ZN(n710) );
  NOR2_X1 U810 ( .A1(G2084), .A2(n765), .ZN(n714) );
  NAND2_X1 U811 ( .A1(n714), .A2(G8), .ZN(n761) );
  NAND2_X1 U812 ( .A1(G8), .A2(n765), .ZN(n799) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n799), .ZN(n759) );
  XOR2_X1 U814 ( .A(G2078), .B(KEYINPUT25), .Z(n969) );
  NOR2_X1 U815 ( .A1(n969), .A2(n765), .ZN(n711) );
  XOR2_X1 U816 ( .A(KEYINPUT93), .B(n711), .Z(n713) );
  INV_X1 U817 ( .A(n765), .ZN(n736) );
  NOR2_X1 U818 ( .A1(n736), .A2(G1961), .ZN(n712) );
  NOR2_X1 U819 ( .A1(n713), .A2(n712), .ZN(n751) );
  AND2_X1 U820 ( .A1(G301), .A2(n751), .ZN(n721) );
  NOR2_X1 U821 ( .A1(n759), .A2(n714), .ZN(n715) );
  NAND2_X1 U822 ( .A1(G8), .A2(n715), .ZN(n718) );
  INV_X1 U823 ( .A(KEYINPUT97), .ZN(n716) );
  NOR2_X1 U824 ( .A1(G168), .A2(n719), .ZN(n720) );
  NOR2_X1 U825 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U826 ( .A1(G2072), .A2(n736), .ZN(n725) );
  INV_X1 U827 ( .A(G1956), .ZN(n944) );
  NOR2_X1 U828 ( .A1(n944), .A2(n736), .ZN(n726) );
  NOR2_X1 U829 ( .A1(n727), .A2(n726), .ZN(n745) );
  INV_X1 U830 ( .A(G299), .ZN(n744) );
  NOR2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n729) );
  XNOR2_X1 U832 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n728) );
  XNOR2_X1 U833 ( .A(n729), .B(n728), .ZN(n749) );
  NOR2_X1 U834 ( .A1(n765), .A2(n968), .ZN(n731) );
  XNOR2_X1 U835 ( .A(n731), .B(n730), .ZN(n733) );
  NAND2_X1 U836 ( .A1(n765), .A2(G1341), .ZN(n732) );
  NAND2_X1 U837 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U838 ( .A1(n1007), .A2(n734), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n1008), .A2(n741), .ZN(n740) );
  NAND2_X1 U840 ( .A1(n765), .A2(G1348), .ZN(n735) );
  XNOR2_X1 U841 ( .A(n735), .B(KEYINPUT96), .ZN(n738) );
  NAND2_X1 U842 ( .A1(n736), .A2(G2067), .ZN(n737) );
  NAND2_X1 U843 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U844 ( .A1(n740), .A2(n739), .ZN(n743) );
  OR2_X1 U845 ( .A1(n1008), .A2(n741), .ZN(n742) );
  NAND2_X1 U846 ( .A1(n743), .A2(n742), .ZN(n747) );
  NAND2_X1 U847 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U848 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U849 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U850 ( .A(n750), .B(KEYINPUT29), .ZN(n753) );
  NOR2_X1 U851 ( .A1(G301), .A2(n751), .ZN(n752) );
  NOR2_X1 U852 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X2 U853 ( .A1(n755), .A2(n754), .ZN(n762) );
  XNOR2_X1 U854 ( .A(n762), .B(n757), .ZN(n758) );
  NOR2_X1 U855 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U856 ( .A1(n761), .A2(n760), .ZN(n777) );
  XNOR2_X1 U857 ( .A(n762), .B(KEYINPUT99), .ZN(n764) );
  AND2_X1 U858 ( .A1(G286), .A2(G8), .ZN(n763) );
  NAND2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n772) );
  INV_X1 U860 ( .A(G8), .ZN(n770) );
  NOR2_X1 U861 ( .A1(G1971), .A2(n799), .ZN(n767) );
  NOR2_X1 U862 ( .A1(G2090), .A2(n765), .ZN(n766) );
  NOR2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U864 ( .A1(n768), .A2(G303), .ZN(n769) );
  OR2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U866 ( .A1(n772), .A2(n771), .ZN(n775) );
  XNOR2_X1 U867 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n773) );
  XNOR2_X1 U868 ( .A(n775), .B(n774), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n779) );
  INV_X1 U870 ( .A(KEYINPUT103), .ZN(n778) );
  INV_X1 U871 ( .A(n792), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G166), .A2(G8), .ZN(n780) );
  NOR2_X1 U873 ( .A1(G2090), .A2(n780), .ZN(n781) );
  NOR2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U875 ( .A(KEYINPUT106), .B(n783), .ZN(n784) );
  INV_X1 U876 ( .A(n799), .ZN(n788) );
  NOR2_X1 U877 ( .A1(n784), .A2(n788), .ZN(n785) );
  XNOR2_X1 U878 ( .A(n785), .B(KEYINPUT107), .ZN(n790) );
  NOR2_X1 U879 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XNOR2_X1 U880 ( .A(n786), .B(KEYINPUT24), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n805) );
  NAND2_X1 U883 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  NOR2_X1 U884 ( .A1(G1976), .A2(G288), .ZN(n797) );
  NOR2_X1 U885 ( .A1(G1971), .A2(G303), .ZN(n791) );
  NOR2_X1 U886 ( .A1(n797), .A2(n791), .ZN(n1004) );
  NAND2_X1 U887 ( .A1(n792), .A2(n1004), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n1000), .A2(n793), .ZN(n794) );
  NOR2_X1 U889 ( .A1(n799), .A2(n794), .ZN(n795) );
  XOR2_X1 U890 ( .A(G1981), .B(KEYINPUT104), .Z(n796) );
  XNOR2_X1 U891 ( .A(G305), .B(n796), .ZN(n994) );
  INV_X1 U892 ( .A(n994), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n797), .A2(KEYINPUT33), .ZN(n798) );
  NOR2_X1 U894 ( .A1(n800), .A2(n513), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U896 ( .A(n803), .B(KEYINPUT105), .ZN(n804) );
  NOR2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U898 ( .A1(n807), .A2(n806), .ZN(n809) );
  XNOR2_X1 U899 ( .A(G1986), .B(G290), .ZN(n1006) );
  NAND2_X1 U900 ( .A1(n1006), .A2(n821), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n824) );
  AND2_X1 U902 ( .A1(n966), .A2(n881), .ZN(n916) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n916), .A2(n810), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n814) );
  AND2_X1 U906 ( .A1(n885), .A2(n968), .ZN(n813) );
  XNOR2_X1 U907 ( .A(n813), .B(KEYINPUT108), .ZN(n922) );
  NOR2_X1 U908 ( .A1(n814), .A2(n922), .ZN(n815) );
  XNOR2_X1 U909 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U911 ( .A1(n818), .A2(n886), .ZN(n924) );
  NAND2_X1 U912 ( .A1(n819), .A2(n924), .ZN(n820) );
  XOR2_X1 U913 ( .A(KEYINPUT109), .B(n820), .Z(n822) );
  NAND2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U916 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U917 ( .A(G301), .ZN(G171) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U920 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(G188) );
  NOR2_X1 U923 ( .A1(n831), .A2(n830), .ZN(G325) );
  XNOR2_X1 U924 ( .A(KEYINPUT111), .B(G325), .ZN(G261) );
  INV_X1 U925 ( .A(n832), .ZN(G319) );
  XNOR2_X1 U926 ( .A(G1986), .B(G2474), .ZN(n842) );
  XOR2_X1 U927 ( .A(G1976), .B(G1956), .Z(n834) );
  XNOR2_X1 U928 ( .A(G1971), .B(G1961), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U930 ( .A(G1966), .B(G1981), .Z(n836) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U933 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U934 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n844) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2072), .Z(n846) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2090), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U943 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U944 ( .A(G2084), .B(G2078), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(G227) );
  NAND2_X1 U946 ( .A1(G100), .A2(n603), .ZN(n852) );
  NAND2_X1 U947 ( .A1(G112), .A2(n871), .ZN(n851) );
  NAND2_X1 U948 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U949 ( .A(n853), .B(KEYINPUT113), .ZN(n855) );
  NAND2_X1 U950 ( .A1(G136), .A2(n605), .ZN(n854) );
  NAND2_X1 U951 ( .A1(n855), .A2(n854), .ZN(n858) );
  NAND2_X1 U952 ( .A1(n872), .A2(G124), .ZN(n856) );
  XOR2_X1 U953 ( .A(KEYINPUT44), .B(n856), .Z(n857) );
  NOR2_X1 U954 ( .A1(n858), .A2(n857), .ZN(G162) );
  NAND2_X1 U955 ( .A1(G103), .A2(n603), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G139), .A2(n605), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n865) );
  NAND2_X1 U958 ( .A1(G115), .A2(n871), .ZN(n862) );
  NAND2_X1 U959 ( .A1(G127), .A2(n872), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(KEYINPUT47), .B(n863), .Z(n864) );
  NOR2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n929) );
  XOR2_X1 U963 ( .A(G162), .B(n929), .Z(n867) );
  XNOR2_X1 U964 ( .A(G160), .B(G164), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n880) );
  NAND2_X1 U966 ( .A1(G106), .A2(n603), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G142), .A2(n605), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n870), .B(KEYINPUT45), .ZN(n877) );
  NAND2_X1 U970 ( .A1(G118), .A2(n871), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G130), .A2(n872), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U973 ( .A(KEYINPUT114), .B(n875), .Z(n876) );
  NAND2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U975 ( .A(n878), .B(KEYINPUT48), .ZN(n879) );
  XOR2_X1 U976 ( .A(n880), .B(n879), .Z(n883) );
  XNOR2_X1 U977 ( .A(n881), .B(KEYINPUT46), .ZN(n882) );
  XNOR2_X1 U978 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n914), .B(n884), .ZN(n888) );
  XNOR2_X1 U980 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n888), .B(n887), .ZN(n889) );
  NOR2_X1 U982 ( .A1(G37), .A2(n889), .ZN(G395) );
  XNOR2_X1 U983 ( .A(n1007), .B(KEYINPUT115), .ZN(n891) );
  XNOR2_X1 U984 ( .A(G171), .B(n1008), .ZN(n890) );
  XNOR2_X1 U985 ( .A(n891), .B(n890), .ZN(n894) );
  XNOR2_X1 U986 ( .A(G286), .B(n892), .ZN(n893) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U988 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U989 ( .A(G2443), .B(G2427), .Z(n897) );
  XNOR2_X1 U990 ( .A(G2438), .B(G2454), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U992 ( .A(n898), .B(G2435), .Z(n900) );
  XNOR2_X1 U993 ( .A(G1341), .B(G1348), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U995 ( .A(G2430), .B(G2446), .Z(n902) );
  XNOR2_X1 U996 ( .A(KEYINPUT110), .B(G2451), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U998 ( .A(n904), .B(n903), .Z(n905) );
  NAND2_X1 U999 ( .A1(G14), .A2(n905), .ZN(n911) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(G225) );
  XOR2_X1 U1006 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1008 ( .A(G132), .ZN(G219) );
  INV_X1 U1009 ( .A(G120), .ZN(G236) );
  INV_X1 U1010 ( .A(G108), .ZN(G238) );
  INV_X1 U1011 ( .A(G82), .ZN(G220) );
  INV_X1 U1012 ( .A(G69), .ZN(G235) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(n911), .ZN(G401) );
  XNOR2_X1 U1015 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n936) );
  NOR2_X1 U1016 ( .A1(n913), .A2(n912), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(G160), .B(G2084), .ZN(n915) );
  NAND2_X1 U1018 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1020 ( .A(KEYINPUT117), .B(n918), .Z(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n927) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n923), .Z(n925) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT118), .B(n928), .ZN(n934) );
  XOR2_X1 U1028 ( .A(G2072), .B(n929), .Z(n931) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n932), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(n936), .B(n935), .ZN(n937) );
  XOR2_X1 U1034 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n985) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n985), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n938), .A2(G29), .ZN(n992) );
  XOR2_X1 U1037 ( .A(G1976), .B(G23), .Z(n940) );
  XOR2_X1 U1038 ( .A(G1971), .B(G22), .Z(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G24), .B(G1986), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1042 ( .A(KEYINPUT58), .B(n943), .Z(n960) );
  XOR2_X1 U1043 ( .A(G1961), .B(G5), .Z(n955) );
  XNOR2_X1 U1044 ( .A(G20), .B(n944), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G19), .ZN(n945) );
  NOR2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1048 ( .A(KEYINPUT125), .B(n947), .Z(n948) );
  NAND2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n952) );
  XOR2_X1 U1050 ( .A(KEYINPUT59), .B(G1348), .Z(n950) );
  XNOR2_X1 U1051 ( .A(G4), .B(n950), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1053 ( .A(KEYINPUT60), .B(n953), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(G21), .B(G1966), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1057 ( .A(KEYINPUT126), .B(n958), .Z(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1059 ( .A(KEYINPUT61), .B(n961), .Z(n963) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT124), .ZN(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n990) );
  XOR2_X1 U1062 ( .A(KEYINPUT122), .B(G34), .Z(n965) );
  XNOR2_X1 U1063 ( .A(G2084), .B(KEYINPUT54), .ZN(n964) );
  XNOR2_X1 U1064 ( .A(n965), .B(n964), .ZN(n983) );
  XNOR2_X1 U1065 ( .A(G2090), .B(G35), .ZN(n981) );
  XNOR2_X1 U1066 ( .A(G25), .B(n966), .ZN(n967) );
  NAND2_X1 U1067 ( .A1(n967), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(G32), .B(n968), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(n969), .B(G27), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(G2067), .B(G26), .ZN(n971) );
  XNOR2_X1 U1071 ( .A(G2072), .B(G33), .ZN(n970) );
  NOR2_X1 U1072 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1073 ( .A(KEYINPUT121), .B(n972), .ZN(n973) );
  NOR2_X1 U1074 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1075 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1077 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  NOR2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n985), .B(n984), .ZN(n987) );
  INV_X1 U1081 ( .A(G29), .ZN(n986) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n988), .ZN(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n1018) );
  XOR2_X1 U1086 ( .A(KEYINPUT56), .B(G16), .Z(n1016) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G299), .ZN(n993) );
  XNOR2_X1 U1088 ( .A(n993), .B(KEYINPUT123), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(G168), .B(G1966), .ZN(n995) );
  NAND2_X1 U1090 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(n996), .B(KEYINPUT57), .ZN(n997) );
  NAND2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n1014) );
  NAND2_X1 U1093 ( .A1(G1971), .A2(G303), .ZN(n999) );
  NAND2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XNOR2_X1 U1095 ( .A(G1961), .B(G301), .ZN(n1001) );
  NOR2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G1341), .B(n1007), .ZN(n1010) );
  XOR2_X1 U1100 ( .A(G1348), .B(n1008), .Z(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(n1019), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

