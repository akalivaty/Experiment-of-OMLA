//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G210), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(G237), .A3(G953), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT75), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT74), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT67), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n196), .A3(G137), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n201), .A2(new_n202), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n196), .B2(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n197), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n204), .A2(new_n209), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT64), .B(G143), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(new_n216), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n218), .A3(G146), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n221), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n223), .A2(new_n225), .A3(new_n216), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(G143), .B2(new_n216), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n214), .A2(new_n215), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n208), .A2(new_n213), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT72), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n221), .A2(new_n227), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT66), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n221), .A2(new_n227), .A3(new_n243), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n201), .A2(new_n206), .A3(new_n207), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n208), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n240), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n232), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT71), .ZN(new_n253));
  INV_X1    g067(.A(new_n251), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n242), .B2(new_n244), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(new_n248), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n239), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT70), .A2(G119), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT70), .A2(G119), .ZN(new_n260));
  OAI21_X1  g074(.A(G116), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G119), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT2), .B(G113), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n264), .B2(new_n265), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n269), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n230), .A2(new_n235), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n237), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n252), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n258), .A2(new_n271), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT76), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n236), .A2(new_n238), .ZN(new_n279));
  AND4_X1   g093(.A1(new_n256), .A2(new_n245), .A3(new_n248), .A4(new_n251), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n256), .B1(new_n255), .B2(new_n248), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n271), .B(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n272), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n277), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n255), .A2(new_n248), .B1(new_n236), .B2(new_n238), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT77), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n271), .B1(new_n287), .B2(new_n288), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n277), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n278), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n252), .A2(new_n293), .A3(new_n274), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(KEYINPUT30), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n194), .B(new_n282), .C1(new_n297), .C2(new_n269), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n294), .B1(new_n258), .B2(new_n293), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n272), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n302), .A2(KEYINPUT31), .A3(new_n194), .A4(new_n282), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n195), .A2(new_n292), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n187), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n278), .A2(new_n194), .A3(new_n286), .A4(new_n291), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n282), .B1(new_n297), .B2(new_n269), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n309), .B2(new_n195), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n271), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n296), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT78), .A3(new_n282), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT78), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n296), .A2(new_n316), .A3(new_n313), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(KEYINPUT28), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n291), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n194), .A2(KEYINPUT29), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n312), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G472), .B1(new_n311), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n300), .A2(new_n303), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n291), .B1(new_n284), .B2(new_n285), .ZN(new_n324));
  AOI211_X1 g138(.A(KEYINPUT76), .B(new_n277), .C1(new_n282), .C2(new_n283), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n195), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n306), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT32), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n307), .A2(new_n322), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT16), .ZN(new_n331));
  INV_X1    g145(.A(G125), .ZN(new_n332));
  OR3_X1    g146(.A1(new_n332), .A2(KEYINPUT16), .A3(G140), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n331), .A2(G146), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G146), .B1(new_n331), .B2(new_n333), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(G128), .B1(new_n259), .B2(new_n260), .ZN(new_n337));
  INV_X1    g151(.A(G119), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G128), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT24), .B(G110), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n345));
  OR2_X1    g159(.A1(KEYINPUT70), .A2(G119), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT70), .A2(G119), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n228), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n337), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n259), .A2(new_n260), .A3(G128), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n340), .A2(new_n349), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G110), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n344), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT80), .B(G110), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n354), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n341), .A2(new_n342), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(KEYINPUT81), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n330), .A2(new_n364), .A3(new_n216), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n330), .B2(new_n216), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(new_n334), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT81), .B1(new_n361), .B2(new_n362), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n359), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT22), .B(G137), .Z(new_n372));
  INV_X1    g186(.A(G953), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n373), .A2(G221), .A3(G234), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n372), .B(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n375), .B(KEYINPUT83), .Z(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n359), .B(new_n375), .C1(new_n369), .C2(new_n370), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(G234), .B2(new_n312), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G902), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n312), .A3(new_n378), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT25), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n377), .A2(KEYINPUT25), .A3(new_n312), .A4(new_n378), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n386), .A2(KEYINPUT84), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(new_n389), .A3(new_n385), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n381), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n383), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n386), .A2(KEYINPUT84), .A3(new_n387), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n381), .A3(new_n390), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT85), .A3(new_n383), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(KEYINPUT9), .B(G234), .Z(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n400), .A2(new_n380), .A3(G953), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n220), .A2(new_n228), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n222), .A2(G128), .ZN(new_n404));
  OAI21_X1  g218(.A(G134), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n226), .A2(G128), .ZN(new_n406));
  INV_X1    g220(.A(new_n404), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n196), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G122), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G116), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n262), .A2(G122), .ZN(new_n412));
  INV_X1    g226(.A(G107), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OR3_X1    g228(.A1(new_n410), .A2(KEYINPUT14), .A3(G116), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n411), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G107), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT94), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT94), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n420), .A3(G107), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n409), .A2(new_n414), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n411), .A2(new_n412), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G107), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n414), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n408), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n226), .A2(KEYINPUT13), .A3(G128), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT93), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n407), .A2(KEYINPUT13), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n428), .A2(new_n429), .B1(new_n406), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n403), .A2(KEYINPUT93), .A3(KEYINPUT13), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n427), .B1(new_n433), .B2(G134), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n402), .B1(new_n423), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n196), .B1(new_n431), .B2(new_n432), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n422), .B(new_n401), .C1(new_n436), .C2(new_n427), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(KEYINPUT95), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT95), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(new_n402), .C1(new_n423), .C2(new_n434), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n312), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n443), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n438), .A2(new_n312), .A3(new_n445), .A4(new_n440), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G952), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(G953), .ZN(new_n449));
  NAND2_X1  g263(.A1(G234), .A2(G237), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT21), .B(G898), .Z(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(G902), .A3(G953), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(G475), .A2(G902), .ZN(new_n455));
  INV_X1    g269(.A(G237), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n456), .A2(new_n373), .A3(G143), .A4(G214), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n456), .A2(new_n373), .A3(G214), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT91), .B(new_n457), .C1(new_n220), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(KEYINPUT18), .A2(G131), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  OAI22_X1  g275(.A1(new_n365), .A2(new_n366), .B1(new_n216), .B2(new_n330), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n457), .B1(new_n220), .B2(new_n458), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G131), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n202), .B(new_n457), .C1(new_n220), .C2(new_n458), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(KEYINPUT17), .A3(G131), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n336), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G113), .B(G122), .ZN(new_n471));
  INV_X1    g285(.A(G104), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n463), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n330), .B(KEYINPUT19), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n216), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n465), .A2(new_n467), .ZN(new_n477));
  INV_X1    g291(.A(new_n334), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n473), .B1(new_n463), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n455), .B1(new_n474), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT20), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n483), .B(new_n455), .C1(new_n474), .C2(new_n480), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n473), .B1(new_n463), .B2(new_n470), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n312), .B1(new_n474), .B2(new_n485), .ZN(new_n486));
  XOR2_X1   g300(.A(KEYINPUT92), .B(G475), .Z(new_n487));
  AOI22_X1  g301(.A1(new_n482), .A2(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n447), .A2(KEYINPUT96), .A3(new_n454), .A4(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n454), .A3(new_n444), .A4(new_n446), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT96), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n413), .A2(G104), .ZN(new_n494));
  OR2_X1    g308(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n495));
  NAND2_X1  g309(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n472), .A2(G107), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n472), .A2(G107), .ZN(new_n499));
  NOR2_X1   g313(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G101), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n496), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n499), .B1(new_n503), .B2(new_n500), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT87), .B(G101), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n495), .A2(new_n494), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n498), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT4), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(G101), .C1(new_n497), .C2(new_n501), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n245), .A2(new_n251), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n494), .A2(new_n498), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G101), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n221), .A2(new_n227), .B1(new_n515), .B2(G128), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n221), .A2(new_n227), .A3(new_n229), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT10), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n248), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n273), .A2(new_n514), .A3(KEYINPUT10), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n511), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(G110), .B(G140), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n373), .A2(G227), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(KEYINPUT89), .A3(new_n526), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n273), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n507), .A2(new_n513), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n221), .A2(new_n227), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n515), .A2(G128), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n532), .B1(new_n535), .B2(new_n230), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n248), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT12), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(KEYINPUT12), .B(new_n248), .C1(new_n531), .C2(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n529), .A2(new_n530), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n523), .ZN(new_n543));
  AND4_X1   g357(.A1(new_n245), .A2(new_n251), .A3(new_n508), .A4(new_n510), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n522), .B1(new_n536), .B2(KEYINPUT10), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n248), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT88), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n511), .A2(new_n520), .A3(new_n522), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n248), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n543), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n542), .B1(new_n551), .B2(new_n526), .ZN(new_n552));
  INV_X1    g366(.A(G469), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n312), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n548), .A2(new_n549), .A3(new_n248), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n549), .B1(new_n548), .B2(new_n248), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n523), .B(new_n526), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n526), .B1(new_n541), .B2(new_n523), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n559), .A3(G469), .ZN(new_n560));
  NAND2_X1  g374(.A1(G469), .A2(G902), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(G214), .B1(G237), .B2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G210), .B1(G237), .B2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n264), .A2(new_n266), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n261), .A2(KEYINPUT5), .A3(new_n263), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n568), .B(G113), .C1(KEYINPUT5), .C2(new_n261), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n514), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n508), .A2(new_n510), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(new_n269), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT6), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G122), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT90), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT90), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n572), .A2(new_n578), .A3(new_n573), .A4(new_n575), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n273), .A2(G125), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n245), .A2(new_n251), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(G125), .ZN(new_n583));
  INV_X1    g397(.A(G224), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G953), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n581), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n255), .B2(new_n332), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n585), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n572), .A2(new_n575), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n570), .B(new_n574), .C1(new_n571), .C2(new_n269), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(KEYINPUT6), .A3(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n580), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n583), .A2(KEYINPUT7), .A3(new_n586), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n574), .B(KEYINPUT8), .ZN(new_n597));
  INV_X1    g411(.A(new_n568), .ZN(new_n598));
  OAI21_X1  g412(.A(G113), .B1(new_n261), .B2(KEYINPUT5), .ZN(new_n599));
  OAI22_X1  g413(.A1(new_n598), .A2(new_n599), .B1(new_n264), .B2(new_n266), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n532), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n569), .A2(new_n567), .B1(new_n513), .B2(new_n507), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n603), .A2(new_n593), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n589), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n596), .A2(new_n604), .A3(new_n590), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n312), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n566), .B1(new_n595), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n580), .A2(new_n591), .A3(new_n594), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(new_n312), .A3(new_n565), .A4(new_n607), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n564), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G221), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n399), .B2(new_n312), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AND4_X1   g429(.A1(new_n493), .A2(new_n562), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n329), .A2(new_n398), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(new_n505), .Z(G3));
  AOI22_X1  g432(.A1(new_n301), .A2(new_n272), .B1(new_n271), .B2(new_n258), .ZN(new_n619));
  AOI21_X1  g433(.A(KEYINPUT31), .B1(new_n619), .B2(new_n194), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n298), .A2(new_n299), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n326), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n312), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n327), .B1(new_n623), .B2(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n562), .A2(new_n615), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n612), .A2(new_n454), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n438), .A2(new_n628), .A3(new_n440), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n435), .A2(KEYINPUT33), .A3(new_n437), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n442), .A2(G902), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n441), .A2(KEYINPUT97), .A3(new_n442), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT97), .B1(new_n441), .B2(new_n442), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n488), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n627), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n624), .A2(new_n398), .A3(new_n626), .A4(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  NOR2_X1   g456(.A1(new_n447), .A2(new_n637), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n627), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n624), .A2(new_n398), .A3(new_n626), .A4(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NOR2_X1   g462(.A1(new_n376), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n371), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n382), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n388), .B2(new_n391), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT98), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n396), .A2(new_n654), .A3(new_n651), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n624), .A2(new_n616), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AND3_X1   g473(.A1(new_n562), .A2(new_n612), .A3(new_n615), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n451), .B(KEYINPUT99), .Z(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(G900), .B2(new_n453), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n643), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n329), .A2(new_n660), .A3(new_n656), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  XNOR2_X1  g480(.A(new_n663), .B(KEYINPUT39), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n626), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n315), .A2(new_n195), .A3(new_n317), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n671), .A3(new_n298), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n312), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n671), .B1(new_n670), .B2(new_n298), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n307), .A2(new_n328), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n447), .A2(new_n488), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n563), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n609), .A2(KEYINPUT38), .A3(new_n611), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT38), .B1(new_n609), .B2(new_n611), .ZN(new_n681));
  NOR4_X1   g495(.A1(new_n652), .A2(new_n679), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n669), .A2(new_n676), .A3(new_n677), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n220), .ZN(G45));
  INV_X1    g498(.A(new_n638), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n663), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n329), .A2(new_n660), .A3(new_n656), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  OAI21_X1  g503(.A(new_n523), .B1(new_n555), .B2(new_n556), .ZN(new_n690));
  INV_X1    g504(.A(new_n526), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n527), .A2(new_n528), .B1(new_n540), .B2(new_n539), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n690), .A2(new_n691), .B1(new_n692), .B2(new_n530), .ZN(new_n693));
  OAI21_X1  g507(.A(G469), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n615), .A3(new_n554), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n329), .A2(new_n398), .A3(new_n639), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND4_X1  g513(.A1(new_n329), .A2(new_n398), .A3(new_n645), .A4(new_n696), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  NOR3_X1   g515(.A1(new_n693), .A2(G469), .A3(G902), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n553), .B1(new_n552), .B2(new_n312), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(KEYINPUT101), .A3(new_n612), .A4(new_n615), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n612), .A2(new_n615), .A3(new_n694), .A4(new_n554), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n329), .A3(new_n493), .A4(new_n656), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  INV_X1    g525(.A(new_n392), .ZN(new_n712));
  OAI21_X1  g526(.A(G472), .B1(new_n304), .B2(G902), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n319), .A2(new_n195), .B1(new_n300), .B2(new_n303), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n714), .B1(new_n715), .B2(new_n306), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n620), .A2(new_n621), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n194), .B1(new_n318), .B2(new_n291), .ZN(new_n718));
  OAI211_X1 g532(.A(KEYINPUT102), .B(new_n305), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n712), .A2(new_n713), .A3(new_n716), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n678), .A2(new_n454), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n706), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  AND3_X1   g538(.A1(new_n713), .A2(new_n716), .A3(new_n719), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n709), .A3(new_n652), .A4(new_n687), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  NAND3_X1  g541(.A1(new_n609), .A2(new_n563), .A3(new_n611), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n561), .B(KEYINPUT103), .Z(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n554), .A2(new_n560), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n609), .A2(new_n733), .A3(new_n563), .A4(new_n611), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n729), .A2(new_n732), .A3(new_n615), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n686), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n329), .A3(new_n712), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n739));
  INV_X1    g553(.A(new_n735), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n329), .A2(new_n739), .A3(new_n398), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n202), .ZN(G33));
  NAND4_X1  g557(.A1(new_n329), .A2(new_n398), .A3(new_n664), .A4(new_n740), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  NAND3_X1  g559(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT45), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n527), .B1(new_n547), .B2(new_n550), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n747), .B1(new_n748), .B2(new_n558), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n749), .A3(G469), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n731), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(KEYINPUT46), .A3(new_n731), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n554), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n615), .A3(new_n667), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT105), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n729), .A2(new_n734), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n441), .A2(new_n442), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT97), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n629), .A2(new_n630), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n762), .A2(new_n633), .B1(new_n763), .B2(new_n631), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n759), .B1(new_n764), .B2(new_n637), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n636), .A2(KEYINPUT43), .A3(new_n488), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n765), .A2(new_n766), .B1(new_n396), .B2(new_n651), .ZN(new_n767));
  INV_X1    g581(.A(G472), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n622), .B2(new_n312), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n327), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT44), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n713), .B1(new_n304), .B2(new_n306), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n767), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n758), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n757), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  NAND4_X1  g591(.A1(new_n685), .A2(new_n729), .A3(new_n663), .A4(new_n734), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n329), .A2(new_n398), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n755), .A2(new_n615), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n755), .A2(new_n782), .A3(new_n615), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NAND2_X1  g599(.A1(new_n448), .A2(new_n373), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n725), .A2(new_n652), .A3(new_n687), .A4(new_n740), .ZN(new_n787));
  INV_X1    g601(.A(new_n447), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n637), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n729), .A2(new_n789), .A3(new_n663), .A4(new_n734), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n329), .A2(new_n626), .A3(new_n656), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n787), .B(new_n744), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n742), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n617), .A2(new_n640), .A3(new_n646), .A4(new_n657), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT106), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n769), .A2(new_n625), .A3(new_n327), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n799), .B(new_n398), .C1(new_n639), .C2(new_n645), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(KEYINPUT106), .A3(new_n617), .A4(new_n657), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n723), .A2(new_n710), .A3(new_n697), .A4(new_n700), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n795), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n665), .A2(new_n688), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n732), .A2(new_n615), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n612), .A2(new_n663), .A3(new_n678), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n808), .A3(new_n652), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n676), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n806), .A2(KEYINPUT52), .A3(new_n726), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n726), .A2(new_n665), .A3(new_n688), .A4(new_n810), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT53), .B1(new_n805), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n794), .A2(new_n742), .A3(new_n803), .ZN(new_n817));
  AND4_X1   g631(.A1(KEYINPUT53), .A2(new_n815), .A3(new_n817), .A4(new_n802), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT54), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n795), .A2(new_n802), .A3(new_n804), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n812), .B(KEYINPUT52), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n815), .A2(new_n817), .A3(KEYINPUT53), .A4(new_n802), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n765), .A2(new_n766), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n661), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n720), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n709), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n758), .A2(KEYINPUT114), .A3(new_n695), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT114), .B1(new_n758), .B2(new_n695), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n676), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n451), .B1(new_n394), .B2(new_n397), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n832), .B(new_n449), .C1(new_n638), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n838), .A2(new_n638), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n449), .A4(new_n832), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n329), .A2(new_n712), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT115), .B1(new_n835), .B2(new_n830), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n846), .B(new_n829), .C1(new_n833), .C2(new_n834), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n844), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT48), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT48), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n850), .B(new_n844), .C1(new_n845), .C2(new_n847), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n840), .A2(new_n843), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n681), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n609), .A2(KEYINPUT38), .A3(new_n611), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n563), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT109), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n696), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n564), .B1(new_n680), .B2(new_n681), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT109), .B1(new_n858), .B2(new_n695), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n831), .A2(KEYINPUT50), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n860), .A2(new_n720), .A3(new_n830), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n864), .B2(KEYINPUT110), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT110), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n831), .A2(new_n866), .A3(new_n860), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT112), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n865), .A2(new_n867), .A3(KEYINPUT112), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n862), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n781), .A2(new_n783), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n704), .A2(new_n614), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n758), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n875), .B2(new_n831), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n764), .A2(new_n488), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n725), .A2(new_n652), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n845), .B2(new_n847), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n876), .A2(new_n881), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n852), .B1(new_n871), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n865), .A2(new_n867), .A3(KEYINPUT112), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n861), .B1(new_n887), .B2(new_n868), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT113), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n881), .A2(new_n884), .A3(new_n882), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n875), .A2(new_n831), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n891), .A2(KEYINPUT108), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(KEYINPUT108), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT113), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n861), .B(new_n895), .C1(new_n887), .C2(new_n868), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n889), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n886), .B1(new_n897), .B2(new_n872), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n827), .B1(new_n898), .B2(KEYINPUT118), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n900), .B(new_n886), .C1(new_n872), .C2(new_n897), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n786), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n704), .B(KEYINPUT49), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n615), .A2(new_n563), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n636), .A2(new_n488), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n904), .B(new_n905), .C1(new_n853), .C2(new_n854), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n836), .A2(new_n903), .A3(new_n712), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n902), .A2(new_n907), .ZN(G75));
  NAND2_X1  g722(.A1(new_n580), .A2(new_n594), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n591), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT119), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n312), .B1(new_n824), .B2(new_n825), .ZN(new_n914));
  AOI211_X1 g728(.A(KEYINPUT55), .B(new_n913), .C1(new_n914), .C2(G210), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT55), .ZN(new_n916));
  OAI211_X1 g730(.A(G210), .B(G902), .C1(new_n816), .C2(new_n818), .ZN(new_n917));
  INV_X1    g731(.A(new_n913), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n911), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n373), .A2(G952), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n188), .B(new_n312), .C1(new_n824), .C2(new_n825), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT55), .B1(new_n923), .B2(new_n913), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n917), .A2(new_n916), .A3(new_n918), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n925), .A3(new_n910), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n920), .A2(new_n922), .A3(new_n926), .ZN(G51));
  XOR2_X1   g741(.A(new_n730), .B(KEYINPUT57), .Z(new_n928));
  OAI21_X1  g742(.A(new_n552), .B1(new_n827), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n914), .A2(G469), .A3(new_n746), .A4(new_n749), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n921), .B1(new_n929), .B2(new_n930), .ZN(G54));
  NAND3_X1  g745(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n474), .A2(new_n480), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n921), .ZN(G60));
  NAND2_X1  g750(.A1(new_n824), .A2(new_n825), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT54), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT59), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n938), .A2(new_n763), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n763), .B1(new_n938), .B2(new_n940), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n921), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n824), .B2(new_n825), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n379), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n921), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n946), .A2(new_n950), .A3(new_n650), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n950), .B1(new_n946), .B2(new_n650), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n949), .B(KEYINPUT61), .C1(new_n951), .C2(new_n952), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(G66));
  AOI21_X1  g771(.A(new_n373), .B1(new_n452), .B2(G224), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n802), .A2(new_n804), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n802), .A2(KEYINPUT121), .A3(new_n804), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n958), .B1(new_n963), .B2(new_n373), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n909), .B1(G898), .B2(new_n373), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n964), .B(new_n965), .Z(G69));
  AOI21_X1  g780(.A(new_n373), .B1(G227), .B2(G900), .ZN(new_n967));
  AND4_X1   g781(.A1(new_n329), .A2(new_n712), .A3(new_n612), .A4(new_n678), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n757), .B1(new_n775), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n742), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n726), .A2(new_n665), .A3(new_n688), .ZN(new_n971));
  INV_X1    g785(.A(new_n744), .ZN(new_n972));
  INV_X1    g786(.A(new_n783), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n782), .B1(new_n755), .B2(new_n615), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n975), .B2(new_n779), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AND4_X1   g793(.A1(new_n738), .A2(new_n784), .A3(new_n741), .A4(new_n744), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n980), .A2(KEYINPUT124), .A3(new_n971), .A4(new_n969), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n373), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n297), .B(new_n475), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(G900), .B2(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n967), .B1(new_n985), .B2(KEYINPUT123), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT122), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n685), .A2(new_n987), .A3(new_n643), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT122), .B1(new_n644), .B2(new_n638), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n988), .A2(new_n758), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n668), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n990), .A2(new_n991), .A3(new_n329), .A4(new_n398), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n771), .A2(new_n774), .ZN(new_n993));
  INV_X1    g807(.A(new_n758), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT105), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n756), .B(new_n996), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n784), .B(new_n992), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n683), .A2(new_n806), .A3(new_n726), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n971), .A2(KEYINPUT62), .A3(new_n683), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n983), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n985), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n986), .B(new_n1005), .Z(G72));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n309), .A2(new_n195), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n298), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n937), .A2(new_n1007), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1007), .B1(new_n937), .B2(new_n1012), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1003), .A2(new_n961), .A3(new_n962), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n1009), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n619), .A2(new_n195), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT125), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1017), .A2(KEYINPUT125), .A3(new_n1018), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT127), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n979), .A2(new_n981), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1009), .B1(new_n1025), .B2(new_n963), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n309), .A2(new_n194), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n921), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1015), .A2(new_n1023), .A3(new_n1024), .A4(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1028), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1030));
  AOI21_X1  g844(.A(KEYINPUT125), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1018), .ZN(new_n1032));
  AOI211_X1 g846(.A(new_n1020), .B(new_n1032), .C1(new_n1016), .C2(new_n1009), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(KEYINPUT127), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1029), .A2(new_n1035), .ZN(G57));
endmodule


