//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT97), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n202), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G71gat), .B(G78gat), .Z(new_n209));
  AND2_X1   g008(.A1(new_n207), .A2(new_n203), .ZN(new_n210));
  OR3_X1    g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n208), .B2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT21), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G231gat), .A2(G233gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(G127gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(G1gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT16), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n220), .B2(new_n219), .ZN(new_n222));
  INV_X1    g021(.A(G8gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n224), .B(KEYINPUT94), .Z(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n223), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n226), .B(KEYINPUT95), .Z(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n214), .B2(new_n213), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n218), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n232));
  INV_X1    g031(.A(G155gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G183gat), .B(G211gat), .Z(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT100), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(G85gat), .A3(G92gat), .A4(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G85gat), .ZN(new_n246));
  INV_X1    g045(.A(G92gat), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n241), .B(new_n242), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G99gat), .A2(G106gat), .ZN(new_n249));
  AOI22_X1  g048(.A1(KEYINPUT8), .A2(new_n249), .B1(new_n246), .B2(new_n247), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n245), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT101), .ZN(new_n252));
  XOR2_X1   g051(.A(G99gat), .B(G106gat), .Z(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n252), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G43gat), .B(G50gat), .Z(new_n256));
  INV_X1    g055(.A(KEYINPUT15), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT92), .B(G36gat), .Z(new_n259));
  INV_X1    g058(.A(G29gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(G29gat), .A2(G36gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT14), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n258), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT93), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n256), .A2(new_n257), .ZN(new_n266));
  OR4_X1    g065(.A1(new_n258), .A2(new_n266), .A3(new_n261), .A4(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n255), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT41), .ZN(new_n270));
  NAND2_X1  g069(.A1(G232gat), .A2(G233gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT98), .Z(new_n272));
  INV_X1    g071(.A(KEYINPUT17), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n265), .A2(KEYINPUT17), .A3(new_n267), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI221_X1 g075(.A(new_n269), .B1(new_n270), .B2(new_n272), .C1(new_n276), .C2(new_n255), .ZN(new_n277));
  XOR2_X1   g076(.A(G190gat), .B(G218gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT102), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n280), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT103), .B1(new_n277), .B2(new_n280), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n272), .A2(new_n270), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT99), .ZN(new_n286));
  XOR2_X1   g085(.A(G134gat), .B(G162gat), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n283), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n281), .A2(KEYINPUT103), .A3(new_n282), .A4(new_n288), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n240), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n213), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT104), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n251), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n255), .B(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G230gat), .A2(G233gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G120gat), .B(G148gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT105), .ZN(new_n302));
  XNOR2_X1  g101(.A(G176gat), .B(G204gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n294), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n300), .B(new_n304), .C1(new_n308), .C2(new_n299), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n299), .B(KEYINPUT106), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n300), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n309), .B1(new_n314), .B2(new_n304), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n293), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  INV_X1    g118(.A(G218gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G211gat), .A2(G218gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(KEYINPUT75), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT22), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n327));
  AND2_X1   g126(.A1(G211gat), .A2(G218gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G211gat), .A2(G218gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n333));
  OAI21_X1  g132(.A(G204gat), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g133(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n335));
  INV_X1    g134(.A(G204gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n331), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n326), .A2(new_n330), .A3(new_n334), .A4(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n334), .A2(new_n337), .A3(new_n323), .A4(new_n325), .ZN(new_n339));
  INV_X1    g138(.A(new_n330), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT83), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT3), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n344), .B2(new_n343), .ZN(new_n346));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347));
  INV_X1    g146(.A(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n233), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n349), .B2(KEYINPUT2), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n351));
  INV_X1    g150(.A(G148gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(G141gat), .ZN(new_n353));
  INV_X1    g152(.A(G141gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(G148gat), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n351), .A2(new_n352), .A3(G141gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n350), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G141gat), .B(G148gat), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n347), .B(new_n349), .C1(new_n358), .C2(KEYINPUT2), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n346), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G228gat), .A2(G233gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n338), .A2(new_n341), .A3(KEYINPUT76), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT76), .B1(new_n338), .B2(new_n341), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n342), .B1(new_n360), .B2(KEYINPUT3), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n343), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n360), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n357), .A2(KEYINPUT80), .A3(new_n359), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n339), .A2(new_n340), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n339), .A2(new_n340), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(new_n363), .A3(new_n367), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n362), .B(KEYINPUT81), .Z(new_n384));
  AOI21_X1  g183(.A(new_n370), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n384), .ZN(new_n386));
  AOI211_X1 g185(.A(KEYINPUT82), .B(new_n386), .C1(new_n377), .C2(new_n382), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n369), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G22gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n390));
  INV_X1    g189(.A(G22gat), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n369), .B(new_n391), .C1(new_n385), .C2(new_n387), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(KEYINPUT31), .B(G50gat), .Z(new_n394));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n393), .A2(new_n397), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n392), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT84), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n366), .ZN(new_n403));
  INV_X1    g202(.A(G226gat), .ZN(new_n404));
  INV_X1    g203(.A(G233gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(KEYINPUT29), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(G169gat), .ZN(new_n410));
  INV_X1    g209(.A(G176gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT66), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT66), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G176gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT23), .ZN(new_n417));
  INV_X1    g216(.A(G169gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT67), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n415), .A2(new_n420), .A3(KEYINPUT67), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n425), .A2(KEYINPUT65), .ZN(new_n426));
  NAND2_X1  g225(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n427));
  MUX2_X1   g226(.A(G183gat), .B(new_n427), .S(G190gat), .Z(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(KEYINPUT65), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT25), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n431), .A2(KEYINPUT68), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT68), .B1(new_n431), .B2(new_n432), .ZN(new_n434));
  INV_X1    g233(.A(new_n425), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n419), .A2(new_n409), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(new_n432), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n438), .A3(new_n420), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n433), .A2(new_n434), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT27), .B(G183gat), .ZN(new_n442));
  INV_X1    g241(.A(G190gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT28), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT69), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n444), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT26), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n419), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(G169gat), .B2(G176gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n419), .B2(new_n448), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n447), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT77), .B1(new_n441), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n431), .A2(new_n432), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n431), .A2(KEYINPUT68), .A3(new_n432), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n439), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT77), .ZN(new_n460));
  INV_X1    g259(.A(new_n453), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n408), .B1(new_n454), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n461), .A3(new_n406), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n403), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n454), .A2(new_n406), .A3(new_n462), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n407), .B1(new_n441), .B2(new_n453), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n366), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT30), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n466), .A2(KEYINPUT30), .A3(new_n469), .A4(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n467), .A2(new_n366), .A3(new_n468), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n440), .B1(new_n455), .B2(new_n456), .ZN(new_n479));
  AOI211_X1 g278(.A(KEYINPUT77), .B(new_n453), .C1(new_n479), .C2(new_n458), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n460), .B1(new_n459), .B2(new_n461), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n407), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n366), .B1(new_n482), .B2(new_n464), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT78), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n485), .A3(new_n469), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n472), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n477), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489));
  XNOR2_X1  g288(.A(G113gat), .B(G120gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT70), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT1), .ZN(new_n493));
  XNOR2_X1  g292(.A(G127gat), .B(G134gat), .ZN(new_n494));
  INV_X1    g293(.A(G120gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n494), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(KEYINPUT1), .B2(new_n490), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT4), .B1(new_n500), .B2(new_n360), .ZN(new_n501));
  INV_X1    g300(.A(new_n376), .ZN(new_n502));
  INV_X1    g301(.A(new_n500), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n501), .B1(new_n504), .B2(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n500), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G225gat), .A2(G233gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n509), .A2(KEYINPUT5), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT5), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n500), .B(new_n360), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(new_n511), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n503), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n500), .A2(new_n360), .ZN(new_n518));
  OAI221_X1 g317(.A(new_n510), .B1(new_n518), .B2(KEYINPUT4), .C1(new_n507), .C2(new_n508), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G1gat), .B(G29gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT0), .ZN(new_n523));
  XNOR2_X1  g322(.A(G57gat), .B(G85gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n489), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n521), .A2(new_n526), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n402), .B1(new_n488), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT71), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n500), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n533), .B(new_n535), .C1(new_n441), .C2(new_n453), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n459), .A2(new_n534), .A3(new_n500), .A4(new_n461), .ZN(new_n537));
  NAND2_X1  g336(.A1(G227gat), .A2(G233gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n538), .B(KEYINPUT64), .Z(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT33), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G43gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(G71gat), .B(G99gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n540), .B(KEYINPUT32), .C1(new_n541), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n540), .B2(KEYINPUT32), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n540), .A2(new_n541), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT72), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT72), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n551), .A3(new_n548), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n546), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n537), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n538), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT34), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n539), .A2(KEYINPUT34), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n532), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n547), .A2(new_n551), .A3(new_n548), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n551), .B1(new_n547), .B2(new_n548), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n545), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(KEYINPUT73), .A3(new_n559), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n560), .B(new_n545), .C1(new_n562), .C2(new_n563), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n561), .A2(KEYINPUT36), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n559), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n566), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n531), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT37), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n454), .A2(new_n462), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n465), .B1(new_n575), .B2(new_n407), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n574), .B(new_n469), .C1(new_n576), .C2(new_n366), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT87), .ZN(new_n578));
  INV_X1    g377(.A(new_n472), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT87), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n466), .A2(new_n580), .A3(new_n574), .A4(new_n469), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n574), .B1(new_n484), .B2(new_n486), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n573), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT88), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT88), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n586), .B(new_n573), .C1(new_n582), .C2(new_n583), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n529), .A2(new_n473), .ZN(new_n588));
  INV_X1    g387(.A(new_n582), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n467), .A2(new_n468), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n574), .B1(new_n590), .B2(new_n403), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n366), .B1(new_n463), .B2(new_n465), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n573), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n588), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n585), .A2(new_n587), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n486), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n485), .B1(new_n466), .B2(new_n469), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n579), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT85), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n598), .A2(new_n599), .A3(new_n475), .A4(new_n476), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT85), .B1(new_n477), .B2(new_n487), .ZN(new_n601));
  INV_X1    g400(.A(new_n509), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n510), .B1(new_n505), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n526), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT39), .B1(new_n515), .B2(new_n511), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n609), .A2(new_n528), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n600), .A2(new_n601), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n402), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n572), .B1(new_n595), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n402), .A2(new_n566), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n615), .A2(KEYINPUT89), .A3(new_n561), .A4(new_n565), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n561), .A2(new_n565), .A3(new_n566), .A4(new_n402), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT89), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT35), .ZN(new_n620));
  NOR4_X1   g419(.A1(new_n477), .A2(new_n487), .A3(new_n529), .A4(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n616), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  AND4_X1   g421(.A1(new_n530), .A2(new_n402), .A3(new_n568), .A4(new_n566), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n600), .A2(new_n601), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT35), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n614), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n229), .A2(new_n275), .A3(new_n274), .ZN(new_n628));
  NAND2_X1  g427(.A1(G229gat), .A2(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n228), .A2(new_n268), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT18), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n228), .B(new_n268), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n629), .B(KEYINPUT13), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n632), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT91), .ZN(new_n639));
  XNOR2_X1  g438(.A(G113gat), .B(G141gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT90), .B(G197gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT11), .B(G169gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n638), .A2(KEYINPUT91), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n627), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n650), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n318), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n529), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  AND4_X1   g457(.A1(new_n601), .A2(new_n655), .A3(new_n600), .A4(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(KEYINPUT42), .ZN(new_n660));
  INV_X1    g459(.A(new_n624), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n223), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT42), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(G1325gat));
  INV_X1    g463(.A(new_n655), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n567), .A2(new_n571), .ZN(new_n666));
  OAI21_X1  g465(.A(G15gat), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n569), .A2(G15gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n667), .B1(new_n665), .B2(new_n668), .ZN(G1326gat));
  INV_X1    g468(.A(new_n402), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  NOR2_X1   g472(.A1(new_n240), .A2(new_n316), .ZN(new_n674));
  INV_X1    g473(.A(new_n292), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n653), .B2(new_n654), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n530), .A2(G29gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT45), .ZN(new_n681));
  INV_X1    g480(.A(new_n676), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n585), .A2(new_n587), .A3(new_n594), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n402), .A3(new_n612), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n625), .B1(new_n684), .B2(new_n572), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n652), .B(new_n649), .C1(new_n685), .C2(new_n622), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT96), .B1(new_n627), .B2(new_n650), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n682), .B(new_n679), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT107), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n680), .A2(new_n681), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n681), .B1(new_n680), .B2(new_n689), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n692), .B(new_n292), .C1(new_n685), .C2(new_n622), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT44), .B1(new_n627), .B2(new_n675), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n650), .A2(new_n674), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT108), .Z(new_n697));
  AND2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(new_n529), .ZN(new_n699));
  OAI22_X1  g498(.A1(new_n690), .A2(new_n691), .B1(new_n699), .B2(new_n260), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n677), .A2(new_n661), .A3(new_n259), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n698), .A2(new_n661), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n702), .B(new_n703), .C1(new_n704), .C2(new_n259), .ZN(G1329gat));
  NAND2_X1  g504(.A1(new_n627), .A2(new_n675), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n692), .ZN(new_n707));
  INV_X1    g506(.A(new_n666), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n627), .A2(KEYINPUT44), .A3(new_n675), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .A4(new_n697), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G43gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n569), .A2(G43gat), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT109), .B1(new_n677), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n682), .B(new_n712), .C1(new_n686), .C2(new_n687), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n711), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g518(.A(KEYINPUT47), .B(new_n711), .C1(new_n713), .C2(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1330gat));
  XOR2_X1   g520(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n722));
  NOR2_X1   g521(.A1(new_n402), .A2(G50gat), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n682), .B(new_n723), .C1(new_n686), .C2(new_n687), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT111), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n670), .A3(new_n709), .A4(new_n697), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G50gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n724), .A2(KEYINPUT111), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n722), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(KEYINPUT48), .A3(new_n724), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  NOR3_X1   g531(.A1(new_n650), .A2(new_n293), .A3(new_n315), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT112), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n622), .B2(new_n685), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n529), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT113), .B(G57gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1332gat));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n661), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT49), .B(G64gat), .Z(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n739), .B2(new_n741), .ZN(G1333gat));
  AOI21_X1  g541(.A(new_n205), .B1(new_n735), .B2(new_n708), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n569), .A2(G71gat), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n735), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n735), .A2(new_n670), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n650), .A2(new_n240), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n316), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n707), .A2(new_n709), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT114), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n707), .A2(new_n754), .A3(new_n709), .A4(new_n751), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(new_n529), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n627), .A2(new_n675), .A3(new_n749), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n292), .B1(new_n685), .B2(new_n622), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n749), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n316), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n529), .A2(new_n246), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n756), .A2(new_n246), .B1(new_n763), .B2(new_n764), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n752), .B2(new_n624), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n661), .A2(new_n247), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n766), .B(new_n767), .C1(new_n763), .C2(new_n768), .ZN(new_n769));
  AOI211_X1 g568(.A(new_n315), .B(new_n768), .C1(new_n759), .C2(new_n761), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n661), .A3(new_n755), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(G92gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n772), .B2(new_n767), .ZN(G1337gat));
  NAND3_X1  g572(.A1(new_n753), .A2(new_n708), .A3(new_n755), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G99gat), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n569), .A2(G99gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n763), .B2(new_n776), .ZN(G1338gat));
  NAND4_X1  g576(.A1(new_n695), .A2(KEYINPUT116), .A3(new_n670), .A4(new_n751), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n707), .A2(new_n670), .A3(new_n709), .A4(new_n751), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n781), .A3(G106gat), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n402), .A2(G106gat), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT51), .B1(new_n760), .B2(new_n749), .ZN(new_n784));
  AND4_X1   g583(.A1(KEYINPUT51), .A2(new_n627), .A3(new_n675), .A4(new_n749), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n316), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT53), .B1(new_n786), .B2(KEYINPUT115), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n762), .A2(new_n788), .A3(new_n316), .A4(new_n783), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n782), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n786), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n753), .A2(new_n670), .A3(new_n755), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(G106gat), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(G1339gat));
  INV_X1    g594(.A(new_n240), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n308), .A2(new_n299), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n306), .A2(new_n310), .A3(new_n307), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(KEYINPUT54), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n308), .A2(new_n800), .A3(new_n311), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n304), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n309), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n304), .A4(new_n801), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n804), .A2(new_n646), .A3(new_n648), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n634), .A2(new_n635), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n629), .B1(new_n628), .B2(new_n630), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n644), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n633), .A2(new_n636), .A3(new_n637), .A4(new_n647), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n316), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n675), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n804), .A2(new_n805), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n290), .A2(new_n291), .A3(new_n809), .A4(new_n810), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n796), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n317), .A2(new_n649), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n661), .A2(new_n530), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n569), .A2(new_n670), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(G113gat), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n822), .A2(new_n823), .A3(new_n649), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n616), .A2(new_n619), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n820), .A2(new_n825), .A3(new_n650), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n824), .B1(new_n823), .B2(new_n826), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n822), .B2(new_n315), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n820), .A2(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n316), .A2(new_n495), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT117), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n828), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT118), .Z(G1341gat));
  OAI21_X1  g632(.A(G127gat), .B1(new_n822), .B2(new_n796), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n796), .A2(G127gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n829), .B2(new_n835), .ZN(G1342gat));
  OR3_X1    g635(.A1(new_n829), .A2(G134gat), .A3(new_n292), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n822), .B2(new_n292), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n670), .A3(new_n666), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n354), .B1(new_n842), .B2(new_n649), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n819), .A2(new_n666), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n402), .B1(new_n816), .B2(new_n817), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n846), .B2(KEYINPUT119), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n845), .B(KEYINPUT57), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(KEYINPUT119), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n649), .A2(new_n354), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n843), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(G1344gat));
  NOR3_X1   g653(.A1(new_n842), .A2(G148gat), .A3(new_n315), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT120), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n849), .A2(new_n315), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G148gat), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n848), .A2(new_n666), .A3(new_n316), .A4(new_n819), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n858), .B1(new_n861), .B2(G148gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n856), .B1(new_n860), .B2(new_n862), .ZN(G1345gat));
  OAI21_X1  g662(.A(G155gat), .B1(new_n849), .B2(new_n796), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n240), .A2(new_n233), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n842), .B2(new_n865), .ZN(G1346gat));
  OAI21_X1  g665(.A(new_n348), .B1(new_n842), .B2(new_n292), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n292), .A2(new_n348), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n849), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n870), .B(new_n871), .ZN(G1347gat));
  NAND3_X1  g671(.A1(new_n818), .A2(new_n661), .A3(new_n623), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(new_n418), .A3(new_n649), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n624), .A2(new_n529), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n818), .A2(new_n825), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n818), .A2(KEYINPUT122), .A3(new_n825), .A4(new_n875), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n650), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n874), .B1(new_n880), .B2(new_n418), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT123), .ZN(G1348gat));
  AOI211_X1 g681(.A(new_n315), .B(new_n873), .C1(new_n412), .C2(new_n414), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n878), .A2(new_n316), .A3(new_n879), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n411), .ZN(G1349gat));
  OAI21_X1  g684(.A(G183gat), .B1(new_n873), .B2(new_n796), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n240), .A2(new_n442), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n876), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g688(.A1(new_n292), .A2(G190gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n878), .A2(new_n879), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT124), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n879), .A3(new_n893), .A4(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G190gat), .B1(new_n873), .B2(new_n292), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT61), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT125), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n895), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1351gat));
  AND2_X1   g701(.A1(new_n666), .A2(new_n875), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n845), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT126), .Z(new_n905));
  AOI21_X1  g704(.A(G197gat), .B1(new_n905), .B2(new_n650), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n848), .A2(new_n903), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n650), .A2(G197gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(G1352gat));
  NAND3_X1  g708(.A1(new_n848), .A2(new_n316), .A3(new_n903), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G204gat), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n845), .A2(new_n336), .A3(new_n316), .A4(new_n903), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n912), .B2(KEYINPUT62), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT62), .ZN(new_n915));
  OAI221_X1 g714(.A(new_n911), .B1(KEYINPUT62), .B2(new_n912), .C1(new_n914), .C2(new_n915), .ZN(G1353gat));
  NAND3_X1  g715(.A1(new_n905), .A2(new_n319), .A3(new_n240), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n848), .A2(new_n240), .A3(new_n903), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT63), .B1(new_n918), .B2(G211gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1354gat));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n320), .A3(new_n675), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n675), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n924), .B2(new_n320), .ZN(G1355gat));
endmodule


