//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n211), .B1(new_n212), .B2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G13), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n214), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n201), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n212), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n206), .A2(new_n207), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n218), .B(new_n230), .C1(new_n233), .C2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G226), .B(G232), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(KEYINPUT8), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT69), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n232), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n208), .A2(G20), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G150), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n231), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G50), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(new_n270), .B2(G20), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(G50), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  OAI211_X1 g0077(.A(G1), .B(G13), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(G223), .A2(G1698), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G222), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n284), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n279), .A2(KEYINPUT68), .A3(G222), .A4(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n278), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  AOI21_X1  g0095(.A(G1), .B1(new_n277), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n278), .A2(G274), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n296), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G226), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(KEYINPUT71), .A2(G179), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT71), .A2(G179), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n294), .B2(new_n302), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n275), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(G190), .B2(new_n303), .ZN(new_n313));
  INV_X1    g0113(.A(new_n268), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n259), .A2(new_n261), .B1(G150), .B2(new_n264), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(new_n263), .ZN(new_n316));
  INV_X1    g0116(.A(new_n274), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT9), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT9), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n269), .A2(new_n319), .A3(new_n274), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n313), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n313), .B2(new_n321), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n310), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G244), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n297), .B1(new_n300), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(G232), .A2(G1698), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n289), .A2(G238), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n279), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G107), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n278), .B1(new_n288), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n327), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G169), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n306), .B2(new_n333), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n256), .A2(new_n254), .ZN(new_n336));
  INV_X1    g0136(.A(new_n264), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n336), .A2(new_n337), .B1(new_n232), .B2(new_n280), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT15), .B(G87), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n260), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n268), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT73), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n271), .A2(G77), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(new_n273), .B2(G77), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n335), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT72), .B1(new_n333), .B2(new_n311), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n333), .A2(G190), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n333), .A2(KEYINPUT72), .A3(G190), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n350), .A2(new_n343), .A3(new_n345), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n325), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n264), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n280), .B2(new_n260), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT76), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n356), .A2(new_n357), .A3(new_n268), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(new_n356), .B2(new_n268), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT11), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT11), .B1(new_n358), .B2(new_n359), .ZN(new_n361));
  OR3_X1    g0161(.A1(new_n271), .A2(KEYINPUT12), .A3(G68), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT12), .B1(new_n271), .B2(G68), .ZN(new_n363));
  AOI22_X1  g0163(.A1(G68), .A2(new_n273), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n301), .A2(new_n289), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n225), .A2(G1698), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n285), .A2(new_n366), .A3(new_n287), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n368), .A2(KEYINPUT74), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT74), .B1(new_n368), .B2(new_n369), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n370), .A2(new_n371), .A3(new_n278), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n297), .B1(new_n300), .B2(new_n220), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT13), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n374), .A2(G190), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT13), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n278), .A2(G274), .A3(new_n296), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(G238), .B2(new_n299), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n371), .A2(new_n278), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n376), .B(new_n378), .C1(new_n379), .C2(new_n370), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n365), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n374), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(KEYINPUT75), .B(KEYINPUT13), .C1(new_n372), .C2(new_n373), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(G200), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(G169), .A3(new_n384), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT14), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT14), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n383), .A2(new_n389), .A3(G169), .A4(new_n384), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n374), .A2(new_n380), .A3(G179), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n365), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n354), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(G20), .B1(G159), .B2(new_n264), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT77), .B1(new_n276), .B2(KEYINPUT3), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT77), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(new_n286), .A3(G33), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n399), .A3(new_n285), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n232), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n202), .B1(new_n401), .B2(KEYINPUT7), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT79), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(KEYINPUT78), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT78), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n397), .A2(new_n399), .A3(new_n405), .A4(new_n285), .ZN(new_n406));
  NOR2_X1   g0206(.A1(KEYINPUT7), .A2(G20), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n402), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n403), .B1(new_n402), .B2(new_n408), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT16), .B(new_n396), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  INV_X1    g0212(.A(new_n396), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT7), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n279), .B2(G20), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n202), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n412), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n411), .A2(new_n268), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n271), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n259), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n273), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(new_n259), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n377), .B1(G232), .B2(new_n299), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n301), .A2(G1698), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G223), .B2(G1698), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n400), .A2(new_n428), .B1(new_n276), .B2(new_n221), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n298), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G169), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n306), .B2(new_n431), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT80), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n432), .B(KEYINPUT80), .C1(new_n306), .C2(new_n431), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n425), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT18), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT81), .ZN(new_n440));
  INV_X1    g0240(.A(G190), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n426), .A2(new_n430), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(G200), .B1(new_n426), .B2(new_n430), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n431), .A2(new_n311), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n426), .A2(new_n430), .A3(new_n441), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(KEYINPUT81), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n419), .A2(new_n448), .A3(new_n424), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n419), .A2(new_n448), .A3(KEYINPUT17), .A4(new_n424), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n425), .A2(new_n453), .A3(new_n437), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n439), .A2(new_n451), .A3(new_n452), .A4(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n394), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n267), .A2(new_n231), .B1(G20), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n232), .C1(G33), .C2(new_n226), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT20), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(KEYINPUT87), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n463), .A2(KEYINPUT87), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n459), .A2(KEYINPUT87), .A3(new_n461), .A4(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n420), .A2(new_n458), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n270), .A2(G33), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n314), .A2(new_n271), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n467), .B(new_n468), .C1(new_n470), .C2(new_n458), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n295), .A2(G1), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G270), .A3(new_n278), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n473), .A2(new_n278), .A3(G274), .A4(new_n474), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n397), .A2(new_n399), .A3(new_n285), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(G257), .A3(new_n289), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n276), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n286), .A2(G33), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT85), .ZN(new_n485));
  AND2_X1   g0285(.A1(G264), .A2(G1698), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n397), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n288), .A2(G303), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n397), .A2(new_n399), .A3(new_n285), .A4(new_n486), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT85), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n481), .A2(new_n487), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n491), .A2(KEYINPUT86), .A3(new_n298), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT86), .B1(new_n491), .B2(new_n298), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n479), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n472), .B1(new_n494), .B2(new_n441), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n487), .A2(new_n490), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n397), .A2(new_n399), .A3(new_n289), .A4(new_n285), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n488), .B1(new_n497), .B2(new_n227), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n298), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT86), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n491), .A2(KEYINPUT86), .A3(new_n298), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n478), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n311), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT88), .B1(new_n495), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n494), .A2(G200), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(G190), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT88), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .A4(new_n472), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n476), .A2(G179), .A3(new_n477), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n472), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n493), .B2(new_n492), .ZN(new_n513));
  OAI211_X1 g0313(.A(KEYINPUT21), .B(G169), .C1(new_n466), .C2(new_n471), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n503), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n472), .A2(new_n308), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT21), .B1(new_n494), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT19), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n221), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n369), .A2(new_n232), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n260), .A2(KEYINPUT19), .A3(new_n226), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n232), .A2(G68), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n524), .A2(new_n525), .B1(new_n400), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n314), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI221_X1 g0329(.A(KEYINPUT83), .B1(new_n400), .B2(new_n526), .C1(new_n524), .C2(new_n525), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n529), .A2(new_n530), .B1(new_n420), .B2(new_n339), .ZN(new_n531));
  INV_X1    g0331(.A(new_n474), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n278), .A2(new_n532), .A3(G250), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n278), .A2(G274), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n532), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G116), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n326), .A2(G1698), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(G238), .B2(G1698), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n400), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n298), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  INV_X1    g0343(.A(new_n470), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G87), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n531), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT84), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT84), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n531), .A2(new_n548), .A3(new_n543), .A4(new_n545), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n535), .B1(new_n298), .B2(new_n540), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G190), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n339), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n531), .A2(new_n554), .B1(new_n550), .B2(new_n306), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G169), .B2(new_n550), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n221), .A2(G20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n279), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT22), .ZN(new_n560));
  OR3_X1    g0360(.A1(new_n537), .A2(KEYINPUT89), .A3(G20), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT89), .B1(new_n537), .B2(G20), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n480), .A2(KEYINPUT22), .A3(new_n558), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT23), .B1(new_n232), .B2(G107), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT90), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT90), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n567), .B(KEYINPUT23), .C1(new_n232), .C2(G107), .ZN(new_n568));
  OR3_X1    g0368(.A1(new_n232), .A2(KEYINPUT23), .A3(G107), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n563), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT24), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n563), .A2(new_n564), .A3(new_n573), .A4(new_n570), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n314), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n420), .A2(KEYINPUT25), .A3(new_n331), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT25), .B1(new_n420), .B2(new_n331), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n578), .A2(new_n579), .B1(new_n470), .B2(new_n331), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n227), .A2(G1698), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G250), .B2(G1698), .ZN(new_n583));
  INV_X1    g0383(.A(G294), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n400), .A2(new_n583), .B1(new_n276), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n298), .B1(new_n474), .B2(new_n473), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n585), .A2(new_n298), .B1(new_n586), .B2(G264), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G190), .A3(new_n477), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n477), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G200), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n576), .A2(new_n581), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT4), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n497), .B2(new_n326), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n289), .A2(KEYINPUT4), .A3(G244), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n222), .B2(new_n289), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n279), .B1(G33), .B2(G283), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n298), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n475), .A2(G257), .A3(new_n278), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT82), .B1(new_n599), .B2(new_n477), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(KEYINPUT82), .A3(new_n477), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT6), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n604), .A2(new_n226), .A3(G107), .ZN(new_n605));
  XNOR2_X1  g0405(.A(G97), .B(G107), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n607), .A2(new_n232), .B1(new_n280), .B2(new_n337), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n331), .B1(new_n415), .B2(new_n416), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n268), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n271), .A2(G97), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n544), .B2(G97), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n603), .A2(new_n308), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n602), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n600), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(new_n306), .A3(new_n598), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n603), .A2(G200), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(G190), .A3(new_n598), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n610), .A2(new_n612), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n587), .A2(G179), .A3(new_n477), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n308), .B1(new_n587), .B2(new_n477), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n575), .A2(new_n580), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n591), .A2(new_n617), .A3(new_n621), .A4(new_n624), .ZN(new_n625));
  NOR4_X1   g0425(.A1(new_n457), .A2(new_n519), .A3(new_n557), .A4(new_n625), .ZN(G372));
  INV_X1    g0426(.A(new_n310), .ZN(new_n627));
  INV_X1    g0427(.A(new_n433), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n419), .B2(new_n424), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT18), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n451), .A2(new_n452), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n347), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n392), .A2(new_n365), .B1(new_n386), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n630), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n313), .A2(new_n321), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n313), .A2(new_n321), .A3(new_n322), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n627), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n557), .B2(new_n617), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT91), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n540), .A2(new_n642), .A3(new_n298), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n540), .B2(new_n298), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n536), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n308), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n529), .A2(new_n530), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n339), .A2(new_n420), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n554), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n550), .A2(new_n306), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n645), .A2(G200), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n652), .A2(new_n531), .A3(new_n545), .A4(new_n551), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(new_n651), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  INV_X1    g0455(.A(new_n617), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n641), .A2(new_n651), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n617), .A2(new_n621), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n591), .A3(new_n654), .ZN(new_n660));
  INV_X1    g0460(.A(new_n624), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n515), .B2(new_n517), .ZN(new_n663));
  INV_X1    g0463(.A(new_n514), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n501), .A2(new_n502), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n494), .A2(new_n664), .B1(new_n665), .B2(new_n512), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT21), .ZN(new_n667));
  INV_X1    g0467(.A(new_n516), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n503), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n669), .A3(KEYINPUT92), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n661), .B1(new_n663), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n660), .B1(new_n671), .B2(KEYINPUT93), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n515), .A2(new_n517), .A3(new_n662), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT92), .B1(new_n666), .B2(new_n669), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n624), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT93), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n658), .B1(new_n672), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n640), .B1(new_n457), .B2(new_n678), .ZN(G369));
  NAND3_X1  g0479(.A1(new_n270), .A2(new_n232), .A3(G13), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n472), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n663), .A2(new_n670), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n519), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n685), .B1(new_n575), .B2(new_n580), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n591), .A2(new_n624), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT94), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n661), .B2(new_n685), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n624), .A2(KEYINPUT94), .A3(new_n686), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n518), .A2(new_n685), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n697), .A2(new_n699), .B1(new_n661), .B2(new_n686), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n216), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n521), .A2(new_n221), .A3(new_n458), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n703), .A2(new_n270), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n234), .B2(new_n703), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT28), .Z(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n542), .A2(new_n511), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n615), .A3(new_n587), .A4(new_n598), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n492), .A2(new_n493), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT30), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n550), .A2(G179), .A3(new_n479), .A4(new_n587), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n603), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n665), .A3(new_n715), .ZN(new_n716));
  AND4_X1   g0516(.A1(new_n306), .A2(new_n603), .A3(new_n645), .A4(new_n589), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n712), .A2(new_n716), .B1(new_n494), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n685), .B1(new_n718), .B2(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n712), .A2(new_n716), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n494), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n720), .A2(KEYINPUT95), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n708), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n557), .A2(new_n625), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n510), .A3(new_n518), .A4(new_n686), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT30), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n715), .B1(new_n714), .B2(new_n665), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n723), .A2(new_n725), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT96), .B1(new_n678), .B2(new_n685), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n641), .A2(new_n651), .A3(new_n657), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT93), .B(new_n624), .C1(new_n673), .C2(new_n674), .ZN(new_n735));
  INV_X1    g0535(.A(new_n660), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n671), .A2(KEYINPUT93), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT96), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(new_n686), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n653), .A2(new_n651), .A3(new_n616), .A4(new_n613), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n745), .A2(KEYINPUT26), .B1(new_n555), .B2(new_n646), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n552), .A2(new_n656), .A3(new_n655), .A4(new_n556), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n515), .A2(new_n517), .A3(new_n661), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n746), .B(new_n747), .C1(new_n660), .C2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT29), .A3(new_n686), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n732), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n707), .B1(new_n751), .B2(G1), .ZN(G364));
  INV_X1    g0552(.A(new_n703), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n214), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n270), .B1(new_n754), .B2(G45), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n691), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G330), .B2(new_n689), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n702), .A2(new_n288), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G355), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G116), .B2(new_n216), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n206), .A2(G45), .A3(new_n207), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n251), .B2(G45), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n404), .A2(new_n406), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n702), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n762), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n231), .B1(G20), .B2(new_n308), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n757), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n441), .A2(G179), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n232), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n232), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n777), .A2(G294), .B1(new_n780), .B2(G303), .ZN(new_n781));
  NOR4_X1   g0581(.A1(new_n232), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n279), .B1(new_n782), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n778), .A2(new_n441), .A3(G200), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n781), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n306), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n232), .A2(new_n441), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n787), .A2(new_n311), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n232), .A2(new_n311), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n787), .A2(G190), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G322), .A2(new_n790), .B1(new_n793), .B2(G326), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n787), .A2(new_n441), .A3(new_n791), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT33), .B(G317), .Z(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n306), .A2(new_n232), .A3(G190), .A4(G200), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT97), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n786), .B(new_n797), .C1(new_n803), .C2(G311), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT98), .Z(new_n805));
  OAI21_X1  g0605(.A(new_n279), .B1(new_n779), .B2(new_n221), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n201), .A2(new_n789), .B1(new_n795), .B2(new_n202), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(G50), .C2(new_n793), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n803), .A2(G77), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n782), .A2(G159), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT32), .Z(new_n811));
  INV_X1    g0611(.A(new_n785), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n777), .A2(G97), .B1(new_n812), .B2(G107), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n808), .A2(new_n809), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n805), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n816));
  INV_X1    g0616(.A(new_n771), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n815), .B2(KEYINPUT99), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n774), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n770), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n689), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n759), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  NOR2_X1   g0623(.A1(new_n347), .A2(new_n685), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n686), .B1(new_n343), .B2(new_n345), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT101), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(KEYINPUT101), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n826), .A2(new_n352), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n824), .B1(new_n828), .B2(new_n347), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n733), .B2(new_n741), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n347), .ZN(new_n831));
  INV_X1    g0631(.A(new_n824), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n685), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n678), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT102), .B1(new_n837), .B2(new_n732), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n757), .B1(new_n837), .B2(new_n732), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT102), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(new_n731), .C1(new_n830), .C2(new_n836), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n817), .A2(new_n769), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n757), .B1(G77), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G303), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n784), .A2(new_n795), .B1(new_n792), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G294), .B2(new_n790), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n785), .A2(new_n221), .B1(new_n779), .B2(new_n331), .ZN(new_n848));
  INV_X1    g0648(.A(new_n782), .ZN(new_n849));
  INV_X1    g0649(.A(G311), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n288), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(G97), .C2(new_n777), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n847), .B(new_n852), .C1(new_n458), .C2(new_n802), .ZN(new_n853));
  XNOR2_X1  g0653(.A(KEYINPUT100), .B(G143), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G137), .A2(new_n793), .B1(new_n790), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(G150), .ZN(new_n856));
  INV_X1    g0656(.A(G159), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n855), .B1(new_n856), .B2(new_n795), .C1(new_n802), .C2(new_n857), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT34), .Z(new_n859));
  NOR2_X1   g0659(.A1(new_n785), .A2(new_n202), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G50), .B2(new_n780), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n777), .A2(G58), .B1(G132), .B2(new_n782), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(new_n765), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n853), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n844), .B1(new_n864), .B2(new_n771), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n769), .B2(new_n829), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n842), .A2(new_n866), .ZN(G384));
  NOR2_X1   g0667(.A1(new_n754), .A2(new_n270), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT95), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n728), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n720), .A2(KEYINPUT95), .A3(new_n721), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(KEYINPUT31), .A3(new_n685), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n723), .A2(new_n725), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n365), .A2(new_n685), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n393), .A2(new_n386), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n386), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n365), .B(new_n685), .C1(new_n392), .C2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n833), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n411), .A2(new_n268), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n402), .A2(new_n408), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT79), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n402), .A2(new_n403), .A3(new_n408), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT16), .B1(new_n885), .B2(new_n396), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n424), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n683), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n425), .A2(new_n453), .A3(new_n437), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n453), .B1(new_n425), .B2(new_n437), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n889), .B1(new_n892), .B2(new_n631), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n887), .A2(new_n433), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n889), .A2(new_n894), .A3(new_n449), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n683), .B1(new_n419), .B2(new_n424), .ZN(new_n896));
  INV_X1    g0696(.A(new_n425), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n448), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT37), .B1(new_n425), .B2(new_n437), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n895), .A2(KEYINPUT37), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n880), .B1(new_n893), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n413), .B1(new_n883), .B2(new_n884), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n314), .B1(new_n902), .B2(KEYINPUT16), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n396), .B1(new_n409), .B2(new_n410), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n412), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n423), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n449), .B1(new_n906), .B2(new_n628), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n683), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n898), .A2(new_n899), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n455), .A2(new_n908), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n901), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n879), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n873), .A2(new_n878), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n916), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n425), .A2(new_n888), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n630), .B2(new_n631), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n919), .B(new_n449), .C1(new_n897), .C2(new_n628), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n921), .A2(KEYINPUT37), .B1(new_n898), .B2(new_n899), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n880), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n913), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n915), .A2(new_n916), .B1(new_n918), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n456), .A3(new_n873), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(G330), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n925), .B1(new_n456), .B2(new_n873), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT103), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n456), .A2(new_n750), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n744), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n640), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n924), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n393), .A2(new_n685), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n913), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n832), .B1(new_n678), .B2(new_n835), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n875), .A2(new_n877), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n914), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n630), .A2(new_n888), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n939), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n934), .B(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n868), .B1(new_n930), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n930), .B2(new_n945), .ZN(new_n947));
  INV_X1    g0747(.A(new_n607), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT35), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(KEYINPUT35), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n949), .A2(G116), .A3(new_n233), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n234), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(G50), .B2(new_n202), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n214), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n952), .A3(new_n955), .ZN(G367));
  AOI21_X1  g0756(.A(new_n686), .B1(new_n531), .B2(new_n545), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT104), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n651), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n654), .B2(new_n958), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n960), .A2(new_n770), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n766), .A2(new_n244), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(new_n772), .C1(new_n216), .C2(new_n339), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n856), .A2(new_n789), .B1(new_n795), .B2(new_n857), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n793), .B2(new_n854), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n776), .A2(new_n202), .B1(new_n785), .B2(new_n280), .ZN(new_n966));
  INV_X1    g0766(.A(G137), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n279), .B1(new_n849), .B2(new_n967), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n966), .B(new_n968), .C1(G58), .C2(new_n780), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n965), .B(new_n969), .C1(new_n207), .C2(new_n802), .ZN(new_n970));
  XOR2_X1   g0770(.A(KEYINPUT111), .B(G317), .Z(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n782), .A2(new_n972), .B1(new_n812), .B2(G97), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n331), .B2(new_n776), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n845), .A2(new_n789), .B1(new_n792), .B2(new_n850), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n974), .A2(new_n765), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n802), .B2(new_n784), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT46), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n779), .B2(new_n458), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n978), .B(new_n980), .C1(new_n584), .C2(new_n795), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT110), .Z(new_n982));
  OAI21_X1  g0782(.A(new_n970), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT47), .Z(new_n984));
  OAI211_X1 g0784(.A(new_n757), .B(new_n963), .C1(new_n984), .C2(new_n817), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n961), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n755), .B(KEYINPUT109), .Z(new_n988));
  AND3_X1   g0788(.A1(new_n689), .A2(KEYINPUT108), .A3(G330), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n697), .B(new_n699), .Z(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(new_n989), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n991), .B1(new_n993), .B2(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n751), .ZN(new_n995));
  INV_X1    g0795(.A(new_n698), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n617), .A2(new_n686), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT105), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n659), .B1(new_n620), .B2(new_n686), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n700), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT44), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n700), .A2(new_n1001), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT107), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT107), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n700), .A2(new_n1001), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT45), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n996), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1010), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1012), .A2(new_n698), .A3(new_n1003), .A4(new_n1008), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n751), .B1(new_n995), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n703), .B(KEYINPUT41), .Z(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n988), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1001), .A2(new_n697), .A3(new_n699), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT42), .Z(new_n1020));
  AOI21_X1  g0820(.A(new_n656), .B1(new_n1001), .B2(new_n661), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n685), .B1(new_n1021), .B2(KEYINPUT106), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(KEYINPUT106), .B2(new_n1021), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT43), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n960), .A2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n960), .A2(new_n1025), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1020), .A2(new_n1023), .A3(new_n1025), .A4(new_n960), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1001), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n698), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1030), .B(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n987), .B1(new_n1018), .B2(new_n1034), .ZN(G387));
  NAND2_X1  g0835(.A1(new_n994), .A2(new_n988), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n766), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n241), .B2(G45), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n704), .B2(new_n760), .ZN(new_n1039));
  AOI211_X1 g0839(.A(G45), .B(new_n704), .C1(G68), .C2(G77), .ZN(new_n1040));
  OR3_X1    g0840(.A1(new_n336), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT50), .B1(new_n336), .B2(G50), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1039), .A2(new_n1043), .B1(G107), .B2(new_n216), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n756), .B1(new_n1044), .B2(new_n772), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n777), .A2(new_n553), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n780), .A2(G77), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n765), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n849), .A2(new_n856), .B1(new_n226), .B2(new_n785), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n795), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n259), .A2(new_n1052), .B1(new_n793), .B2(G159), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n207), .C2(new_n789), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G68), .B2(new_n803), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT112), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G311), .A2(new_n1052), .B1(new_n790), .B2(new_n972), .ZN(new_n1057));
  INV_X1    g0857(.A(G322), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n792), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n803), .B2(G303), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT48), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(KEYINPUT48), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n777), .A2(G283), .B1(new_n780), .B2(G294), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT49), .Z(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n782), .A2(G326), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1049), .B(new_n1067), .C1(new_n458), .C2(new_n785), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1065), .B2(KEYINPUT113), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1056), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1045), .B1(new_n697), .B2(new_n820), .C1(new_n1070), .C2(new_n817), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n995), .A2(new_n703), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n994), .A2(new_n751), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1036), .B(new_n1071), .C1(new_n1072), .C2(new_n1073), .ZN(G393));
  INV_X1    g0874(.A(new_n1014), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n988), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n772), .B1(new_n226), .B2(new_n216), .C1(new_n1037), .C2(new_n248), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n757), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n288), .B1(new_n785), .B2(new_n331), .C1(new_n849), .C2(new_n1058), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n776), .A2(new_n458), .B1(new_n779), .B2(new_n784), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n845), .B2(new_n795), .ZN(new_n1082));
  INV_X1    g0882(.A(G317), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n850), .A2(new_n789), .B1(new_n792), .B2(new_n1083), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1085));
  AOI21_X1  g0885(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n584), .B2(new_n802), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n812), .A2(G87), .B1(new_n782), .B2(new_n854), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n202), .B2(new_n779), .C1(new_n280), .C2(new_n776), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G50), .B2(new_n1052), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n765), .C1(new_n336), .C2(new_n802), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n856), .A2(new_n792), .B1(new_n789), .B2(new_n857), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  OAI21_X1  g0893(.A(new_n1087), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1078), .B1(new_n1094), .B2(new_n771), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1001), .B2(new_n820), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n995), .A2(new_n1014), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n703), .B1(new_n995), .B2(new_n1014), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1076), .B(new_n1096), .C1(new_n1097), .C2(new_n1098), .ZN(G390));
  NAND3_X1  g0899(.A1(new_n749), .A2(new_n686), .A3(new_n829), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n832), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n941), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n937), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n924), .A3(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n730), .A2(G330), .A3(new_n829), .A4(new_n941), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n913), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT39), .B1(new_n923), .B2(new_n913), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1104), .B(new_n1105), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n936), .A2(new_n938), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n824), .B1(new_n739), .B2(new_n834), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n941), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1103), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n937), .B1(new_n923), .B2(new_n913), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1111), .A2(new_n1114), .B1(new_n1102), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n873), .A2(G330), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n878), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1110), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n873), .A2(G330), .A3(new_n829), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n1113), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1101), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n1105), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n730), .A2(G330), .A3(new_n829), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1117), .A2(new_n878), .B1(new_n1124), .B2(new_n1113), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n1112), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1117), .A2(new_n456), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1126), .A2(new_n933), .A3(new_n640), .A4(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n753), .B1(new_n1119), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1113), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1118), .A2(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1105), .A2(new_n1122), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1131), .A2(new_n940), .B1(new_n1132), .B2(new_n1121), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT29), .B1(new_n733), .B2(new_n741), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n640), .B(new_n1127), .C1(new_n1134), .C2(new_n931), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1104), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n878), .A3(new_n1117), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1138), .A3(new_n1110), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1129), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT115), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT115), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1129), .A2(new_n1142), .A3(new_n1139), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1110), .B(new_n988), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n757), .B1(new_n259), .B2(new_n843), .ZN(new_n1146));
  INV_X1    g0946(.A(G128), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n779), .A2(new_n856), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT53), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n792), .A2(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n279), .B1(new_n776), .B2(new_n857), .C1(new_n1151), .C2(new_n849), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(G50), .C2(new_n812), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n967), .B2(new_n795), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G132), .B2(new_n790), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1153), .B(new_n1156), .C1(new_n802), .C2(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n288), .B1(new_n779), .B2(new_n221), .C1(new_n849), .C2(new_n584), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n860), .B(new_n1159), .C1(G77), .C2(new_n777), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n331), .A2(new_n795), .B1(new_n789), .B2(new_n458), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G283), .B2(new_n793), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(new_n226), .C2(new_n802), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1146), .B1(new_n1164), .B2(new_n771), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1108), .B2(new_n769), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1145), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT116), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT116), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1145), .A2(new_n1169), .A3(new_n1166), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1144), .A2(new_n1172), .ZN(G378));
  NAND3_X1  g0973(.A1(new_n879), .A2(new_n924), .A3(KEYINPUT40), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n917), .B1(new_n913), .B2(new_n901), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(G330), .C1(new_n1175), .C2(KEYINPUT40), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1177));
  NAND2_X1  g0977(.A1(new_n325), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1177), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n639), .A2(new_n310), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n275), .A2(new_n888), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1181), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1181), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1185), .B1(new_n1190), .B2(new_n1182), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1176), .A2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n939), .A2(new_n942), .A3(new_n943), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n915), .A2(new_n916), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(G330), .A4(new_n1174), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1193), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1194), .B1(new_n1197), .B2(new_n1193), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1195), .A2(new_n768), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n757), .B1(G50), .B2(new_n843), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n777), .A2(G150), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n779), .B2(new_n1157), .C1(new_n1151), .C2(new_n792), .ZN(new_n1204));
  INV_X1    g1004(.A(G132), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1147), .A2(new_n789), .B1(new_n795), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n803), .C2(G137), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT59), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n812), .A2(G159), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n782), .C2(G124), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n792), .A2(new_n458), .B1(new_n776), .B2(new_n202), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT117), .Z(new_n1215));
  OAI22_X1  g1015(.A1(new_n226), .A2(new_n795), .B1(new_n789), .B2(new_n331), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G41), .B1(new_n782), .B2(G283), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1047), .B(new_n1217), .C1(new_n201), .C2(new_n785), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1216), .A2(new_n1218), .A3(new_n765), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1215), .B(new_n1219), .C1(new_n802), .C2(new_n339), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT58), .ZN(new_n1221));
  AOI21_X1  g1021(.A(G41), .B1(new_n765), .B2(G33), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1213), .B(new_n1221), .C1(G50), .C2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1202), .B1(new_n1223), .B2(new_n771), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1200), .A2(new_n988), .B1(new_n1201), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1135), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1119), .B2(new_n1133), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1195), .B1(new_n925), .B2(G330), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1176), .A2(new_n1192), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n944), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1193), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(KEYINPUT57), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n703), .B1(new_n1228), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1227), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1225), .B1(new_n1234), .B2(new_n1235), .ZN(G375));
  OAI21_X1  g1036(.A(new_n757), .B1(G68), .B2(new_n843), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n802), .A2(new_n856), .B1(new_n207), .B2(new_n776), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT122), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n765), .B1(new_n201), .B2(new_n785), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT123), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G132), .A2(new_n793), .B1(new_n790), .B2(G137), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n780), .A2(G159), .B1(G128), .B2(new_n782), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(new_n795), .C2(new_n1157), .ZN(new_n1244));
  OR3_X1    g1044(.A1(new_n1239), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n803), .A2(G107), .B1(G116), .B2(new_n1052), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1246), .A2(KEYINPUT120), .B1(G294), .B2(new_n793), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(KEYINPUT120), .B2(new_n1246), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT121), .Z(new_n1249));
  OAI21_X1  g1049(.A(new_n288), .B1(new_n849), .B2(new_n845), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1046), .B1(new_n226), .B2(new_n779), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(G77), .C2(new_n812), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n784), .B2(new_n789), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1245), .B1(new_n1249), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1237), .B1(new_n1254), .B2(new_n771), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n769), .B2(new_n941), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n988), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1256), .B1(new_n1133), .B2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT124), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1128), .A2(new_n1017), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(G381));
  NOR3_X1   g1062(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(G390), .A2(G384), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n751), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n1075), .B2(new_n994), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1257), .B1(new_n1267), .B2(new_n1016), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1034), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n986), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1201), .A2(new_n1224), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(new_n1257), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT57), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1198), .A2(new_n1199), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n753), .B1(new_n1275), .B2(new_n1227), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1228), .B2(new_n1272), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1273), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1167), .B1(new_n1129), .B2(new_n1139), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1265), .A2(new_n1270), .A3(new_n1278), .A4(new_n1279), .ZN(G407));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n684), .A3(new_n1279), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(G213), .A3(new_n1281), .ZN(G409));
  INV_X1    g1082(.A(G390), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G390), .B(new_n987), .C1(new_n1018), .C2(new_n1034), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1270), .B2(G390), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(G393), .B(new_n822), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1286), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1284), .A2(new_n1289), .A3(new_n1285), .A4(new_n1287), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1200), .A2(new_n1017), .A3(new_n1227), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1225), .A2(new_n1294), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1278), .A2(G378), .B1(new_n1279), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G213), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(G343), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1258), .B(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1133), .A2(new_n1135), .A3(KEYINPUT60), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n703), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1128), .A2(KEYINPUT60), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1260), .B2(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(KEYINPUT126), .B(G384), .C1(new_n1300), .C2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1260), .B1(new_n1136), .B2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n703), .A3(new_n1301), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n842), .A2(new_n1310), .A3(new_n866), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1306), .A2(new_n1309), .A3(new_n1259), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1305), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT62), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1296), .A2(new_n1298), .A3(new_n1314), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1228), .A2(new_n1272), .A3(new_n1016), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1279), .B1(new_n1316), .B2(new_n1273), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1171), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(G375), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1317), .B(KEYINPUT125), .C1(G375), .C2(new_n1318), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1298), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1321), .A2(new_n1313), .A3(new_n1322), .A4(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT62), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1315), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1298), .A2(G2897), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1313), .B(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT61), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1293), .B1(new_n1326), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1324), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1328), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1319), .A2(KEYINPUT63), .A3(new_n1313), .A4(new_n1323), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1293), .A2(KEYINPUT61), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1334), .A2(new_n1336), .A3(new_n1337), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1332), .A2(new_n1339), .ZN(G405));
  INV_X1    g1140(.A(new_n1313), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1293), .A2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1291), .A2(new_n1313), .A3(new_n1292), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(G375), .A2(new_n1318), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1345), .B1(G375), .B2(new_n1279), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1344), .B(new_n1346), .ZN(G402));
endmodule


