//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n207), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT0), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT67), .Z(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT66), .B(G77), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n220), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT65), .B(G238), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G68), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n214), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n218), .B1(new_n217), .B2(new_n216), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G200), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  INV_X1    g0051(.A(G223), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1698), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT75), .ZN(new_n257));
  OR2_X1    g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT75), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(new_n261), .A3(new_n253), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g0063(.A(G226), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G87), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n251), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n251), .A2(new_n269), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(new_n273), .B2(G232), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n249), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G190), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n266), .B1(new_n262), .B2(new_n257), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n277), .B(new_n274), .C1(new_n278), .C2(new_n251), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n206), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT69), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G1), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G20), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT69), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n281), .A2(new_n287), .A3(new_n206), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n283), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n212), .B2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n284), .A2(new_n207), .A3(G1), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT16), .ZN(new_n297));
  INV_X1    g0097(.A(G68), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n258), .A2(new_n207), .A3(new_n259), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT7), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n254), .A2(new_n255), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n298), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(G58), .B(G68), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G20), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT70), .ZN(new_n307));
  INV_X1    g0107(.A(G33), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n207), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G159), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n306), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n297), .B1(new_n304), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT7), .B1(new_n302), .B2(new_n207), .ZN(new_n316));
  NOR4_X1   g0116(.A1(new_n254), .A2(new_n255), .A3(new_n300), .A4(G20), .ZN(new_n317));
  OAI21_X1  g0117(.A(G68), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n311), .A2(G159), .B1(new_n305), .B2(G20), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(KEYINPUT16), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n315), .A2(new_n320), .A3(new_n282), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n280), .A2(new_n296), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT17), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n282), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n318), .A2(new_n319), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n297), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n295), .B1(new_n327), .B2(new_n320), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT17), .A3(new_n280), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n268), .B2(new_n275), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n333), .B(new_n274), .C1(new_n278), .C2(new_n251), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n321), .A2(new_n296), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(KEYINPUT18), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT18), .B1(new_n335), .B2(new_n336), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT76), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n332), .A2(new_n334), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT18), .ZN(new_n342));
  NOR4_X1   g0142(.A1(new_n328), .A2(new_n341), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n330), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G1698), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n260), .A2(G226), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n260), .A2(G232), .A3(G1698), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n206), .B1(G33), .B2(G41), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT13), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n271), .B1(new_n273), .B2(G238), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(new_n352), .B2(new_n354), .ZN(new_n356));
  OAI21_X1  g0156(.A(G169), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT14), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n352), .A2(new_n354), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT13), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(G169), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(G179), .A3(new_n361), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n358), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n285), .A2(G20), .A3(new_n298), .ZN(new_n367));
  XOR2_X1   g0167(.A(new_n367), .B(KEYINPUT12), .Z(new_n368));
  NOR2_X1   g0168(.A1(new_n293), .A2(new_n282), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n298), .B1(new_n212), .B2(G20), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n207), .A2(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n202), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(G20), .B2(new_n298), .ZN(new_n374));
  INV_X1    g0174(.A(G50), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n312), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n283), .A2(new_n288), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT11), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(KEYINPUT11), .A3(new_n377), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n371), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n366), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n362), .A2(new_n249), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n360), .A2(new_n277), .A3(new_n361), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n312), .A2(new_n290), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n223), .A2(new_n207), .B1(new_n391), .B2(new_n372), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n282), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT71), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n395), .B(new_n282), .C1(new_n390), .C2(new_n392), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n202), .B1(new_n212), .B2(G20), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n369), .A2(new_n398), .B1(new_n223), .B2(new_n293), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n271), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n272), .B2(new_n221), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n260), .A2(new_n225), .A3(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n260), .A2(G232), .A3(new_n346), .ZN(new_n404));
  INV_X1    g0204(.A(G107), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n403), .B(new_n404), .C1(new_n405), .C2(new_n260), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n402), .B1(new_n406), .B2(new_n351), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G179), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n331), .B2(new_n407), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n400), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n407), .A2(new_n277), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n407), .A2(G200), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n397), .B(new_n399), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  AND4_X1   g0214(.A1(new_n345), .A2(new_n385), .A3(new_n389), .A4(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n252), .A2(new_n346), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n346), .A2(G222), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n260), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n302), .A2(new_n222), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n251), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G226), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n401), .B1(new_n272), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G179), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n331), .B2(new_n423), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n289), .B(G50), .C1(G1), .C2(new_n207), .ZN(new_n426));
  INV_X1    g0226(.A(G150), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n312), .A2(new_n427), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n290), .A2(new_n372), .B1(new_n207), .B2(new_n201), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n377), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n293), .A2(new_n375), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n423), .A2(G190), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n249), .B2(new_n423), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT72), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n426), .A2(new_n430), .A3(KEYINPUT72), .A4(new_n431), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT9), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n436), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT10), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(KEYINPUT9), .A3(new_n439), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT73), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n442), .A2(KEYINPUT73), .A3(new_n443), .A4(new_n444), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n442), .A2(new_n444), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT10), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n434), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n415), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n346), .A2(G244), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n258), .B2(new_n259), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT4), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT77), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n454), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n221), .A2(G1698), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n458), .C1(new_n255), .C2(new_n254), .ZN(new_n461));
  OAI211_X1 g0261(.A(G250), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n351), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G41), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n212), .B(G45), .C1(new_n465), .C2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G41), .ZN(new_n468));
  OAI211_X1 g0268(.A(G257), .B(new_n251), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT78), .B1(new_n467), .B2(G41), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT78), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(new_n465), .A3(KEYINPUT5), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n467), .A2(G41), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(new_n212), .A3(G45), .A4(G274), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(G169), .B1(new_n464), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n286), .A2(G97), .ZN(new_n480));
  OAI21_X1  g0280(.A(G107), .B1(new_n316), .B2(new_n317), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n202), .B1(new_n309), .B2(new_n310), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  AND2_X1   g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  NOR2_X1   g0284(.A1(G97), .A2(G107), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n405), .A2(KEYINPUT6), .A3(G97), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n482), .B1(new_n488), .B2(G20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n481), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n480), .B1(new_n490), .B2(new_n282), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n212), .A2(G33), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n283), .A2(new_n286), .A3(new_n288), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G97), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n479), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n464), .A2(new_n333), .A3(new_n478), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT80), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n464), .A2(new_n478), .A3(KEYINPUT80), .A4(new_n333), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT81), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n496), .B2(new_n501), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n464), .A2(G190), .A3(new_n478), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n491), .A2(new_n505), .A3(new_n495), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT79), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n464), .A2(new_n478), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(G200), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n507), .A3(G200), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n506), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n503), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT20), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n207), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G97), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n454), .B1(new_n517), .B2(G33), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n518), .B2(new_n207), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n514), .B1(new_n519), .B2(new_n325), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n308), .A2(G97), .ZN(new_n521));
  AOI21_X1  g0321(.A(G20), .B1(new_n521), .B2(new_n454), .ZN(new_n522));
  OAI211_X1 g0322(.A(KEYINPUT20), .B(new_n282), .C1(new_n522), .C2(new_n516), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n515), .B1(new_n212), .B2(G33), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n369), .A2(new_n525), .B1(new_n515), .B2(new_n293), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n474), .A2(new_n476), .ZN(new_n527));
  OAI211_X1 g0327(.A(G270), .B(new_n251), .C1(new_n466), .C2(new_n468), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n346), .A2(G257), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G264), .A2(G1698), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n258), .A2(new_n259), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G303), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n254), .A2(new_n255), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n351), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT85), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G257), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G1698), .ZN(new_n539));
  AND2_X1   g0339(.A1(G264), .A2(G1698), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n539), .A2(new_n540), .B1(new_n254), .B2(new_n255), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n258), .A2(G303), .A3(new_n259), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(KEYINPUT85), .A3(new_n351), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n529), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  INV_X1    g0346(.A(new_n528), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(new_n477), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT85), .B1(new_n543), .B2(new_n351), .ZN(new_n549));
  AOI211_X1 g0349(.A(new_n536), .B(new_n251), .C1(new_n541), .C2(new_n542), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n524), .B(new_n526), .C1(new_n546), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n524), .A2(new_n526), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n545), .A2(G179), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n551), .A2(new_n554), .A3(KEYINPUT21), .A4(G169), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n551), .A2(G169), .A3(new_n554), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT86), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n553), .B(new_n557), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n308), .A2(new_n515), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n207), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT23), .B1(new_n405), .B2(G20), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n568), .A2(new_n207), .A3(G107), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n566), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n207), .B(G87), .C1(new_n254), .C2(new_n255), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT22), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n260), .A2(new_n573), .A3(new_n207), .A4(G87), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n325), .B1(new_n575), .B2(KEYINPUT24), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT24), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n572), .A2(new_n574), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(new_n570), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n285), .A2(G20), .A3(new_n405), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n581), .B(KEYINPUT25), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n494), .B2(G107), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT87), .ZN(new_n585));
  INV_X1    g0385(.A(G250), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(G1698), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G257), .A2(G1698), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n587), .A2(new_n589), .B1(new_n254), .B2(new_n255), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G294), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n251), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(G264), .B(new_n251), .C1(new_n466), .C2(new_n468), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n585), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n588), .B1(new_n586), .B2(G1698), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n260), .A2(new_n596), .B1(G33), .B2(G294), .ZN(new_n597));
  OAI211_X1 g0397(.A(KEYINPUT87), .B(new_n593), .C1(new_n597), .C2(new_n251), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n527), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n592), .A2(new_n594), .A3(new_n477), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n599), .A2(new_n333), .B1(new_n331), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n584), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n584), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n249), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT88), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n599), .A2(KEYINPUT88), .A3(new_n249), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n600), .A2(new_n277), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n603), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G45), .ZN(new_n612));
  OAI21_X1  g0412(.A(G250), .B1(new_n612), .B2(G1), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n212), .A2(G45), .A3(G274), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n251), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n346), .A2(G238), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G244), .A2(G1698), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n565), .B1(new_n260), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n616), .B1(new_n620), .B2(new_n251), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G169), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n333), .B2(new_n621), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT19), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n207), .B1(new_n349), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(G87), .A2(G97), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n405), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n207), .B(G68), .C1(new_n254), .C2(new_n255), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n624), .B1(new_n349), .B2(G20), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n282), .B1(new_n293), .B2(new_n391), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n391), .B2(new_n493), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n351), .B1(new_n613), .B2(new_n614), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n260), .A2(new_n619), .ZN(new_n636));
  INV_X1    g0436(.A(new_n565), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n635), .B1(new_n638), .B2(new_n351), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(KEYINPUT83), .A3(G190), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT83), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n621), .B2(G200), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n621), .A2(new_n277), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT82), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n289), .A2(new_n645), .A3(G87), .A4(new_n492), .ZN(new_n646));
  INV_X1    g0446(.A(G87), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT82), .B1(new_n493), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n632), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n634), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n634), .B(KEYINPUT84), .C1(new_n644), .C2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n513), .A2(new_n564), .A3(new_n611), .A4(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n453), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g0456(.A(new_n656), .B(KEYINPUT89), .Z(G372));
  OAI21_X1  g0457(.A(new_n342), .B1(new_n328), .B2(new_n341), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n337), .ZN(new_n659));
  INV_X1    g0459(.A(new_n410), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n389), .A2(new_n660), .B1(new_n366), .B2(new_n384), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n661), .B2(new_n330), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n449), .A2(new_n451), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n434), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n653), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n646), .A2(new_n632), .A3(new_n648), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n258), .A2(new_n259), .B1(new_n617), .B2(new_n618), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n351), .B1(new_n667), .B2(new_n565), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n249), .B1(new_n668), .B2(new_n616), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n669), .A2(new_n641), .B1(new_n277), .B2(new_n621), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n666), .A2(new_n670), .A3(new_n640), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT84), .B1(new_n671), .B2(new_n634), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n503), .A2(new_n504), .B1(new_n665), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT26), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n503), .A2(new_n504), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n650), .B1(new_n610), .B2(new_n604), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n490), .A2(new_n282), .ZN(new_n677));
  INV_X1    g0477(.A(new_n480), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n495), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n511), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n680), .B(new_n505), .C1(new_n681), .C2(new_n509), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n557), .B(new_n602), .C1(new_n561), .C2(new_n562), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n675), .A2(new_n676), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n671), .A2(new_n496), .A3(new_n501), .A4(new_n634), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(KEYINPUT26), .ZN(new_n686));
  INV_X1    g0486(.A(new_n634), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n674), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n664), .B1(new_n453), .B2(new_n690), .ZN(G369));
  NAND2_X1  g0491(.A1(new_n285), .A2(new_n207), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT90), .ZN(new_n694));
  INV_X1    g0494(.A(G213), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n692), .B2(KEYINPUT27), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n694), .A2(G343), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n554), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n563), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n557), .B1(new_n561), .B2(new_n562), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n584), .A2(new_n697), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n611), .A2(new_n704), .B1(new_n603), .B2(new_n697), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n697), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n603), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n700), .A2(new_n708), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n608), .A2(new_n609), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT88), .B1(new_n599), .B2(new_n249), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n604), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n602), .A3(new_n704), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n709), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n709), .C1(new_n710), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n707), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT92), .Z(G399));
  INV_X1    g0521(.A(new_n215), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G1), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n626), .A2(new_n405), .A3(new_n515), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n725), .A2(new_n726), .B1(new_n210), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n595), .A2(new_n598), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n729), .A2(new_n639), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n551), .A2(new_n333), .ZN(new_n731));
  INV_X1    g0531(.A(new_n508), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n732), .A3(new_n639), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n545), .A2(G179), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n639), .A2(G179), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n599), .A2(new_n738), .A3(new_n551), .A4(new_n508), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n733), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n697), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n741), .A2(KEYINPUT31), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n655), .B2(new_n697), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n741), .A2(KEYINPUT31), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G330), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT26), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n654), .B(new_n749), .C1(new_n504), .C2(new_n503), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n687), .B1(new_n685), .B2(KEYINPUT26), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n684), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(KEYINPUT29), .A3(new_n708), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT93), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n752), .A2(new_n755), .A3(KEYINPUT29), .A4(new_n708), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT29), .B1(new_n689), .B2(new_n708), .ZN(new_n758));
  OAI211_X1 g0558(.A(KEYINPUT94), .B(new_n748), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT94), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n758), .B1(new_n754), .B2(new_n756), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n761), .B2(new_n747), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n728), .B1(new_n763), .B2(G1), .ZN(G364));
  NOR2_X1   g0564(.A1(new_n284), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n725), .B1(G45), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n703), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n702), .A2(G330), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n702), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n206), .B1(G20), .B2(new_n331), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n722), .A2(new_n260), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n244), .A2(new_n612), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n210), .A2(new_n612), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n722), .A2(new_n302), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G355), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G116), .B2(new_n215), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n776), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n207), .A2(new_n277), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(new_n249), .A3(G179), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n333), .A2(new_n249), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n789), .A2(new_n647), .B1(new_n791), .B2(new_n375), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n207), .A2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n794), .A2(G179), .A3(new_n249), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n792), .B1(G107), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G179), .A2(G200), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n207), .B1(new_n797), .B2(G190), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G97), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n793), .A2(new_n797), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n313), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT32), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n793), .A2(G179), .A3(new_n249), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n786), .A2(G179), .A3(new_n249), .ZN(new_n805));
  INV_X1    g0605(.A(G58), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n223), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n790), .A2(new_n793), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n302), .B(new_n807), .C1(G68), .C2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n796), .A2(new_n800), .A3(new_n803), .A4(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT33), .B(G317), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n808), .B1(new_n813), .B2(KEYINPUT97), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(KEYINPUT97), .B2(new_n813), .ZN(new_n815));
  INV_X1    g0615(.A(new_n804), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n788), .A2(G303), .B1(G311), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n805), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n795), .A2(G283), .B1(new_n818), .B2(G322), .ZN(new_n819));
  INV_X1    g0619(.A(new_n801), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n260), .B1(new_n820), .B2(G329), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n815), .A2(new_n817), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G326), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n791), .A2(new_n823), .B1(new_n798), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT96), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n811), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n775), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n785), .A2(new_n828), .A3(new_n766), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n768), .A2(new_n769), .B1(new_n774), .B2(new_n829), .ZN(G396));
  NAND2_X1  g0630(.A1(new_n689), .A2(new_n708), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n400), .A2(new_n697), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n413), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n410), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n660), .A2(new_n708), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n831), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n766), .B1(new_n838), .B2(new_n747), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n747), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n775), .A2(new_n770), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n767), .B1(new_n202), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n795), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n298), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G50), .B2(new_n788), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n806), .B2(new_n798), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n302), .B1(new_n820), .B2(G132), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(KEYINPUT99), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n791), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G137), .A2(new_n849), .B1(new_n816), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G143), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n851), .B2(new_n805), .C1(new_n427), .C2(new_n808), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT34), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n848), .B(new_n853), .C1(KEYINPUT99), .C2(new_n847), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n533), .A2(new_n791), .B1(new_n804), .B2(new_n515), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n260), .B(new_n855), .C1(G107), .C2(new_n788), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n818), .A2(G294), .B1(new_n809), .B2(G283), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n795), .A2(G87), .B1(G311), .B2(new_n820), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n856), .A2(new_n800), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT98), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n854), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n775), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n842), .B1(new_n837), .B2(new_n771), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n840), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT100), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n866), .B(new_n867), .ZN(G384));
  OAI21_X1  g0668(.A(new_n222), .B1(new_n806), .B2(new_n298), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n869), .A2(new_n210), .B1(G50), .B2(new_n298), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(G1), .A3(new_n284), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n486), .A2(new_n487), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT35), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n515), .B(new_n209), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n873), .B2(new_n872), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT36), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  INV_X1    g0678(.A(new_n377), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n326), .B2(new_n297), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n295), .B1(new_n880), .B2(new_n320), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n694), .A2(new_n696), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT101), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n315), .A2(new_n320), .A3(new_n377), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n296), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT101), .ZN(new_n886));
  INV_X1    g0686(.A(new_n882), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n340), .A2(new_n344), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n328), .A2(KEYINPUT17), .A3(new_n280), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT17), .B1(new_n328), .B2(new_n280), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n890), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n336), .A2(new_n334), .A3(new_n332), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n336), .A2(new_n887), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n896), .A2(new_n322), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n335), .A2(new_n885), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n883), .A2(new_n322), .A3(new_n901), .A4(new_n888), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n900), .B1(KEYINPUT37), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n895), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n658), .A2(KEYINPUT76), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n343), .B1(new_n906), .B2(new_n337), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n889), .B1(new_n907), .B2(new_n330), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n899), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n384), .A2(new_n697), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n385), .A2(new_n913), .A3(new_n389), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n384), .B(new_n697), .C1(new_n366), .C2(new_n388), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n836), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n654), .A2(new_n602), .A3(new_n713), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n496), .A2(new_n501), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT81), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n682), .A3(new_n920), .ZN(new_n921));
  NOR4_X1   g0721(.A1(new_n917), .A2(new_n921), .A3(new_n563), .A4(new_n697), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n741), .A2(KEYINPUT31), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n916), .B(new_n744), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n924), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT102), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n328), .A2(new_n341), .A3(new_n342), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n324), .B(new_n329), .C1(new_n928), .C2(new_n338), .ZN(new_n929));
  INV_X1    g0729(.A(new_n897), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n896), .A2(new_n322), .A3(new_n897), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT37), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n929), .A2(new_n930), .B1(new_n932), .B2(new_n899), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n927), .B1(new_n933), .B2(KEYINPUT38), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n910), .B(KEYINPUT38), .C1(new_n345), .C2(new_n890), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n932), .A2(new_n899), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n897), .B1(new_n894), .B2(new_n659), .ZN(new_n937));
  OAI211_X1 g0737(.A(KEYINPUT102), .B(new_n904), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n926), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n925), .B1(KEYINPUT40), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n453), .ZN(new_n942));
  INV_X1    g0742(.A(new_n745), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n941), .A2(new_n746), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n942), .A2(new_n943), .A3(G330), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n945), .B1(new_n949), .B2(KEYINPUT104), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT104), .B2(new_n949), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT105), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n385), .A2(new_n697), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT39), .ZN(new_n954));
  AND4_X1   g0754(.A1(new_n954), .A2(new_n934), .A3(new_n935), .A4(new_n938), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n904), .B1(new_n895), .B2(new_n903), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n956), .B2(new_n935), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n953), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n914), .A2(new_n915), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n689), .A2(new_n708), .A3(new_n837), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n961), .B2(new_n835), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n905), .B2(new_n911), .ZN(new_n963));
  INV_X1    g0763(.A(new_n659), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n882), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n958), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT103), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT39), .B1(new_n905), .B2(new_n911), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n934), .A2(new_n935), .A3(new_n938), .A4(new_n954), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n970), .A2(new_n953), .B1(new_n964), .B2(new_n882), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT103), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n972), .A3(new_n963), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n761), .A2(new_n942), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n664), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n974), .B(new_n976), .Z(new_n977));
  AND2_X1   g0777(.A1(new_n952), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT106), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n212), .B2(new_n765), .C1(new_n952), .C2(new_n977), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n878), .B1(new_n981), .B2(new_n982), .ZN(G367));
  OR2_X1    g0783(.A1(new_n778), .A2(new_n239), .ZN(new_n984));
  INV_X1    g0784(.A(new_n391), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n772), .B(new_n775), .C1(new_n722), .C2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n767), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n788), .A2(G116), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT46), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n798), .A2(new_n405), .ZN(new_n990));
  INV_X1    g0790(.A(G311), .ZN(new_n991));
  XNOR2_X1  g0791(.A(KEYINPUT108), .B(G317), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n791), .A2(new_n991), .B1(new_n801), .B2(new_n992), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n260), .B(new_n993), .C1(G97), .C2(new_n795), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n805), .A2(new_n533), .B1(new_n808), .B2(new_n824), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G283), .B2(new_n816), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n989), .A2(new_n990), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n805), .A2(new_n427), .B1(new_n791), .B2(new_n851), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n375), .A2(new_n804), .B1(new_n808), .B2(new_n313), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n799), .A2(G68), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n302), .B1(new_n788), .B2(G58), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT109), .B(G137), .Z(new_n1003));
  AOI22_X1  g0803(.A1(new_n795), .A2(new_n222), .B1(new_n820), .B2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT47), .B1(new_n997), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n997), .A2(KEYINPUT47), .A3(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n775), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n697), .A2(new_n649), .ZN(new_n1009));
  MUX2_X1   g0809(.A(new_n634), .B(new_n650), .S(new_n1009), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n987), .B1(new_n1006), .B2(new_n1008), .C1(new_n1011), .C2(new_n773), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n765), .A2(G45), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(G1), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n679), .A2(new_n697), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n919), .A2(new_n682), .A3(new_n920), .A4(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n496), .A2(new_n501), .A3(new_n697), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n716), .A2(new_n718), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT44), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT44), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n716), .A2(new_n1022), .A3(new_n718), .A4(new_n1019), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1019), .B1(new_n716), .B2(new_n718), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(KEYINPUT45), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT45), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1026), .B(new_n1019), .C1(new_n716), .C2(new_n718), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1021), .B(new_n1023), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n706), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1024), .B(KEYINPUT45), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n707), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n705), .A2(new_n710), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n714), .B2(new_n710), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(new_n703), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n763), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n723), .B(KEYINPUT41), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1014), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT107), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n710), .A2(new_n714), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n1018), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT42), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1018), .A2(new_n603), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n697), .B1(new_n1045), .B2(new_n675), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1041), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n706), .A2(new_n1018), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1051), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1012), .B1(new_n1039), .B2(new_n1054), .ZN(G387));
  INV_X1    g0855(.A(new_n1036), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n763), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n759), .A2(new_n762), .A3(new_n1036), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n723), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n789), .A2(new_n223), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G159), .B2(new_n849), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n799), .A2(new_n985), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n298), .A2(new_n804), .B1(new_n808), .B2(new_n290), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n805), .A2(new_n375), .B1(new_n801), .B2(new_n427), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n302), .B1(new_n795), .B2(G97), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1061), .A2(new_n1062), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n260), .B1(new_n795), .B2(G116), .ZN(new_n1068));
  INV_X1    g0868(.A(G283), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n789), .A2(new_n824), .B1(new_n798), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n804), .A2(new_n533), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n805), .A2(new_n992), .B1(new_n808), .B2(new_n991), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G322), .C2(new_n849), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1070), .B1(new_n1073), .B2(KEYINPUT48), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(KEYINPUT48), .B2(new_n1073), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT49), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1068), .B1(new_n823), .B2(new_n801), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1067), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT112), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n775), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n782), .A2(new_n726), .B1(new_n405), .B2(new_n722), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n236), .A2(new_n612), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n290), .A2(G50), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT50), .ZN(new_n1087));
  AOI211_X1 g0887(.A(G45), .B(new_n726), .C1(G68), .C2(G77), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n778), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT110), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1084), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT111), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n776), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1083), .A2(new_n1095), .A3(new_n766), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n705), .B2(new_n772), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1056), .B2(new_n1014), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1059), .A2(new_n1098), .ZN(G393));
  INV_X1    g0899(.A(new_n1033), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1036), .B1(new_n759), .B2(new_n762), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n724), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1032), .A2(KEYINPUT113), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT113), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1030), .A2(new_n1031), .A3(new_n1104), .A4(new_n707), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1029), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1057), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1103), .A2(new_n1029), .A3(new_n1014), .A4(new_n1105), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n776), .B1(new_n517), .B2(new_n215), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n777), .B2(new_n247), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n816), .A2(G294), .B1(new_n820), .B2(G322), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1069), .B2(new_n789), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n260), .B(new_n1113), .C1(G107), .C2(new_n795), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n808), .A2(new_n533), .B1(new_n798), .B2(new_n515), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT114), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n818), .A2(G311), .B1(new_n849), .B2(G317), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT52), .Z(new_n1120));
  NAND4_X1  g0920(.A1(new_n1114), .A2(new_n1117), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n805), .A2(new_n313), .B1(new_n791), .B2(new_n427), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT51), .Z(new_n1123));
  NOR2_X1   g0923(.A1(new_n801), .A2(new_n851), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n290), .A2(new_n804), .B1(new_n808), .B2(new_n375), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(G68), .C2(new_n788), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n799), .A2(G77), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n302), .B1(new_n795), .B2(G87), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1121), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n767), .B(new_n1111), .C1(new_n1130), .C2(new_n775), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1018), .B2(new_n773), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1108), .A2(new_n1109), .A3(new_n1132), .ZN(G390));
  OAI211_X1 g0933(.A(new_n968), .B(new_n969), .C1(new_n962), .C2(new_n953), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n752), .A2(new_n708), .A3(new_n834), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n835), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n959), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n953), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n939), .A3(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n743), .A2(G330), .A3(new_n744), .A4(new_n916), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1134), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n975), .A2(new_n664), .A3(new_n948), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n743), .A2(G330), .A3(new_n744), .A4(new_n837), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n960), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n1136), .A3(new_n1140), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n926), .A2(G330), .B1(new_n1143), .B2(new_n960), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n961), .A2(new_n835), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT115), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1140), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(KEYINPUT115), .B(new_n1140), .C1(new_n1134), .C2(new_n1139), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1141), .B(new_n1149), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT116), .B1(new_n1156), .B2(new_n724), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT116), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1158), .A3(new_n723), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1141), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1149), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n968), .A2(new_n770), .A3(new_n969), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n818), .A2(G116), .B1(new_n809), .B2(G107), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n517), .B2(new_n804), .C1(new_n1069), .C2(new_n791), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n844), .B(new_n1166), .C1(G294), .C2(new_n820), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n260), .B1(new_n788), .B2(G87), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT117), .Z(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(new_n1127), .A3(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n843), .A2(new_n375), .B1(new_n804), .B2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n302), .B(new_n1172), .C1(G132), .C2(new_n818), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n799), .A2(G159), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n788), .A2(G150), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT53), .Z(new_n1176));
  INV_X1    g0976(.A(G128), .ZN(new_n1177));
  INV_X1    g0977(.A(G125), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n791), .A2(new_n1177), .B1(new_n801), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n809), .B2(new_n1003), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .A4(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n864), .B1(new_n1170), .B2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n767), .B(new_n1182), .C1(new_n290), .C2(new_n841), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT118), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1164), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1014), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1185), .B1(new_n1160), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1163), .A2(new_n1188), .ZN(G378));
  NAND2_X1  g0989(.A1(new_n440), .A2(new_n887), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n452), .B(new_n1190), .Z(new_n1191));
  XOR2_X1   g0991(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n967), .A2(new_n973), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n967), .B2(new_n973), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n946), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1142), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1155), .A2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1191), .B(new_n1192), .Z(new_n1199));
  AOI21_X1  g0999(.A(new_n972), .B1(new_n971), .B2(new_n963), .ZN(new_n1200));
  AND4_X1   g1000(.A1(new_n972), .A2(new_n958), .A3(new_n963), .A4(new_n965), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n967), .A2(new_n973), .A3(new_n1193), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n947), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1196), .A2(new_n1198), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT57), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1196), .A2(new_n1198), .A3(new_n1207), .A4(new_n1204), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n724), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1196), .A2(new_n1014), .A3(new_n1204), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n767), .B1(new_n375), .B2(new_n841), .ZN(new_n1211));
  INV_X1    g1011(.A(G137), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1178), .A2(new_n791), .B1(new_n804), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1171), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n788), .A2(new_n1214), .B1(G132), .B2(new_n809), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1177), .B2(new_n805), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1213), .B(new_n1216), .C1(G150), .C2(new_n799), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n308), .B(new_n465), .C1(new_n843), .C2(new_n313), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G124), .B2(new_n820), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1060), .B1(G107), .B2(new_n818), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n843), .A2(new_n806), .B1(new_n515), .B2(new_n791), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n391), .A2(new_n804), .B1(new_n808), .B2(new_n517), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n302), .A2(new_n465), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G283), .B2(new_n820), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1224), .A2(new_n1001), .A3(new_n1227), .A4(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT58), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1228), .B(new_n375), .C1(G33), .C2(G41), .ZN(new_n1234));
  AND4_X1   g1034(.A1(new_n1223), .A2(new_n1232), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1211), .B1(new_n1235), .B2(new_n864), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1193), .B2(new_n770), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT119), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1210), .A2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1209), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(G375));
  OR2_X1    g1041(.A1(new_n1148), .A2(new_n1186), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n789), .A2(new_n517), .B1(new_n1069), .B2(new_n805), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n260), .B(new_n1243), .C1(G116), .C2(new_n809), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n795), .A2(G77), .B1(G303), .B2(new_n820), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G294), .A2(new_n849), .B1(new_n816), .B2(G107), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1244), .A2(new_n1062), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n804), .A2(new_n427), .B1(new_n801), .B2(new_n1177), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n302), .B(new_n1248), .C1(G58), .C2(new_n795), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n799), .A2(G50), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1003), .A2(new_n818), .B1(new_n849), .B2(G132), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n788), .A2(G159), .B1(new_n809), .B2(new_n1214), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n864), .B1(new_n1247), .B2(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n767), .B(new_n1254), .C1(new_n298), .C2(new_n841), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n959), .B2(new_n771), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1242), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1161), .A2(new_n1038), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(G381));
  AND2_X1   g1061(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1187), .B1(new_n1262), .B2(new_n1157), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1240), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(G396), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1059), .A2(new_n1265), .A3(new_n1098), .ZN(new_n1266));
  OR4_X1    g1066(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1266), .ZN(new_n1267));
  OR3_X1    g1067(.A1(new_n1264), .A2(G387), .A3(new_n1267), .ZN(G407));
  NOR2_X1   g1068(.A1(new_n695), .A2(G343), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1264), .A2(new_n1270), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT120), .Z(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1266), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1109), .A2(new_n1132), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1107), .B2(new_n1102), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT124), .B1(G387), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(new_n1277), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G387), .A2(KEYINPUT124), .A3(new_n1277), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1275), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(G387), .A2(new_n1277), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(G387), .A2(new_n1277), .B1(new_n1274), .B2(new_n1266), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1283), .A2(new_n1284), .A3(KEYINPUT125), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT125), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1282), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n723), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1259), .A2(KEYINPUT60), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT60), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1142), .A2(new_n1148), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1288), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(G384), .A3(new_n1258), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n866), .B(KEYINPUT100), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1292), .B2(new_n1257), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1209), .A2(new_n1263), .A3(new_n1239), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1239), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1196), .A2(new_n1198), .A3(new_n1038), .A4(new_n1204), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G378), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1270), .B(new_n1299), .C1(new_n1300), .C2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT121), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n723), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(G378), .A3(new_n1301), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1263), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT121), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1311), .A2(new_n1312), .A3(new_n1270), .A4(new_n1299), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT62), .B1(new_n1305), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1270), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1269), .A2(G2897), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT123), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1294), .A2(new_n1297), .A3(new_n1316), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT122), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT122), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1294), .A2(new_n1297), .A3(new_n1322), .A4(new_n1316), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT123), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1325), .B(new_n1317), .C1(new_n1295), .C2(new_n1298), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1319), .A2(new_n1324), .A3(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT61), .B1(new_n1315), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1304), .A2(KEYINPUT62), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1287), .B1(new_n1314), .B2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  OAI21_X1  g1132(.A(KEYINPUT126), .B1(new_n1304), .B2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1269), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT126), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1334), .A2(new_n1335), .A3(KEYINPUT63), .A4(new_n1299), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1333), .A2(new_n1336), .ZN(new_n1337));
  AOI211_X1 g1137(.A(KEYINPUT61), .B(new_n1287), .C1(new_n1315), .C2(new_n1327), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1305), .A2(new_n1313), .A3(new_n1332), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1337), .A2(new_n1338), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1331), .A2(new_n1340), .ZN(G405));
  NAND2_X1  g1141(.A1(G375), .A2(G378), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1264), .ZN(new_n1343));
  OR2_X1    g1143(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1343), .B1(new_n1282), .B2(new_n1344), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1299), .A2(KEYINPUT127), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1342), .A2(new_n1287), .A3(new_n1264), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1345), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1346), .B1(new_n1345), .B2(new_n1347), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(G402));
endmodule


