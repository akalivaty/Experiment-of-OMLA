

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754;

  NAND2_X1 U375 ( .A1(n359), .A2(n395), .ZN(n530) );
  NAND2_X2 U376 ( .A1(n376), .A2(n589), .ZN(n379) );
  XNOR2_X2 U377 ( .A(n409), .B(n444), .ZN(n376) );
  XNOR2_X2 U378 ( .A(n530), .B(n374), .ZN(n411) );
  NAND2_X1 U379 ( .A1(n572), .A2(n696), .ZN(n592) );
  INV_X1 U380 ( .A(G953), .ZN(n748) );
  AND2_X2 U381 ( .A1(n402), .A2(n363), .ZN(n391) );
  AND2_X2 U382 ( .A1(n518), .A2(n517), .ZN(n353) );
  XNOR2_X1 U383 ( .A(n404), .B(G110), .ZN(n467) );
  INV_X1 U384 ( .A(KEYINPUT22), .ZN(n352) );
  BUF_X1 U385 ( .A(n616), .Z(n746) );
  XNOR2_X1 U386 ( .A(n390), .B(KEYINPUT45), .ZN(n615) );
  INV_X1 U387 ( .A(G119), .ZN(n404) );
  XNOR2_X1 U388 ( .A(KEYINPUT69), .B(G101), .ZN(n457) );
  XNOR2_X2 U389 ( .A(n353), .B(n352), .ZN(n524) );
  XNOR2_X1 U390 ( .A(n390), .B(KEYINPUT45), .ZN(n354) );
  INV_X1 U391 ( .A(n550), .ZN(n355) );
  XNOR2_X1 U392 ( .A(n369), .B(n432), .ZN(n519) );
  NAND2_X4 U393 ( .A1(n382), .A2(n380), .ZN(n656) );
  XNOR2_X1 U394 ( .A(n580), .B(KEYINPUT46), .ZN(n581) );
  OR2_X1 U395 ( .A1(n626), .A2(n393), .ZN(n375) );
  NAND2_X1 U396 ( .A1(G469), .A2(n473), .ZN(n393) );
  XNOR2_X1 U397 ( .A(G134), .B(G131), .ZN(n436) );
  XNOR2_X1 U398 ( .A(G128), .B(KEYINPUT94), .ZN(n422) );
  XNOR2_X1 U399 ( .A(G146), .B(G125), .ZN(n458) );
  XOR2_X1 U400 ( .A(KEYINPUT8), .B(KEYINPUT71), .Z(n428) );
  NOR2_X2 U401 ( .A1(n746), .A2(n416), .ZN(n716) );
  NAND2_X1 U402 ( .A1(n354), .A2(KEYINPUT2), .ZN(n416) );
  AND2_X1 U403 ( .A1(n364), .A2(n372), .ZN(n578) );
  NOR2_X1 U404 ( .A1(n721), .A2(G953), .ZN(n406) );
  NOR2_X1 U405 ( .A1(n585), .A2(KEYINPUT47), .ZN(n586) );
  INV_X1 U406 ( .A(G237), .ZN(n472) );
  XNOR2_X1 U407 ( .A(n572), .B(n389), .ZN(n697) );
  INV_X1 U408 ( .A(KEYINPUT38), .ZN(n389) );
  XNOR2_X1 U409 ( .A(G137), .B(KEYINPUT5), .ZN(n448) );
  XOR2_X1 U410 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n449) );
  XOR2_X1 U411 ( .A(G119), .B(G113), .Z(n447) );
  NOR2_X1 U412 ( .A1(G953), .A2(G237), .ZN(n488) );
  NAND2_X1 U413 ( .A1(G234), .A2(G237), .ZN(n479) );
  XNOR2_X1 U414 ( .A(n388), .B(KEYINPUT110), .ZN(n700) );
  NAND2_X1 U415 ( .A1(n697), .A2(n696), .ZN(n388) );
  NOR2_X1 U416 ( .A1(n587), .A2(n552), .ZN(n553) );
  XNOR2_X1 U417 ( .A(n487), .B(n486), .ZN(n518) );
  NAND2_X1 U418 ( .A1(n485), .A2(n358), .ZN(n487) );
  INV_X1 U419 ( .A(KEYINPUT1), .ZN(n374) );
  XNOR2_X1 U420 ( .A(G122), .B(G107), .ZN(n504) );
  XNOR2_X1 U421 ( .A(n415), .B(G116), .ZN(n466) );
  XNOR2_X1 U422 ( .A(KEYINPUT88), .B(KEYINPUT3), .ZN(n415) );
  AND2_X1 U423 ( .A1(n503), .A2(G221), .ZN(n370) );
  XNOR2_X1 U424 ( .A(G143), .B(G131), .ZN(n492) );
  XOR2_X1 U425 ( .A(G140), .B(G122), .Z(n493) );
  XNOR2_X1 U426 ( .A(G110), .B(G104), .ZN(n439) );
  NAND2_X1 U427 ( .A1(n381), .A2(n397), .ZN(n380) );
  NOR2_X1 U428 ( .A1(n716), .A2(KEYINPUT65), .ZN(n397) );
  BUF_X1 U429 ( .A(n518), .Z(n533) );
  INV_X1 U430 ( .A(KEYINPUT70), .ZN(n385) );
  XOR2_X1 U431 ( .A(G134), .B(G116), .Z(n507) );
  XNOR2_X1 U432 ( .A(n579), .B(KEYINPUT40), .ZN(n752) );
  AND2_X1 U433 ( .A1(n407), .A2(n405), .ZN(n722) );
  AND2_X1 U434 ( .A1(n719), .A2(n406), .ZN(n405) );
  XNOR2_X1 U435 ( .A(n718), .B(KEYINPUT83), .ZN(n407) );
  AND2_X1 U436 ( .A1(n638), .A2(n528), .ZN(n356) );
  XOR2_X1 U437 ( .A(n437), .B(KEYINPUT93), .Z(n357) );
  XOR2_X1 U438 ( .A(n484), .B(KEYINPUT92), .Z(n358) );
  AND2_X1 U439 ( .A1(n375), .A2(n394), .ZN(n359) );
  OR2_X1 U440 ( .A1(G902), .A2(n724), .ZN(n360) );
  XOR2_X1 U441 ( .A(n449), .B(n448), .Z(n361) );
  AND2_X1 U442 ( .A1(G217), .A2(n433), .ZN(n362) );
  AND2_X1 U443 ( .A1(n541), .A2(n662), .ZN(n363) );
  NOR2_X1 U444 ( .A1(n683), .A2(n386), .ZN(n364) );
  BUF_X1 U445 ( .A(n530), .Z(n576) );
  INV_X1 U446 ( .A(n576), .ZN(n373) );
  XOR2_X1 U447 ( .A(KEYINPUT66), .B(KEYINPUT32), .Z(n365) );
  XOR2_X1 U448 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n366) );
  XOR2_X1 U449 ( .A(n614), .B(KEYINPUT68), .Z(n367) );
  XNOR2_X1 U450 ( .A(n742), .B(n442), .ZN(n626) );
  AND2_X1 U451 ( .A1(n367), .A2(KEYINPUT65), .ZN(n368) );
  NAND2_X1 U452 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U453 ( .A1(n657), .A2(n473), .ZN(n369) );
  XNOR2_X1 U454 ( .A(n371), .B(n370), .ZN(n657) );
  XNOR2_X1 U455 ( .A(n426), .B(n740), .ZN(n371) );
  NOR2_X1 U456 ( .A1(n752), .A2(n753), .ZN(n582) );
  NOR2_X1 U457 ( .A1(n583), .A2(n584), .ZN(n421) );
  NAND2_X1 U458 ( .A1(n421), .A2(n599), .ZN(n420) );
  AND2_X1 U459 ( .A1(n577), .A2(n373), .ZN(n372) );
  INV_X1 U460 ( .A(n411), .ZN(n526) );
  AND2_X1 U461 ( .A1(n376), .A2(n558), .ZN(n692) );
  NOR2_X1 U462 ( .A1(n574), .A2(n377), .ZN(n674) );
  INV_X1 U463 ( .A(n485), .ZN(n377) );
  XNOR2_X2 U464 ( .A(n592), .B(KEYINPUT19), .ZN(n485) );
  XNOR2_X1 U465 ( .A(n378), .B(n366), .ZN(n513) );
  NAND2_X1 U466 ( .A1(n704), .A2(n533), .ZN(n378) );
  XNOR2_X2 U467 ( .A(n379), .B(KEYINPUT33), .ZN(n704) );
  NAND2_X1 U468 ( .A1(n384), .A2(n367), .ZN(n381) );
  AND2_X2 U469 ( .A1(n383), .A2(n396), .ZN(n382) );
  NAND2_X1 U470 ( .A1(n384), .A2(n368), .ZN(n383) );
  XNOR2_X2 U471 ( .A(n612), .B(n417), .ZN(n384) );
  INV_X1 U472 ( .A(n697), .ZN(n386) );
  INV_X1 U473 ( .A(n387), .ZN(n683) );
  NAND2_X1 U474 ( .A1(n411), .A2(n387), .ZN(n409) );
  XNOR2_X2 U475 ( .A(n410), .B(n385), .ZN(n387) );
  AND2_X1 U476 ( .A1(n387), .A2(n531), .ZN(n532) );
  XNOR2_X2 U477 ( .A(n477), .B(n476), .ZN(n572) );
  NAND2_X1 U478 ( .A1(n615), .A2(n542), .ZN(n544) );
  NAND2_X2 U479 ( .A1(n392), .A2(n391), .ZN(n390) );
  AND2_X2 U480 ( .A1(n400), .A2(n399), .ZN(n392) );
  NAND2_X1 U481 ( .A1(n443), .A2(G902), .ZN(n394) );
  NAND2_X1 U482 ( .A1(n626), .A2(n443), .ZN(n395) );
  NAND2_X1 U483 ( .A1(n716), .A2(KEYINPUT65), .ZN(n396) );
  XNOR2_X1 U484 ( .A(n467), .B(n437), .ZN(n425) );
  NAND2_X1 U485 ( .A1(n401), .A2(KEYINPUT44), .ZN(n400) );
  INV_X1 U486 ( .A(n654), .ZN(n401) );
  XNOR2_X2 U487 ( .A(n515), .B(n514), .ZN(n654) );
  NAND2_X1 U488 ( .A1(n639), .A2(n638), .ZN(n398) );
  AND2_X1 U489 ( .A1(n639), .A2(n356), .ZN(n403) );
  NAND2_X1 U490 ( .A1(n398), .A2(KEYINPUT44), .ZN(n399) );
  NAND2_X1 U491 ( .A1(n654), .A2(n403), .ZN(n402) );
  XNOR2_X2 U492 ( .A(G140), .B(G137), .ZN(n437) );
  XNOR2_X2 U493 ( .A(n408), .B(KEYINPUT4), .ZN(n460) );
  XNOR2_X1 U494 ( .A(n408), .B(n504), .ZN(n506) );
  XNOR2_X2 U495 ( .A(G143), .B(G128), .ZN(n408) );
  NAND2_X1 U496 ( .A1(n519), .A2(n685), .ZN(n410) );
  NOR2_X1 U497 ( .A1(n412), .A2(n574), .ZN(n575) );
  NOR2_X1 U498 ( .A1(n412), .A2(n720), .ZN(n721) );
  NOR2_X1 U499 ( .A1(n695), .A2(n412), .ZN(n707) );
  XNOR2_X1 U500 ( .A(n573), .B(KEYINPUT41), .ZN(n412) );
  XNOR2_X1 U501 ( .A(n466), .B(n413), .ZN(n470) );
  XNOR2_X1 U502 ( .A(n495), .B(n414), .ZN(n413) );
  INV_X1 U503 ( .A(KEYINPUT16), .ZN(n414) );
  XNOR2_X2 U504 ( .A(G113), .B(G104), .ZN(n495) );
  INV_X1 U505 ( .A(KEYINPUT81), .ZN(n417) );
  NAND2_X1 U506 ( .A1(n418), .A2(n609), .ZN(n616) );
  XNOR2_X1 U507 ( .A(n420), .B(n419), .ZN(n418) );
  INV_X1 U508 ( .A(KEYINPUT48), .ZN(n419) );
  INV_X1 U509 ( .A(KEYINPUT82), .ZN(n543) );
  INV_X1 U510 ( .A(KEYINPUT64), .ZN(n580) );
  INV_X1 U511 ( .A(KEYINPUT44), .ZN(n528) );
  INV_X1 U512 ( .A(n635), .ZN(n597) );
  XNOR2_X1 U513 ( .A(n559), .B(KEYINPUT30), .ZN(n560) );
  XNOR2_X1 U514 ( .A(n561), .B(n560), .ZN(n564) );
  BUF_X1 U515 ( .A(n656), .Z(n723) );
  INV_X1 U516 ( .A(KEYINPUT63), .ZN(n624) );
  XOR2_X1 U517 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n423) );
  XNOR2_X1 U518 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U519 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U520 ( .A(n458), .B(KEYINPUT10), .ZN(n740) );
  NAND2_X1 U521 ( .A1(G234), .A2(n748), .ZN(n427) );
  XNOR2_X1 U522 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U523 ( .A(KEYINPUT79), .B(n429), .ZN(n503) );
  INV_X1 U524 ( .A(G902), .ZN(n473) );
  XOR2_X1 U525 ( .A(KEYINPUT25), .B(KEYINPUT95), .Z(n431) );
  XNOR2_X1 U526 ( .A(G902), .B(KEYINPUT15), .ZN(n613) );
  NAND2_X1 U527 ( .A1(n613), .A2(G234), .ZN(n430) );
  XNOR2_X1 U528 ( .A(n430), .B(KEYINPUT20), .ZN(n433) );
  XNOR2_X1 U529 ( .A(n431), .B(n362), .ZN(n432) );
  AND2_X1 U530 ( .A1(n433), .A2(G221), .ZN(n435) );
  XNOR2_X1 U531 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n434) );
  XNOR2_X1 U532 ( .A(n435), .B(n434), .ZN(n685) );
  XNOR2_X2 U533 ( .A(n460), .B(n436), .ZN(n453) );
  XNOR2_X2 U534 ( .A(n453), .B(n357), .ZN(n742) );
  XNOR2_X1 U535 ( .A(n457), .B(G146), .ZN(n445) );
  NAND2_X1 U536 ( .A1(n748), .A2(G227), .ZN(n438) );
  XNOR2_X1 U537 ( .A(n438), .B(G107), .ZN(n440) );
  XNOR2_X1 U538 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U539 ( .A(n445), .B(n441), .ZN(n442) );
  INV_X1 U540 ( .A(G469), .ZN(n443) );
  INV_X1 U541 ( .A(KEYINPUT74), .ZN(n444) );
  XNOR2_X1 U542 ( .A(n445), .B(n466), .ZN(n452) );
  NAND2_X1 U543 ( .A1(n488), .A2(G210), .ZN(n446) );
  XNOR2_X1 U544 ( .A(n447), .B(n446), .ZN(n450) );
  XNOR2_X1 U545 ( .A(n450), .B(n361), .ZN(n451) );
  XNOR2_X1 U546 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U547 ( .A(n453), .B(n454), .ZN(n619) );
  NAND2_X1 U548 ( .A1(n619), .A2(n473), .ZN(n455) );
  XNOR2_X2 U549 ( .A(n455), .B(G472), .ZN(n558) );
  XNOR2_X1 U550 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n456) );
  XNOR2_X1 U551 ( .A(n558), .B(n456), .ZN(n589) );
  XNOR2_X1 U552 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U553 ( .A(n460), .B(n459), .ZN(n465) );
  XOR2_X1 U554 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n463) );
  NAND2_X1 U555 ( .A1(G224), .A2(n748), .ZN(n461) );
  XNOR2_X1 U556 ( .A(n461), .B(KEYINPUT89), .ZN(n462) );
  XNOR2_X1 U557 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U558 ( .A(n465), .B(n464), .ZN(n471) );
  INV_X1 U559 ( .A(n467), .ZN(n468) );
  XNOR2_X1 U560 ( .A(n468), .B(n504), .ZN(n469) );
  XNOR2_X1 U561 ( .A(n470), .B(n469), .ZN(n728) );
  XNOR2_X1 U562 ( .A(n471), .B(n728), .ZN(n646) );
  INV_X1 U563 ( .A(n613), .ZN(n542) );
  OR2_X2 U564 ( .A1(n646), .A2(n542), .ZN(n477) );
  NAND2_X1 U565 ( .A1(n473), .A2(n472), .ZN(n478) );
  NAND2_X1 U566 ( .A1(n478), .A2(G210), .ZN(n475) );
  INV_X1 U567 ( .A(KEYINPUT76), .ZN(n474) );
  XNOR2_X1 U568 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U569 ( .A1(n478), .A2(G214), .ZN(n696) );
  XNOR2_X1 U570 ( .A(n479), .B(KEYINPUT14), .ZN(n481) );
  NAND2_X1 U571 ( .A1(G952), .A2(n481), .ZN(n710) );
  NOR2_X1 U572 ( .A1(G953), .A2(n710), .ZN(n548) );
  NOR2_X1 U573 ( .A1(G898), .A2(n748), .ZN(n480) );
  XOR2_X1 U574 ( .A(KEYINPUT90), .B(n480), .Z(n729) );
  NAND2_X1 U575 ( .A1(G902), .A2(n481), .ZN(n545) );
  NOR2_X1 U576 ( .A1(n729), .A2(n545), .ZN(n482) );
  XOR2_X1 U577 ( .A(KEYINPUT91), .B(n482), .Z(n483) );
  NOR2_X1 U578 ( .A1(n548), .A2(n483), .ZN(n484) );
  INV_X1 U579 ( .A(KEYINPUT0), .ZN(n486) );
  XNOR2_X1 U580 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n500) );
  XOR2_X1 U581 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n490) );
  NAND2_X1 U582 ( .A1(G214), .A2(n488), .ZN(n489) );
  XNOR2_X1 U583 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U584 ( .A(n491), .B(KEYINPUT12), .Z(n498) );
  XNOR2_X1 U585 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U586 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U587 ( .A(n740), .B(n496), .ZN(n497) );
  XNOR2_X1 U588 ( .A(n498), .B(n497), .ZN(n641) );
  NOR2_X1 U589 ( .A1(G902), .A2(n641), .ZN(n499) );
  XNOR2_X1 U590 ( .A(n500), .B(n499), .ZN(n502) );
  INV_X1 U591 ( .A(G475), .ZN(n501) );
  XNOR2_X1 U592 ( .A(n502), .B(n501), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n503), .A2(G217), .ZN(n510) );
  XOR2_X1 U594 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n505) );
  XNOR2_X1 U595 ( .A(n506), .B(n505), .ZN(n508) );
  XNOR2_X1 U596 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U597 ( .A(n510), .B(n509), .ZN(n724) );
  XNOR2_X1 U598 ( .A(G478), .B(n360), .ZN(n535) );
  NAND2_X1 U599 ( .A1(n537), .A2(n535), .ZN(n512) );
  INV_X1 U600 ( .A(KEYINPUT104), .ZN(n511) );
  XNOR2_X1 U601 ( .A(n512), .B(n511), .ZN(n568) );
  NAND2_X1 U602 ( .A1(n513), .A2(n568), .ZN(n515) );
  INV_X1 U603 ( .A(KEYINPUT35), .ZN(n514) );
  OR2_X1 U604 ( .A1(n537), .A2(n535), .ZN(n699) );
  INV_X1 U605 ( .A(n685), .ZN(n516) );
  NOR2_X1 U606 ( .A1(n699), .A2(n516), .ZN(n517) );
  XNOR2_X1 U607 ( .A(n589), .B(KEYINPUT75), .ZN(n521) );
  INV_X1 U608 ( .A(n526), .ZN(n595) );
  INV_X1 U609 ( .A(n519), .ZN(n550) );
  AND2_X1 U610 ( .A1(n595), .A2(n550), .ZN(n520) );
  NAND2_X1 U611 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X2 U612 ( .A1(n524), .A2(n522), .ZN(n523) );
  XNOR2_X2 U613 ( .A(n523), .B(n365), .ZN(n639) );
  NOR2_X1 U614 ( .A1(n355), .A2(n558), .ZN(n525) );
  NAND2_X1 U615 ( .A1(n526), .A2(n525), .ZN(n527) );
  OR2_X1 U616 ( .A1(n524), .A2(n527), .ZN(n638) );
  NAND2_X1 U617 ( .A1(n692), .A2(n533), .ZN(n529) );
  XNOR2_X1 U618 ( .A(n529), .B(KEYINPUT31), .ZN(n680) );
  NOR2_X1 U619 ( .A1(n576), .A2(n558), .ZN(n531) );
  NAND2_X1 U620 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U621 ( .A(n534), .B(KEYINPUT99), .ZN(n667) );
  OR2_X1 U622 ( .A1(n680), .A2(n667), .ZN(n538) );
  INV_X1 U623 ( .A(n535), .ZN(n536) );
  NOR2_X1 U624 ( .A1(n537), .A2(n536), .ZN(n679) );
  XOR2_X1 U625 ( .A(KEYINPUT102), .B(n679), .Z(n608) );
  NAND2_X1 U626 ( .A1(n537), .A2(n536), .ZN(n588) );
  AND2_X1 U627 ( .A1(n608), .A2(n588), .ZN(n701) );
  INV_X1 U628 ( .A(n701), .ZN(n557) );
  NAND2_X1 U629 ( .A1(n538), .A2(n557), .ZN(n541) );
  NOR2_X1 U630 ( .A1(n589), .A2(n550), .ZN(n539) );
  NAND2_X1 U631 ( .A1(n539), .A2(n526), .ZN(n540) );
  OR2_X1 U632 ( .A1(n524), .A2(n540), .ZN(n662) );
  XNOR2_X1 U633 ( .A(n544), .B(n543), .ZN(n611) );
  INV_X1 U634 ( .A(KEYINPUT28), .ZN(n554) );
  OR2_X1 U635 ( .A1(n748), .A2(n545), .ZN(n546) );
  NOR2_X1 U636 ( .A1(G900), .A2(n546), .ZN(n547) );
  NOR2_X1 U637 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U638 ( .A(KEYINPUT77), .B(n549), .ZN(n562) );
  AND2_X1 U639 ( .A1(n562), .A2(n550), .ZN(n551) );
  NAND2_X1 U640 ( .A1(n685), .A2(n551), .ZN(n587) );
  INV_X1 U641 ( .A(n558), .ZN(n552) );
  XNOR2_X1 U642 ( .A(n554), .B(n553), .ZN(n555) );
  NOR2_X1 U643 ( .A1(n555), .A2(n576), .ZN(n556) );
  XNOR2_X1 U644 ( .A(n556), .B(KEYINPUT109), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n674), .A2(n557), .ZN(n585) );
  NAND2_X1 U646 ( .A1(n585), .A2(KEYINPUT47), .ZN(n570) );
  NAND2_X1 U647 ( .A1(n558), .A2(n696), .ZN(n561) );
  XOR2_X1 U648 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n559) );
  INV_X1 U649 ( .A(n562), .ZN(n563) );
  NOR2_X1 U650 ( .A1(n564), .A2(n563), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n577), .A2(n373), .ZN(n565) );
  NOR2_X1 U652 ( .A1(n565), .A2(n683), .ZN(n566) );
  BUF_X1 U653 ( .A(n572), .Z(n604) );
  NAND2_X1 U654 ( .A1(n566), .A2(n604), .ZN(n567) );
  XOR2_X1 U655 ( .A(KEYINPUT108), .B(n567), .Z(n569) );
  NAND2_X1 U656 ( .A1(n569), .A2(n568), .ZN(n673) );
  NAND2_X1 U657 ( .A1(n570), .A2(n673), .ZN(n571) );
  XNOR2_X1 U658 ( .A(n571), .B(KEYINPUT78), .ZN(n584) );
  NOR2_X1 U659 ( .A1(n700), .A2(n699), .ZN(n573) );
  XNOR2_X1 U660 ( .A(n575), .B(KEYINPUT42), .ZN(n753) );
  XNOR2_X1 U661 ( .A(n578), .B(KEYINPUT39), .ZN(n607) );
  NOR2_X1 U662 ( .A1(n607), .A2(n588), .ZN(n579) );
  XNOR2_X1 U663 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U664 ( .A(KEYINPUT73), .B(n586), .Z(n598) );
  INV_X1 U665 ( .A(n587), .ZN(n591) );
  XNOR2_X1 U666 ( .A(n588), .B(KEYINPUT105), .ZN(n677) );
  AND2_X1 U667 ( .A1(n589), .A2(n677), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n601) );
  NOR2_X1 U669 ( .A1(n601), .A2(n592), .ZN(n594) );
  XNOR2_X1 U670 ( .A(KEYINPUT84), .B(KEYINPUT36), .ZN(n593) );
  XNOR2_X1 U671 ( .A(n594), .B(n593), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n635) );
  NOR2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  INV_X1 U674 ( .A(n696), .ZN(n600) );
  NOR2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n602), .A2(n526), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT43), .ZN(n606) );
  INV_X1 U678 ( .A(n604), .ZN(n605) );
  AND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n636) );
  NOR2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n682) );
  NOR2_X1 U681 ( .A1(n636), .A2(n682), .ZN(n609) );
  INV_X1 U682 ( .A(n616), .ZN(n610) );
  INV_X1 U683 ( .A(KEYINPUT2), .ZN(n713) );
  NOR2_X1 U684 ( .A1(n613), .A2(n713), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n656), .A2(G472), .ZN(n621) );
  XOR2_X1 U686 ( .A(KEYINPUT87), .B(KEYINPUT111), .Z(n617) );
  XNOR2_X1 U687 ( .A(n617), .B(KEYINPUT62), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n621), .B(n620), .ZN(n623) );
  INV_X1 U690 ( .A(G952), .ZN(n622) );
  AND2_X1 U691 ( .A1(n622), .A2(G953), .ZN(n727) );
  NOR2_X2 U692 ( .A1(n623), .A2(n727), .ZN(n625) );
  XNOR2_X1 U693 ( .A(n625), .B(n624), .ZN(G57) );
  NAND2_X1 U694 ( .A1(n656), .A2(G469), .ZN(n630) );
  XOR2_X1 U695 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n627) );
  XNOR2_X1 U696 ( .A(n627), .B(KEYINPUT58), .ZN(n628) );
  XNOR2_X1 U697 ( .A(n626), .B(n628), .ZN(n629) );
  XNOR2_X1 U698 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X2 U699 ( .A1(n631), .A2(n727), .ZN(n633) );
  INV_X1 U700 ( .A(KEYINPUT121), .ZN(n632) );
  XNOR2_X1 U701 ( .A(n633), .B(n632), .ZN(G54) );
  XOR2_X1 U702 ( .A(G125), .B(KEYINPUT37), .Z(n634) );
  XNOR2_X1 U703 ( .A(n635), .B(n634), .ZN(G27) );
  XNOR2_X1 U704 ( .A(G140), .B(KEYINPUT116), .ZN(n637) );
  XOR2_X1 U705 ( .A(n637), .B(n636), .Z(G42) );
  XNOR2_X1 U706 ( .A(n638), .B(G110), .ZN(G12) );
  XNOR2_X1 U707 ( .A(n639), .B(G119), .ZN(G21) );
  NAND2_X1 U708 ( .A1(n656), .A2(G475), .ZN(n643) );
  XNOR2_X1 U709 ( .A(KEYINPUT67), .B(KEYINPUT59), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(n644) );
  NOR2_X2 U712 ( .A1(n644), .A2(n727), .ZN(n645) );
  XNOR2_X1 U713 ( .A(n645), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U714 ( .A1(n656), .A2(G210), .ZN(n651) );
  XNOR2_X1 U715 ( .A(KEYINPUT86), .B(KEYINPUT54), .ZN(n648) );
  XNOR2_X1 U716 ( .A(KEYINPUT55), .B(KEYINPUT85), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n646), .B(n649), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X2 U720 ( .A1(n652), .A2(n727), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n653), .B(KEYINPUT56), .ZN(G51) );
  BUF_X1 U722 ( .A(n654), .Z(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(G122), .ZN(G24) );
  NAND2_X1 U724 ( .A1(n723), .A2(G217), .ZN(n660) );
  BUF_X1 U725 ( .A(n657), .Z(n658) );
  XOR2_X1 U726 ( .A(n658), .B(KEYINPUT122), .Z(n659) );
  XNOR2_X1 U727 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U728 ( .A1(n661), .A2(n727), .ZN(G66) );
  XNOR2_X1 U729 ( .A(G101), .B(n662), .ZN(G3) );
  NAND2_X1 U730 ( .A1(n667), .A2(n677), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n663), .B(G104), .ZN(G6) );
  XOR2_X1 U732 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n665) );
  XNOR2_X1 U733 ( .A(G107), .B(KEYINPUT112), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n665), .B(n664), .ZN(n666) );
  XOR2_X1 U735 ( .A(KEYINPUT26), .B(n666), .Z(n669) );
  NAND2_X1 U736 ( .A1(n667), .A2(n679), .ZN(n668) );
  XNOR2_X1 U737 ( .A(n669), .B(n668), .ZN(G9) );
  XOR2_X1 U738 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n671) );
  NAND2_X1 U739 ( .A1(n674), .A2(n679), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U741 ( .A(G128), .B(n672), .ZN(G30) );
  XNOR2_X1 U742 ( .A(G143), .B(n673), .ZN(G45) );
  XOR2_X1 U743 ( .A(G146), .B(KEYINPUT115), .Z(n676) );
  NAND2_X1 U744 ( .A1(n674), .A2(n677), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n676), .B(n675), .ZN(G48) );
  NAND2_X1 U746 ( .A1(n680), .A2(n677), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n678), .B(G113), .ZN(G15) );
  NAND2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n681), .B(G116), .ZN(G18) );
  XOR2_X1 U750 ( .A(G134), .B(n682), .Z(G36) );
  NAND2_X1 U751 ( .A1(n683), .A2(n526), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n684), .B(KEYINPUT50), .ZN(n689) );
  NOR2_X1 U753 ( .A1(n685), .A2(n355), .ZN(n686) );
  XOR2_X1 U754 ( .A(KEYINPUT49), .B(n686), .Z(n687) );
  XNOR2_X1 U755 ( .A(KEYINPUT117), .B(n687), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n558), .A2(n690), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(KEYINPUT118), .ZN(n693) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U760 ( .A(KEYINPUT51), .B(n694), .Z(n695) );
  NOR2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n705) );
  INV_X1 U765 ( .A(n704), .ZN(n720) );
  NOR2_X1 U766 ( .A1(n705), .A2(n720), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U768 ( .A(n708), .B(KEYINPUT52), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U770 ( .A(KEYINPUT119), .B(n711), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n354), .A2(KEYINPUT2), .ZN(n712) );
  XOR2_X1 U772 ( .A(KEYINPUT80), .B(n712), .Z(n715) );
  NAND2_X1 U773 ( .A1(n746), .A2(n713), .ZN(n714) );
  NAND2_X1 U774 ( .A1(n715), .A2(n714), .ZN(n717) );
  NOR2_X1 U775 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U776 ( .A(KEYINPUT53), .B(n722), .ZN(G75) );
  NAND2_X1 U777 ( .A1(n723), .A2(G478), .ZN(n725) );
  XNOR2_X1 U778 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n727), .A2(n726), .ZN(G63) );
  XNOR2_X1 U780 ( .A(n728), .B(G101), .ZN(n730) );
  NAND2_X1 U781 ( .A1(n730), .A2(n729), .ZN(n739) );
  INV_X1 U782 ( .A(n354), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n731), .A2(G953), .ZN(n737) );
  XOR2_X1 U784 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n733) );
  NAND2_X1 U785 ( .A1(G224), .A2(G953), .ZN(n732) );
  XNOR2_X1 U786 ( .A(n733), .B(n732), .ZN(n734) );
  NAND2_X1 U787 ( .A1(G898), .A2(n734), .ZN(n735) );
  XOR2_X1 U788 ( .A(KEYINPUT124), .B(n735), .Z(n736) );
  NOR2_X1 U789 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U790 ( .A(n739), .B(n738), .ZN(G69) );
  XNOR2_X1 U791 ( .A(n740), .B(KEYINPUT125), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(n747) );
  XNOR2_X1 U793 ( .A(n747), .B(KEYINPUT126), .ZN(n743) );
  XNOR2_X1 U794 ( .A(G227), .B(n743), .ZN(n744) );
  NAND2_X1 U795 ( .A1(G900), .A2(n744), .ZN(n745) );
  NAND2_X1 U796 ( .A1(n745), .A2(G953), .ZN(n751) );
  XNOR2_X1 U797 ( .A(n747), .B(n746), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U799 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U800 ( .A(n752), .B(G131), .Z(G33) );
  XNOR2_X1 U801 ( .A(G137), .B(KEYINPUT127), .ZN(n754) );
  XNOR2_X1 U802 ( .A(n754), .B(n753), .ZN(G39) );
endmodule

