//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT65), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n207), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n203), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n226), .A2(G50), .A3(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n210), .B(new_n221), .C1(new_n224), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G97), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT73), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G223), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n249), .B1(new_n202), .B2(new_n247), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT67), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n260), .B(new_n257), .C1(G41), .C2(G45), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n259), .A2(G274), .A3(new_n254), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n254), .A2(new_n258), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT68), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n254), .A2(new_n265), .A3(new_n258), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G226), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n256), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n201), .A2(new_n203), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n273), .A2(G20), .B1(G150), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT69), .A2(G58), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT69), .A2(G58), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT8), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(KEYINPUT8), .B2(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n223), .A2(G33), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n222), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G50), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n283), .A2(new_n222), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(G1), .B2(new_n223), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n290), .B2(G50), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n269), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n272), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n292), .A2(new_n297), .B1(new_n269), .B2(G200), .ZN(new_n298));
  INV_X1    g0098(.A(new_n292), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n270), .A2(G190), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n298), .A2(new_n304), .A3(new_n300), .A4(new_n301), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n296), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G20), .A2(G77), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT15), .B(G87), .ZN(new_n309));
  INV_X1    g0109(.A(new_n274), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT8), .B(G58), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n308), .B1(new_n309), .B2(new_n281), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n312), .A2(new_n284), .ZN(new_n313));
  INV_X1    g0113(.A(new_n286), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n202), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n289), .B2(new_n202), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT71), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n316), .B1(new_n284), .B2(new_n312), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n267), .A2(G244), .ZN(new_n322));
  INV_X1    g0122(.A(G107), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n250), .A2(new_n215), .B1(new_n323), .B2(new_n247), .ZN(new_n324));
  INV_X1    g0124(.A(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n329), .A2(new_n213), .A3(G1698), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n255), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n322), .A2(new_n331), .A3(new_n262), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n293), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n321), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT72), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n332), .A2(G179), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT72), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n321), .A2(new_n337), .A3(new_n333), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n321), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n332), .A2(KEYINPUT70), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT70), .B1(new_n332), .B2(new_n341), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n332), .A2(G200), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n340), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n246), .B1(new_n307), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n280), .A2(new_n314), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n289), .B2(new_n280), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT7), .B1(new_n329), .B2(new_n223), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  AOI211_X1 g0152(.A(new_n352), .B(G20), .C1(new_n326), .C2(new_n328), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G159), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n310), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT69), .B(G58), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n225), .B1(new_n357), .B2(new_n214), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n358), .B2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n288), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n354), .A2(KEYINPUT16), .A3(new_n359), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n350), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n254), .A2(G232), .A3(new_n258), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n262), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(G179), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n326), .A2(new_n328), .A3(G226), .A4(G1698), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n326), .A2(new_n328), .A3(G223), .A4(new_n248), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G87), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT79), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n371), .A2(new_n372), .A3(new_n255), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n372), .B1(new_n371), .B2(new_n255), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n367), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n371), .A2(new_n255), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n293), .B1(new_n377), .B2(new_n366), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n348), .B1(new_n364), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n203), .B1(new_n278), .B2(G68), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n381), .A2(new_n223), .B1(new_n355), .B2(new_n310), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n352), .B1(new_n247), .B2(G20), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n327), .A2(G33), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n385));
  OAI211_X1 g0185(.A(KEYINPUT7), .B(new_n223), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n214), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n361), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(new_n363), .A3(new_n284), .ZN(new_n389));
  INV_X1    g0189(.A(new_n350), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n375), .A2(new_n378), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT18), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n380), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n339), .A4(new_n345), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n396), .A2(KEYINPUT81), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n262), .A2(new_n341), .A3(new_n365), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n376), .A2(KEYINPUT79), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n371), .A2(new_n372), .A3(new_n255), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n262), .A2(new_n365), .ZN(new_n403));
  AOI21_X1  g0203(.A(G200), .B1(new_n403), .B2(new_n376), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT80), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n399), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n373), .B2(new_n374), .ZN(new_n407));
  INV_X1    g0207(.A(G200), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n377), .B2(new_n366), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT80), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n391), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n396), .A2(KEYINPUT81), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n398), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n402), .A2(KEYINPUT80), .A3(new_n404), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n410), .B1(new_n407), .B2(new_n409), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n364), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n397), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n347), .A2(new_n394), .A3(new_n395), .A4(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n247), .A2(G232), .A3(G1698), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n247), .A2(G226), .A3(new_n248), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G97), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n255), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n264), .A2(G238), .A3(new_n266), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n262), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT74), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(KEYINPUT74), .A3(new_n262), .ZN(new_n432));
  AOI211_X1 g0232(.A(KEYINPUT13), .B(new_n427), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n432), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(new_n426), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G190), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n214), .A2(G20), .ZN(new_n439));
  INV_X1    g0239(.A(G50), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n439), .B1(new_n281), .B2(new_n202), .C1(new_n310), .C2(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n441), .A2(new_n284), .ZN(new_n442));
  XOR2_X1   g0242(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n443));
  OR2_X1    g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT12), .B1(new_n314), .B2(new_n214), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n314), .A2(KEYINPUT12), .A3(new_n214), .ZN(new_n447));
  AOI211_X1 g0247(.A(new_n446), .B(new_n447), .C1(new_n290), .C2(G68), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT76), .ZN(new_n450));
  OAI21_X1  g0250(.A(G200), .B1(new_n433), .B2(new_n436), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n438), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT77), .B(KEYINPUT14), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n437), .B2(new_n293), .ZN(new_n455));
  INV_X1    g0255(.A(new_n432), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT74), .B1(new_n428), .B2(new_n262), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n426), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT13), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n435), .A2(new_n434), .A3(new_n426), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(G179), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT78), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT78), .A4(G179), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT14), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(KEYINPUT77), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(G169), .B(new_n467), .C1(new_n433), .C2(new_n436), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n455), .A2(new_n463), .A3(new_n464), .A4(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n450), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n452), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  INV_X1    g0274(.A(G41), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G41), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n474), .A2(new_n476), .A3(new_n478), .A4(G274), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n257), .B(G45), .C1(new_n475), .C2(KEYINPUT5), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n477), .A2(G41), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n254), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G257), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n326), .A2(new_n328), .A3(G244), .A4(new_n248), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G283), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n255), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT83), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT83), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n494), .A3(new_n255), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n484), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT84), .B1(new_n496), .B2(new_n408), .ZN(new_n497));
  INV_X1    g0297(.A(new_n484), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n491), .A2(new_n494), .A3(new_n255), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n494), .B1(new_n491), .B2(new_n255), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT84), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(G200), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n243), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n323), .A2(KEYINPUT6), .A3(G97), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(G20), .B1(G77), .B2(new_n274), .ZN(new_n508));
  OAI21_X1  g0308(.A(G107), .B1(new_n351), .B2(new_n353), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n284), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n257), .A2(G33), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n286), .A2(new_n512), .A3(new_n222), .A4(new_n283), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G97), .ZN(new_n514));
  INV_X1    g0314(.A(G97), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n286), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT82), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n492), .A2(new_n498), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(new_n341), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n497), .A2(new_n503), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n293), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n519), .B(new_n524), .C1(new_n501), .C2(G179), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n247), .A2(new_n223), .A3(G68), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n223), .B1(new_n424), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G87), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n515), .A3(new_n323), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n527), .B1(new_n281), .B2(new_n515), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n526), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n284), .B1(new_n314), .B2(new_n309), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n513), .A2(new_n529), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n247), .A2(G238), .A3(new_n248), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n247), .A2(G244), .A3(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G116), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n255), .ZN(new_n541));
  INV_X1    g0341(.A(G250), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n257), .B2(G45), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT85), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n254), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n254), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(KEYINPUT85), .B1(G274), .B2(new_n474), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n541), .A2(G190), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n545), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n255), .B2(new_n540), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n536), .B(new_n548), .C1(new_n408), .C2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n293), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n534), .B1(new_n309), .B2(new_n513), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n541), .A2(new_n271), .A3(new_n545), .A4(new_n547), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n326), .A2(new_n328), .A3(G250), .A4(new_n248), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT88), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n247), .A2(KEYINPUT88), .A3(G250), .A4(new_n248), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G294), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n326), .A2(new_n328), .A3(G257), .A4(G1698), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT89), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n563), .A2(new_n562), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(KEYINPUT89), .A3(new_n561), .A4(new_n560), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n255), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n482), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G264), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n479), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G200), .ZN(new_n573));
  OR3_X1    g0373(.A1(new_n286), .A2(KEYINPUT25), .A3(G107), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT25), .B1(new_n286), .B2(G107), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(new_n575), .C1(new_n323), .C2(new_n513), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n576), .B(KEYINPUT87), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT23), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n223), .B2(G107), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n323), .A2(KEYINPUT23), .A3(G20), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(G20), .B2(new_n539), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n326), .A2(new_n328), .A3(new_n223), .A4(G87), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT22), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT22), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n247), .A2(new_n585), .A3(new_n223), .A4(G87), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n582), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n284), .B1(new_n587), .B2(KEYINPUT24), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(KEYINPUT24), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n577), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n569), .A2(G190), .A3(new_n479), .A4(new_n571), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n573), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n523), .A2(new_n525), .A3(new_n557), .A4(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G116), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n314), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n513), .B2(new_n595), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(G20), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n284), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT86), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n284), .A2(KEYINPUT86), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n489), .B(new_n223), .C1(G33), .C2(new_n515), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT20), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n284), .A2(KEYINPUT86), .A3(new_n599), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT86), .B1(new_n284), .B2(new_n599), .ZN(new_n608));
  OAI211_X1 g0408(.A(KEYINPUT20), .B(new_n605), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n598), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(G303), .B1(new_n384), .B2(new_n385), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n326), .A2(new_n328), .A3(G257), .A4(new_n248), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n326), .A2(new_n328), .A3(G264), .A4(G1698), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n255), .ZN(new_n616));
  OAI211_X1 g0416(.A(G270), .B(new_n254), .C1(new_n480), .C2(new_n481), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n617), .A2(new_n479), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n293), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n611), .A2(KEYINPUT21), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n597), .B1(new_n624), .B2(new_n609), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n616), .A2(new_n618), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G169), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n621), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n626), .A2(new_n271), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n611), .A2(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n620), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT87), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n576), .B(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n590), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(new_n588), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n569), .A2(new_n271), .A3(new_n479), .A4(new_n571), .ZN(new_n636));
  INV_X1    g0436(.A(new_n479), .ZN(new_n637));
  INV_X1    g0437(.A(new_n571), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n254), .B1(new_n564), .B2(new_n565), .ZN(new_n639));
  AOI211_X1 g0439(.A(new_n637), .B(new_n638), .C1(new_n639), .C2(new_n568), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n635), .B(new_n636), .C1(new_n640), .C2(G169), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n626), .A2(G200), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n625), .B(new_n642), .C1(new_n341), .C2(new_n626), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n631), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NOR4_X1   g0444(.A1(new_n421), .A2(new_n472), .A3(new_n594), .A4(new_n644), .ZN(G372));
  NOR2_X1   g0445(.A1(new_n421), .A2(new_n472), .ZN(new_n646));
  INV_X1    g0446(.A(new_n556), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT82), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n517), .B(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n288), .B1(new_n508), .B2(new_n509), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n484), .B1(new_n491), .B2(new_n255), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n649), .A2(new_n650), .B1(G169), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n271), .B2(new_n496), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n557), .A2(KEYINPUT26), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n551), .A2(new_n556), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n656), .B2(new_n525), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n647), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n620), .A2(new_n628), .A3(new_n630), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n659), .B(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(new_n641), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n658), .B1(new_n662), .B2(new_n594), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n646), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n293), .B1(new_n459), .B2(new_n460), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n468), .B1(new_n665), .B2(new_n453), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n463), .A2(new_n464), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n470), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(new_n339), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n438), .A2(new_n450), .A3(new_n451), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n420), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n394), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n303), .A2(new_n305), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n296), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n664), .A2(new_n674), .ZN(G369));
  AND2_X1   g0475(.A1(new_n223), .A2(G13), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n257), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n625), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n661), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n685), .B(new_n643), .C1(new_n631), .C2(new_n684), .ZN(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n641), .A2(new_n682), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n593), .B1(new_n591), .B2(new_n683), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n641), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n659), .A2(new_n683), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT91), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n691), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n641), .A2(new_n682), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n692), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n208), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n530), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n228), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n631), .A2(new_n641), .A3(new_n643), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n511), .B(new_n518), .C1(new_n341), .C2(new_n520), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n501), .A2(G200), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(KEYINPUT84), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n653), .B1(new_n710), .B2(new_n503), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n635), .B1(new_n640), .B2(G190), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n656), .B1(new_n712), .B2(new_n573), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n707), .A2(new_n711), .A3(new_n713), .A4(new_n683), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT31), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n552), .A2(new_n271), .A3(new_n626), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(new_n572), .A3(new_n501), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n569), .A2(new_n550), .A3(new_n571), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT92), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT92), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n569), .A2(new_n550), .A3(new_n720), .A4(new_n571), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n520), .A2(new_n271), .A3(new_n626), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n719), .A2(KEYINPUT30), .A3(new_n721), .A4(new_n722), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n683), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(KEYINPUT31), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n715), .A2(new_n728), .B1(new_n729), .B2(KEYINPUT93), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n727), .A2(KEYINPUT31), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT93), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n687), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT29), .B1(new_n663), .B2(new_n683), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n631), .A2(new_n641), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n658), .B1(new_n594), .B2(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n737), .A2(KEYINPUT29), .A3(new_n683), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT94), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n738), .A2(KEYINPUT94), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n734), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n706), .B1(new_n741), .B2(G1), .ZN(G364));
  AOI21_X1  g0542(.A(new_n257), .B1(new_n676), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n701), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n700), .A2(new_n329), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n747), .A2(G355), .B1(new_n595), .B2(new_n700), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n241), .A2(G45), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n700), .A2(new_n247), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n228), .B2(G45), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n222), .B1(G20), .B2(new_n293), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n746), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n341), .A2(G20), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n271), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n329), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n408), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n760), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G329), .A2(new_n767), .B1(new_n770), .B2(G283), .ZN(new_n771));
  INV_X1    g0571(.A(G303), .ZN(new_n772));
  NAND2_X1  g0572(.A1(G20), .A2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G326), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n271), .A2(new_n408), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n774), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n771), .B1(new_n772), .B2(new_n775), .C1(new_n776), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n223), .B1(new_n765), .B2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n764), .B(new_n779), .C1(G294), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n760), .A2(new_n777), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT33), .B(G317), .Z(new_n784));
  NAND2_X1  g0584(.A1(new_n761), .A2(new_n774), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT96), .Z(new_n788));
  AND2_X1   g0588(.A1(new_n780), .A2(KEYINPUT95), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n780), .A2(KEYINPUT95), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G97), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n767), .A2(G159), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  INV_X1    g0595(.A(new_n778), .ZN(new_n796));
  INV_X1    g0596(.A(new_n775), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G50), .A2(new_n796), .B1(new_n797), .B2(G87), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n798), .B(new_n247), .C1(new_n202), .C2(new_n762), .ZN(new_n799));
  INV_X1    g0599(.A(new_n783), .ZN(new_n800));
  INV_X1    g0600(.A(new_n785), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n800), .A2(G68), .B1(new_n801), .B2(new_n278), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n323), .B2(new_n769), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n795), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n782), .A2(new_n788), .B1(new_n793), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n756), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n758), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n686), .B2(new_n755), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n688), .A2(new_n745), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n686), .A2(new_n687), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NAND2_X1  g0612(.A1(new_n663), .A2(new_n683), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n321), .A2(new_n682), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n338), .A2(new_n336), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n337), .B1(new_n321), .B2(new_n333), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n345), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT97), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n339), .A2(new_n814), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n339), .A2(KEYINPUT97), .A3(new_n345), .A4(new_n814), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n813), .B(new_n823), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n594), .A2(new_n644), .A3(new_n682), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT31), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n728), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n729), .A2(KEYINPUT93), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n733), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G330), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n745), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n830), .B2(new_n824), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n756), .A2(new_n753), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n745), .B1(new_n834), .B2(G77), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n769), .A2(new_n529), .B1(new_n766), .B2(new_n763), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n778), .A2(new_n772), .B1(new_n775), .B2(new_n323), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n762), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n247), .B1(new_n839), .B2(G116), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n800), .A2(G283), .B1(new_n801), .B2(G294), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n793), .A2(new_n838), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n762), .A2(new_n355), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  INV_X1    g0644(.A(G143), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n783), .A2(new_n844), .B1(new_n785), .B2(new_n845), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n843), .B(new_n846), .C1(G137), .C2(new_n796), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT34), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n247), .B1(new_n775), .B2(new_n440), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n769), .A2(new_n214), .B1(new_n766), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(new_n278), .C2(new_n781), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n847), .A2(KEYINPUT34), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n842), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n835), .B1(new_n855), .B2(new_n756), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n822), .B2(new_n754), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n832), .A2(new_n857), .ZN(G384));
  OAI211_X1 g0658(.A(G116), .B(new_n224), .C1(new_n507), .C2(KEYINPUT35), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(KEYINPUT35), .B2(new_n507), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT36), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n229), .B(G77), .C1(new_n214), .C2(new_n357), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n201), .A2(G68), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n257), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n470), .A2(new_n682), .ZN(new_n866));
  INV_X1    g0666(.A(new_n666), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n463), .A2(new_n464), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n450), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n471), .A2(new_n866), .B1(new_n869), .B2(new_n682), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n663), .A2(new_n683), .A3(new_n822), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n339), .A2(new_n682), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n870), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  INV_X1    g0675(.A(new_n680), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n391), .B1(new_n392), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n875), .B1(new_n418), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n418), .A2(new_n877), .A3(new_n875), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT99), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n880), .A2(KEYINPUT98), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n880), .B2(KEYINPUT98), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n379), .A2(new_n680), .B1(new_n389), .B2(new_n390), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n412), .A2(KEYINPUT37), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT98), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT99), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n880), .A2(KEYINPUT98), .A3(new_n881), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n878), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n397), .B1(new_n418), .B2(new_n413), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n412), .A2(new_n398), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n394), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n391), .A2(new_n876), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n884), .A2(new_n890), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n884), .A2(new_n890), .A3(KEYINPUT38), .A4(new_n896), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n874), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n394), .B2(new_n876), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(KEYINPUT39), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n893), .A2(new_n895), .B1(new_n879), .B2(new_n880), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT101), .B1(new_n905), .B2(KEYINPUT38), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT101), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n894), .B1(new_n420), .B2(new_n394), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n886), .A2(new_n878), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n907), .B(new_n898), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n900), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n904), .B1(KEYINPUT39), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n469), .A2(new_n470), .A3(new_n683), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT100), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n903), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n739), .A2(new_n646), .A3(new_n740), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n674), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n727), .B1(new_n714), .B2(KEYINPUT31), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n822), .B1(new_n920), .B2(new_n731), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n870), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n901), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n900), .A2(new_n906), .A3(new_n910), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n827), .A2(new_n729), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n668), .A2(new_n670), .A3(new_n866), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n469), .A2(new_n470), .A3(new_n682), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n927), .A2(KEYINPUT40), .A3(new_n822), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT102), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT102), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n922), .A2(new_n911), .A3(new_n933), .A4(KEYINPUT40), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n925), .A2(G330), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n646), .A2(G330), .A3(new_n927), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n922), .A2(new_n911), .A3(KEYINPUT40), .ZN(new_n938));
  AOI22_X1  g0738(.A1(KEYINPUT102), .A2(new_n938), .B1(new_n923), .B2(new_n924), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n939), .A2(new_n646), .A3(new_n927), .A4(new_n934), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n919), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n257), .B2(new_n676), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n919), .B1(new_n937), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n865), .B1(new_n942), .B2(new_n943), .ZN(G367));
  OR2_X1    g0744(.A1(new_n536), .A2(new_n683), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n556), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n557), .A2(new_n945), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n946), .B1(new_n947), .B2(KEYINPUT103), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(KEYINPUT103), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n519), .A2(new_n682), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n711), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n525), .B2(new_n683), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n691), .A3(new_n694), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n525), .B1(new_n952), .B2(new_n641), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n683), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n950), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT104), .Z(new_n961));
  INV_X1    g0761(.A(new_n953), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n692), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n964), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n701), .B(KEYINPUT41), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT107), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n688), .A2(new_n971), .B1(new_n691), .B2(new_n694), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n695), .B(KEYINPUT106), .Z(new_n973));
  NOR3_X1   g0773(.A1(new_n686), .A2(KEYINPUT107), .A3(new_n687), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n972), .B2(new_n973), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n741), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT108), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(KEYINPUT108), .A3(new_n741), .ZN(new_n981));
  INV_X1    g0781(.A(new_n692), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n698), .A2(new_n953), .ZN(new_n983));
  XOR2_X1   g0783(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n697), .A2(KEYINPUT44), .A3(new_n962), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT44), .B1(new_n697), .B2(new_n962), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n982), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n985), .A2(new_n991), .A3(new_n692), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n980), .A2(new_n981), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n970), .B1(new_n993), .B2(new_n741), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n967), .B(new_n968), .C1(new_n744), .C2(new_n994), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n237), .A2(new_n700), .A3(new_n247), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n757), .B1(new_n208), .B2(new_n309), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n745), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(G283), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n515), .A2(new_n769), .B1(new_n762), .B2(new_n999), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n247), .B(new_n1000), .C1(G303), .C2(new_n801), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n797), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT46), .B1(new_n797), .B2(G116), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G107), .B2(new_n781), .ZN(new_n1004));
  INV_X1    g0804(.A(G317), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n766), .A2(new_n1005), .B1(new_n778), .B2(new_n763), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G294), .B2(new_n800), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n791), .A2(new_n214), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n357), .A2(new_n775), .B1(new_n785), .B2(new_n844), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n329), .B(new_n1010), .C1(G77), .C2(new_n770), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n201), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n839), .A2(new_n1012), .B1(new_n796), .B2(G143), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G159), .A2(new_n800), .B1(new_n767), .B2(G137), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1008), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT109), .Z(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(KEYINPUT47), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n806), .B1(new_n1017), .B2(KEYINPUT47), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n998), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n755), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n949), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n995), .A2(new_n1022), .ZN(G387));
  AOI21_X1  g0823(.A(new_n702), .B1(new_n977), .B2(new_n741), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n741), .B2(new_n977), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n977), .A2(new_n744), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n329), .B1(new_n766), .B2(new_n776), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n839), .A2(G303), .B1(new_n801), .B2(G317), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT110), .B(G322), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1028), .B1(new_n763), .B2(new_n783), .C1(new_n778), .C2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  INV_X1    g0831(.A(G294), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1031), .B1(new_n999), .B2(new_n780), .C1(new_n1032), .C2(new_n775), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT49), .Z(new_n1034));
  AOI211_X1 g0834(.A(new_n1027), .B(new_n1034), .C1(G116), .C2(new_n770), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n766), .A2(new_n844), .B1(new_n778), .B2(new_n355), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G50), .B2(new_n801), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n329), .B1(new_n770), .B2(G97), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n839), .A2(G68), .B1(new_n797), .B2(G77), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n791), .A2(new_n309), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n280), .A2(new_n783), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n756), .B1(new_n1035), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n234), .A2(G45), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n703), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1045), .A2(new_n750), .B1(new_n1046), .B2(new_n747), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n311), .A2(G50), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1048), .A2(KEYINPUT50), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(KEYINPUT50), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n703), .B(new_n473), .C1(new_n214), .C2(new_n202), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1047), .A2(new_n1052), .B1(G107), .B2(new_n208), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n746), .B1(new_n1053), .B2(new_n757), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1044), .B(new_n1054), .C1(new_n691), .C2(new_n1021), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1026), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1025), .A2(new_n1056), .ZN(G393));
  NAND3_X1  g0857(.A1(new_n990), .A2(KEYINPUT111), .A3(new_n992), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT111), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n985), .A2(new_n991), .A3(new_n1059), .A4(new_n692), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(new_n978), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n993), .A2(new_n1061), .A3(new_n701), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n839), .A2(G294), .B1(new_n800), .B2(G303), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n595), .B2(new_n780), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT112), .Z(new_n1065));
  OAI21_X1  g0865(.A(new_n329), .B1(new_n769), .B2(new_n323), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n766), .A2(new_n1029), .B1(new_n775), .B2(new_n999), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT52), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n778), .A2(new_n1005), .B1(new_n785), .B2(new_n763), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1066), .B(new_n1067), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1065), .B(new_n1070), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n800), .A2(new_n1012), .B1(new_n797), .B2(G68), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n845), .B2(new_n766), .C1(new_n311), .C2(new_n762), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n329), .B(new_n1073), .C1(G87), .C2(new_n770), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n792), .A2(G77), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n778), .A2(new_n844), .B1(new_n785), .B2(new_n355), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n806), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n244), .A2(new_n750), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n756), .B(new_n755), .C1(G97), .C2(new_n700), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n746), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT113), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n755), .B2(new_n962), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n744), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1062), .A2(new_n1086), .ZN(G390));
  NAND3_X1  g0887(.A1(new_n822), .A2(new_n737), .A3(new_n683), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n873), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n915), .B1(new_n1089), .B2(new_n930), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n911), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n829), .A2(G330), .A3(new_n822), .A4(new_n930), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n874), .A2(new_n915), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n1092), .C1(new_n912), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT39), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n899), .B2(new_n900), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1095), .B2(new_n926), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1093), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1097), .A2(new_n1098), .B1(new_n911), .B2(new_n1090), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n921), .A2(new_n870), .A3(new_n687), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1094), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n871), .A2(new_n873), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n930), .B1(new_n734), .B2(new_n822), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1103), .B1(new_n1104), .B2(new_n1100), .ZN(new_n1105));
  OAI211_X1 g0905(.A(G330), .B(new_n822), .C1(new_n920), .C2(new_n731), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1089), .B1(new_n870), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1092), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT114), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT114), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1092), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1105), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n917), .A2(new_n674), .A3(new_n936), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n702), .B1(new_n1102), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1102), .B2(new_n1115), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1102), .A2(new_n743), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n746), .B1(new_n280), .B2(new_n833), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n769), .A2(new_n214), .B1(new_n766), .B2(new_n1032), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n247), .B(new_n1120), .C1(G87), .C2(new_n797), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G283), .A2(new_n796), .B1(new_n801), .B2(G116), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n839), .A2(G97), .B1(new_n800), .B2(G107), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1121), .A2(new_n1075), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n785), .A2(new_n850), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n247), .B1(new_n778), .B2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT54), .B(G143), .Z(new_n1128));
  AOI211_X1 g0928(.A(new_n1125), .B(new_n1127), .C1(new_n839), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n792), .A2(G159), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n775), .A2(new_n844), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  INV_X1    g0932(.A(G137), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n783), .A2(new_n1133), .B1(new_n769), .B2(new_n201), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G125), .B2(new_n767), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1124), .A2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1119), .B1(new_n806), .B2(new_n1137), .C1(new_n912), .C2(new_n754), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1117), .A2(new_n1118), .A3(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT119), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT55), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n306), .B(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n299), .B2(new_n680), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n306), .B(KEYINPUT55), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n299), .A2(new_n680), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1143), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1144), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1140), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n935), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n939), .A2(G330), .A3(new_n1151), .A4(new_n934), .ZN(new_n1154));
  AOI211_X1 g0954(.A(KEYINPUT120), .B(new_n916), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n916), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1153), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT120), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n744), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n753), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n767), .A2(G283), .B1(new_n801), .B2(G107), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n357), .B2(new_n769), .C1(new_n309), .C2(new_n762), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n329), .A2(new_n475), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n800), .B2(G97), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n202), .B2(new_n775), .C1(new_n595), .C2(new_n778), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1163), .A2(new_n1166), .A3(new_n1009), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1164), .B(new_n440), .C1(G33), .C2(G41), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT115), .Z(new_n1171));
  NOR2_X1   g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT117), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n762), .A2(new_n1133), .B1(new_n785), .B2(new_n1126), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G125), .B2(new_n796), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n800), .A2(G132), .B1(new_n797), .B2(new_n1128), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n844), .C2(new_n791), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n770), .A2(G159), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1173), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1172), .B2(KEYINPUT117), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n756), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n746), .B1(new_n201), .B2(new_n833), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1161), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1160), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1114), .B1(new_n1102), .B2(new_n1115), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1154), .A2(new_n1153), .A3(new_n916), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n916), .B1(new_n1154), .B2(new_n1153), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1191), .B(KEYINPUT57), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1195), .A2(new_n701), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1191), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1190), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(G375));
  NAND4_X1  g1001(.A1(new_n1113), .A2(new_n1105), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1115), .A2(new_n969), .A3(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G97), .A2(new_n797), .B1(new_n801), .B2(G283), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n323), .B2(new_n762), .C1(new_n1032), .C2(new_n778), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n329), .B1(new_n769), .B2(new_n202), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n783), .A2(new_n595), .B1(new_n766), .B2(new_n772), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1205), .A2(new_n1041), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT121), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n766), .A2(new_n1126), .B1(new_n778), .B2(new_n850), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n329), .B(new_n1210), .C1(new_n278), .C2(new_n770), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n792), .A2(G50), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n839), .A2(G150), .B1(new_n801), .B2(G137), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n800), .A2(new_n1128), .B1(new_n797), .B2(G159), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1208), .B2(KEYINPUT121), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n756), .B1(new_n1209), .B2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n745), .C1(G68), .C2(new_n834), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n870), .B2(new_n753), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1112), .B2(new_n744), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1203), .A2(new_n1220), .ZN(G381));
  OR2_X1    g1021(.A1(new_n1200), .A2(KEYINPUT122), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1025), .A2(new_n811), .A3(new_n1056), .ZN(new_n1223));
  INV_X1    g1023(.A(G384), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G378), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1200), .A2(KEYINPUT122), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1222), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT123), .ZN(G407));
  NAND3_X1  g1030(.A1(new_n1222), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1231));
  OAI211_X1 g1031(.A(G407), .B(G213), .C1(G343), .C2(new_n1231), .ZN(G409));
  AND2_X1   g1032(.A1(new_n935), .A2(new_n1152), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n935), .A2(new_n1152), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1158), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n916), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1157), .A2(new_n1158), .A3(new_n1156), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1188), .B1(new_n1238), .B2(new_n744), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1191), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1195), .A2(new_n701), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G378), .B(new_n1239), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1157), .A2(new_n1156), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1192), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1188), .B1(new_n1244), .B2(new_n744), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1197), .B2(new_n970), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1227), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1242), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n870), .B1(new_n830), .B2(new_n823), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1101), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1250), .A2(new_n1103), .B1(KEYINPUT114), .B2(new_n1108), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1251), .A2(KEYINPUT60), .A3(new_n1113), .A4(new_n1111), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1202), .A2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1252), .A2(new_n1254), .A3(new_n701), .A4(new_n1115), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1255), .A2(G384), .A3(new_n1220), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G384), .B1(new_n1255), .B2(new_n1220), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G213), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(G343), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1248), .A2(new_n1258), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT62), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1260), .A2(G2897), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(KEYINPUT124), .B(new_n1266), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT124), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1255), .A2(new_n1220), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1224), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1255), .A2(G384), .A3(new_n1220), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1266), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1268), .B1(new_n1269), .B2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1238), .A2(new_n969), .A3(new_n1191), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G378), .B1(new_n1277), .B2(new_n1245), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(new_n1200), .B2(G378), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1279), .B2(new_n1260), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1248), .A2(new_n1281), .A3(new_n1258), .A4(new_n1261), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1263), .A2(new_n1264), .A3(new_n1280), .A4(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1248), .A2(new_n1261), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT61), .B1(new_n1286), .B2(new_n1276), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1287), .A2(new_n1263), .A3(KEYINPUT126), .A4(new_n1282), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n811), .B1(new_n1025), .B2(new_n1056), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1223), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(G390), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1062), .B(new_n1086), .C1(new_n1223), .C2(new_n1289), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n995), .A2(new_n1291), .A3(new_n1022), .A4(new_n1292), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  XOR2_X1   g1096(.A(new_n1296), .B(KEYINPUT127), .Z(new_n1297));
  NAND3_X1  g1097(.A1(new_n1285), .A2(new_n1288), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1280), .A2(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1262), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1294), .A2(new_n1264), .A3(new_n1295), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT125), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1300), .B(new_n1302), .C1(new_n1303), .C2(new_n1262), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(G405));
  NOR2_X1   g1105(.A1(new_n1200), .A2(G378), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1242), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(new_n1258), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1309), .B(new_n1296), .ZN(G402));
endmodule


