//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1228, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n211), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n209), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n203), .A2(G50), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n214), .B1(KEYINPUT1), .B2(new_n221), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(new_n222), .ZN(new_n243));
  NAND2_X1  g0043(.A1(G33), .A2(G41), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n246));
  AND2_X1   g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(KEYINPUT68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n245), .A2(new_n246), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT68), .ZN(new_n250));
  OAI21_X1  g0050(.A(G238), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1698), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n257), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n256), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n245), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT13), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n243), .B2(new_n244), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n246), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n208), .B(KEYINPUT64), .C1(G41), .C2(G45), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n252), .A2(new_n262), .A3(new_n263), .A4(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(new_n248), .B2(new_n251), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT13), .B1(new_n271), .B2(new_n261), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(G190), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n222), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G50), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n209), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G77), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n280), .A2(new_n281), .B1(new_n209), .B2(G68), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n275), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT11), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n208), .A2(G20), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT65), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n275), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G68), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n202), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT12), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n283), .A2(new_n284), .ZN(new_n296));
  AND4_X1   g0096(.A1(new_n285), .A2(new_n293), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n273), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n270), .B2(new_n272), .ZN(new_n300));
  OR3_X1    g0100(.A1(new_n298), .A2(KEYINPUT69), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT69), .B1(new_n298), .B2(new_n300), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n297), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n270), .A2(G179), .A3(new_n272), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n270), .B2(new_n272), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n305), .B(new_n306), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n292), .A2(G50), .ZN(new_n314));
  XOR2_X1   g0114(.A(KEYINPUT8), .B(G58), .Z(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(new_n280), .ZN(new_n317));
  OAI21_X1  g0117(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n318));
  INV_X1    g0118(.A(G150), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n277), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n275), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n289), .A2(new_n278), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n314), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n255), .B2(new_n256), .ZN(new_n325));
  AND2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n325), .A2(G223), .B1(new_n328), .B2(G77), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n257), .A2(G222), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(G226), .B2(new_n247), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n323), .A2(KEYINPUT9), .B1(new_n336), .B2(G190), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n314), .A2(new_n321), .A3(new_n322), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT9), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(new_n335), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n338), .A2(new_n339), .B1(new_n340), .B2(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT10), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n323), .B1(new_n307), .B2(new_n340), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(G179), .B2(new_n340), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT66), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n315), .B1(new_n347), .B2(new_n276), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n347), .B2(new_n276), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT15), .B(G87), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n350), .A2(new_n280), .B1(new_n209), .B2(new_n281), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n275), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n288), .A2(G77), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n292), .B2(G77), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n325), .A2(G238), .B1(new_n328), .B2(G107), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n259), .A2(G232), .A3(new_n324), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n332), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n334), .B1(G244), .B2(new_n247), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n356), .B1(new_n299), .B2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(KEYINPUT67), .B1(G190), .B2(new_n363), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT67), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n356), .B(new_n366), .C1(new_n299), .C2(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n362), .A2(new_n307), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n355), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  OR3_X1    g0173(.A1(new_n313), .A2(new_n346), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n255), .A2(new_n209), .A3(new_n256), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT7), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n255), .A2(new_n377), .A3(new_n209), .A4(new_n256), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(G68), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  XNOR2_X1  g0180(.A(G58), .B(G68), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G20), .B1(G159), .B2(new_n276), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n380), .B1(new_n379), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n275), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n315), .A2(new_n288), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n292), .B2(new_n315), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n245), .A2(G232), .A3(new_n246), .ZN(new_n388));
  INV_X1    g0188(.A(G87), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n254), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(G223), .A2(G1698), .ZN(new_n391));
  INV_X1    g0191(.A(G226), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(G1698), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n390), .B1(new_n393), .B2(new_n259), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n269), .B(new_n388), .C1(new_n394), .C2(new_n245), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n299), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(G1698), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(G223), .B2(G1698), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n398), .A2(new_n328), .B1(new_n254), .B2(new_n389), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n332), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(new_n269), .A4(new_n388), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n385), .A2(new_n387), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT71), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n385), .A2(new_n403), .A3(KEYINPUT71), .A4(new_n387), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n395), .A2(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n369), .B2(new_n395), .ZN(new_n411));
  INV_X1    g0211(.A(new_n275), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n379), .A2(new_n382), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT16), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n387), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n411), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT18), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n385), .A2(new_n387), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n411), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n404), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n409), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n374), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(G250), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n428));
  OAI211_X1 g0228(.A(G257), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G294), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n332), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n208), .A2(G45), .ZN(new_n433));
  OR2_X1    g0233(.A1(KEYINPUT5), .A2(G41), .ZN(new_n434));
  NAND2_X1  g0234(.A1(KEYINPUT5), .A2(G41), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n265), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT5), .B(G41), .ZN(new_n438));
  INV_X1    g0238(.A(G45), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n438), .A2(new_n440), .B1(new_n243), .B2(new_n244), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G264), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n432), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT78), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n431), .A2(new_n332), .B1(new_n441), .B2(G264), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT78), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n437), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(G169), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n443), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G179), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n209), .B(G87), .C1(new_n326), .C2(new_n327), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT22), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT24), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  INV_X1    g0256(.A(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(G20), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT73), .B(G116), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n254), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n461), .B2(new_n209), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n453), .A2(new_n454), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n454), .B1(new_n453), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n275), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT25), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n288), .B2(G107), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n288), .A2(new_n466), .A3(G107), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n208), .A2(G33), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n288), .A2(new_n470), .A3(new_n222), .A4(new_n274), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n468), .A2(new_n469), .B1(new_n457), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n451), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n444), .A2(new_n447), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n477), .A2(new_n401), .B1(new_n299), .B2(new_n443), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n478), .B2(new_n474), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n462), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT24), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n453), .A2(new_n454), .A3(new_n462), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n472), .B1(new_n485), .B2(new_n275), .ZN(new_n486));
  AOI21_X1  g0286(.A(G190), .B1(new_n444), .B2(new_n447), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n449), .A2(G200), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n486), .B(KEYINPUT79), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n475), .B1(new_n479), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT74), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n440), .A2(G274), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n433), .A2(G250), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n332), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G244), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n495));
  OAI211_X1 g0295(.A(G238), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(new_n254), .C2(new_n460), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n494), .B1(new_n497), .B2(new_n332), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n491), .B1(new_n499), .B2(new_n401), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n259), .A2(new_n209), .A3(G68), .ZN(new_n501));
  NAND3_X1  g0301(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n209), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n206), .B2(G87), .ZN(new_n504));
  INV_X1    g0304(.A(G97), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n280), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n501), .B(new_n504), .C1(KEYINPUT19), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n275), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n350), .A2(new_n289), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n471), .A2(new_n389), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n499), .A2(G200), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n498), .A2(KEYINPUT74), .A3(G190), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n500), .A2(new_n511), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n508), .B(new_n509), .C1(new_n350), .C2(new_n471), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n498), .A2(new_n369), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(G169), .C2(new_n498), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n514), .A2(new_n517), .A3(KEYINPUT75), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT75), .B1(new_n514), .B2(new_n517), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n209), .C1(G33), .C2(new_n505), .ZN(new_n522));
  INV_X1    g0322(.A(G116), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n275), .B(new_n522), .C1(new_n527), .C2(new_n209), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT20), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n460), .A2(G20), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(KEYINPUT20), .A3(new_n275), .A4(new_n522), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT76), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n290), .A2(new_n534), .A3(G116), .A4(new_n470), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT76), .B1(new_n471), .B2(new_n523), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n531), .ZN(new_n538));
  INV_X1    g0338(.A(G13), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G1), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n533), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n441), .A2(G270), .B1(new_n265), .B2(new_n436), .ZN(new_n543));
  OAI211_X1 g0343(.A(G264), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n544));
  OAI211_X1 g0344(.A(G257), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n255), .A2(G303), .A3(new_n256), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n332), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n307), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n542), .A2(KEYINPUT21), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT21), .B1(new_n542), .B2(new_n549), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n543), .A2(new_n548), .A3(G179), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n530), .A2(new_n532), .B1(new_n540), .B2(new_n538), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n537), .B2(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n543), .A2(new_n548), .A3(G190), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(new_n553), .A3(new_n537), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n299), .B1(new_n543), .B2(new_n548), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT77), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n542), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT77), .ZN(new_n561));
  INV_X1    g0361(.A(new_n558), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n556), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(G244), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n565));
  NOR2_X1   g0365(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G250), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n567), .A2(new_n521), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n566), .ZN(new_n570));
  INV_X1    g0370(.A(new_n565), .ZN(new_n571));
  AND2_X1   g0371(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n245), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n441), .A2(G257), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n437), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n307), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n568), .A2(new_n521), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n572), .B1(new_n257), .B2(G244), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n567), .C1(new_n579), .C2(new_n566), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n576), .B1(new_n580), .B2(new_n332), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n369), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT6), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n505), .A2(new_n457), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n205), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n457), .A2(KEYINPUT6), .A3(G97), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n376), .A2(G107), .A3(new_n378), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n412), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n289), .A2(new_n505), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n471), .B2(new_n505), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n577), .B(new_n582), .C1(new_n590), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n581), .A2(G190), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n590), .A2(new_n592), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n594), .B(new_n595), .C1(new_n299), .C2(new_n581), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n555), .A2(new_n564), .A3(new_n593), .A4(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n427), .A2(new_n490), .A3(new_n520), .A4(new_n597), .ZN(G372));
  NAND2_X1  g0398(.A1(new_n497), .A2(new_n332), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n494), .A2(KEYINPUT80), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n494), .A2(KEYINPUT80), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n307), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n515), .A3(new_n516), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT82), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n451), .A2(new_n474), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n607), .B(KEYINPUT81), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n555), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n602), .A2(G200), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n500), .A2(new_n511), .A3(new_n610), .A4(new_n513), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n604), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n593), .A2(new_n596), .ZN(new_n613));
  AOI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n479), .C2(new_n489), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n606), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n518), .A2(new_n519), .A3(new_n593), .ZN(new_n616));
  XNOR2_X1  g0416(.A(KEYINPUT83), .B(KEYINPUT26), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n612), .A2(new_n593), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT26), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n427), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n345), .ZN(new_n625));
  INV_X1    g0425(.A(new_n312), .ZN(new_n626));
  INV_X1    g0426(.A(new_n372), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n303), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n424), .B1(new_n406), .B2(new_n407), .ZN(new_n629));
  INV_X1    g0429(.A(new_n425), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n423), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n625), .B1(new_n633), .B2(new_n343), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n624), .A2(new_n634), .ZN(G369));
  NAND2_X1  g0435(.A1(new_n540), .A2(new_n209), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(G343), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n490), .B1(new_n486), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n607), .B2(new_n643), .ZN(new_n645));
  INV_X1    g0445(.A(new_n555), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n643), .A2(new_n560), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n555), .A2(new_n564), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n647), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n650), .A2(new_n651), .A3(G330), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n650), .B2(G330), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n645), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT85), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT85), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n608), .A2(new_n642), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n646), .A2(new_n643), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n490), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n657), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n212), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G1), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n225), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n607), .A2(new_n555), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n614), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI22_X1  g0473(.A1(new_n616), .A2(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n614), .A2(KEYINPUT89), .A3(new_n670), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n673), .A2(new_n674), .A3(new_n605), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT90), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(KEYINPUT29), .A4(new_n643), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n676), .A2(KEYINPUT29), .A3(new_n643), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n642), .B1(new_n615), .B2(new_n622), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT90), .B1(new_n680), .B2(KEYINPUT29), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n678), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n498), .A2(new_n445), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT86), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n552), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n498), .A2(new_n445), .A3(KEYINPUT86), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n686), .A2(new_n687), .A3(new_n581), .A4(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  AOI21_X1  g0490(.A(G179), .B1(new_n543), .B2(new_n548), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n602), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n581), .A2(new_n449), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n689), .A2(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT87), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n574), .A2(new_n552), .A3(new_n576), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n697), .A2(KEYINPUT30), .A3(new_n688), .A4(new_n686), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n694), .B2(new_n695), .ZN(new_n699));
  OAI211_X1 g0499(.A(KEYINPUT31), .B(new_n642), .C1(new_n696), .C2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n490), .A2(new_n597), .A3(new_n520), .A4(new_n643), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n689), .A2(new_n690), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n693), .A2(new_n692), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n698), .A3(KEYINPUT88), .A4(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n642), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT88), .B1(new_n694), .B2(new_n698), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n702), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n700), .A2(new_n701), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n683), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n669), .B1(new_n712), .B2(G1), .ZN(G364));
  NOR2_X1   g0513(.A1(new_n652), .A2(new_n653), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n539), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n208), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n664), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n714), .B(new_n719), .C1(G330), .C2(new_n650), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n663), .A2(new_n328), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  XOR2_X1   g0522(.A(G355), .B(KEYINPUT91), .Z(new_n723));
  OAI22_X1  g0523(.A1(new_n722), .A2(new_n723), .B1(G116), .B2(new_n212), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n663), .A2(new_n259), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n225), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n726), .B1(new_n439), .B2(new_n727), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n238), .A2(new_n439), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G13), .A2(G33), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n222), .B1(G20), .B2(new_n307), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n718), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n209), .A2(G190), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n739), .A2(new_n369), .A3(G200), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G311), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n369), .A2(new_n299), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n738), .ZN(new_n744));
  XOR2_X1   g0544(.A(KEYINPUT33), .B(G317), .Z(new_n745));
  OAI22_X1  g0545(.A1(new_n741), .A2(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n209), .A2(new_n401), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n743), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n259), .B(new_n746), .C1(G326), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n747), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n751), .A2(new_n299), .A3(G179), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n751), .A2(new_n369), .A3(G200), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G303), .A2(new_n752), .B1(new_n753), .B2(G322), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n739), .A2(G179), .A3(new_n299), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n755), .A2(G283), .B1(G329), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n209), .B1(new_n756), .B2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G294), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n750), .A2(new_n754), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n753), .A2(G58), .B1(new_n749), .B2(G50), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n740), .A2(KEYINPUT92), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n740), .A2(KEYINPUT92), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n764), .B1(new_n767), .B2(new_n281), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(KEYINPUT93), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n760), .B(KEYINPUT94), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n758), .A2(G159), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  INV_X1    g0573(.A(new_n752), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n774), .A2(new_n389), .B1(new_n744), .B2(new_n202), .ZN(new_n775));
  INV_X1    g0575(.A(new_n755), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n259), .B1(new_n776), .B2(new_n457), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n773), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n769), .A2(new_n771), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n768), .A2(KEYINPUT93), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n763), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n737), .B1(new_n781), .B2(new_n734), .ZN(new_n782));
  INV_X1    g0582(.A(new_n733), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n650), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n720), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NOR2_X1   g0586(.A1(new_n372), .A2(new_n642), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n355), .A2(new_n642), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n368), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(new_n789), .B2(new_n372), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n680), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n718), .B1(new_n791), .B2(new_n710), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n710), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n734), .A2(new_n731), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT95), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n719), .B1(new_n796), .B2(new_n281), .ZN(new_n797));
  INV_X1    g0597(.A(new_n734), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n755), .A2(G87), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n748), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n259), .B(new_n801), .C1(G294), .C2(new_n753), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n774), .A2(new_n457), .B1(new_n757), .B2(new_n742), .ZN(new_n803));
  INV_X1    g0603(.A(new_n744), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G283), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n767), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n527), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n753), .A2(G143), .B1(new_n749), .B2(G137), .ZN(new_n809));
  INV_X1    g0609(.A(G159), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n319), .B2(new_n744), .C1(new_n767), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT34), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n752), .A2(G50), .B1(G132), .B2(new_n758), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n328), .B1(new_n755), .B2(G68), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n201), .C2(new_n760), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n811), .B2(new_n812), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n808), .A2(new_n771), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n797), .B1(new_n798), .B2(new_n818), .C1(new_n790), .C2(new_n732), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n793), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G384));
  INV_X1    g0621(.A(new_n587), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT35), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n523), .B(new_n224), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n824), .A2(KEYINPUT96), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(KEYINPUT96), .B2(new_n824), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT36), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n727), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n278), .A2(G68), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n208), .B(G13), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n626), .A2(new_n643), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT38), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n416), .A2(KEYINPUT97), .A3(new_n417), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT97), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n385), .B2(new_n387), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n639), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n834), .B1(new_n426), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n411), .B1(new_n835), .B2(new_n837), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n838), .A2(new_n841), .A3(new_n406), .A4(new_n407), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT37), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n416), .A2(new_n417), .B1(new_n411), .B2(new_n639), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT37), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n406), .A2(new_n844), .A3(new_n845), .A4(new_n407), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT98), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT98), .ZN(new_n848));
  AND4_X1   g0648(.A1(new_n845), .A2(new_n406), .A3(new_n407), .A4(new_n844), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(new_n842), .C2(KEYINPUT37), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n411), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT97), .B1(new_n416), .B2(new_n417), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n385), .A2(new_n836), .A3(new_n387), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n408), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n845), .B1(new_n856), .B2(new_n838), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n848), .B1(new_n857), .B2(new_n849), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n843), .A2(KEYINPUT98), .A3(new_n846), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n858), .A2(new_n859), .B1(new_n426), .B2(new_n839), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n851), .B1(new_n860), .B2(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n419), .A2(new_n422), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n629), .A2(new_n863), .A3(new_n630), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT38), .B1(new_n864), .B2(new_n838), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n858), .B2(new_n859), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n420), .A2(new_n639), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n844), .A2(new_n404), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n426), .A2(new_n869), .B1(new_n846), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n867), .B1(new_n872), .B2(KEYINPUT38), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT99), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT99), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n846), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n864), .B2(new_n868), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT39), .B1(new_n877), .B2(new_n834), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n851), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT100), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n862), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n862), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n833), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n787), .B1(new_n680), .B2(new_n790), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n297), .A2(new_n643), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n303), .A2(new_n312), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n303), .B2(new_n312), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n891), .A2(new_n861), .B1(new_n863), .B2(new_n640), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n682), .A2(new_n427), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n634), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n790), .B1(new_n888), .B2(new_n889), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT101), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n703), .A2(new_n698), .A3(new_n704), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT88), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n901), .A2(KEYINPUT31), .A3(new_n642), .A4(new_n705), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n701), .A2(new_n708), .A3(new_n898), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n701), .A2(new_n708), .A3(new_n902), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT101), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n897), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n861), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n877), .A2(new_n834), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n908), .B1(new_n851), .B2(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n907), .A2(new_n908), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n905), .A2(new_n903), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n427), .A3(new_n912), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n847), .A2(new_n850), .B1(new_n864), .B2(new_n838), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n866), .B1(new_n914), .B2(new_n834), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n789), .A2(new_n372), .ZN(new_n916));
  INV_X1    g0716(.A(new_n787), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n303), .A2(new_n312), .A3(new_n887), .ZN(new_n919));
  INV_X1    g0719(.A(new_n889), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n912), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n908), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n906), .A2(new_n910), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n427), .A2(new_n912), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n913), .A2(new_n927), .A3(G330), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n896), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n208), .B2(new_n715), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n896), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n831), .B1(new_n930), .B2(new_n931), .ZN(G367));
  OAI211_X1 g0732(.A(new_n593), .B(new_n596), .C1(new_n595), .C2(new_n643), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n593), .B2(new_n643), .ZN(new_n934));
  NOR2_X1   g0734(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n661), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n936), .B(new_n937), .Z(new_n938));
  NAND2_X1  g0738(.A1(new_n661), .A2(new_n934), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT45), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n657), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(new_n657), .A3(new_n940), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n660), .A2(new_n490), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n645), .B2(new_n660), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(new_n714), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n711), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n664), .B(KEYINPUT41), .Z(new_n951));
  OAI21_X1  g0751(.A(new_n716), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n942), .A2(new_n934), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n660), .A2(new_n934), .A3(new_n490), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n593), .B1(new_n933), .B2(new_n607), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n954), .A2(KEYINPUT42), .B1(new_n643), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(KEYINPUT42), .B2(new_n954), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT43), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n643), .A2(new_n511), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n612), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n606), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n957), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n958), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n953), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n952), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n752), .A2(KEYINPUT46), .A3(G116), .ZN(new_n967));
  INV_X1    g0767(.A(new_n753), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n967), .B1(new_n748), .B2(new_n742), .C1(new_n800), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n755), .A2(G97), .ZN(new_n970));
  INV_X1    g0770(.A(G294), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n970), .B1(new_n971), .B2(new_n744), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n259), .B(new_n972), .C1(G317), .C2(new_n758), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n774), .A2(new_n460), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n973), .B1(KEYINPUT46), .B2(new_n974), .C1(new_n457), .C2(new_n760), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n969), .B(new_n975), .C1(G283), .C2(new_n807), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT104), .Z(new_n977));
  INV_X1    g0777(.A(G143), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n968), .A2(new_n319), .B1(new_n748), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n328), .B(new_n979), .C1(G58), .C2(new_n752), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n770), .A2(G68), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n807), .A2(G50), .ZN(new_n982));
  INV_X1    g0782(.A(G137), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n744), .A2(new_n810), .B1(new_n757), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G77), .B2(new_n755), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n977), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n734), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n961), .A2(new_n733), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n735), .B1(new_n212), .B2(new_n350), .C1(new_n726), .C2(new_n234), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n991), .A2(KEYINPUT103), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(KEYINPUT103), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n992), .A2(new_n993), .A3(new_n719), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n966), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(G387));
  NAND2_X1  g0797(.A1(new_n663), .A2(new_n457), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n231), .A2(new_n439), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n315), .A2(new_n278), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT50), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n666), .B(new_n439), .C1(new_n202), .C2(new_n281), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n725), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n998), .B1(new_n666), .B2(new_n722), .C1(new_n999), .C2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n719), .B1(new_n1004), .B2(new_n735), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT105), .Z(new_n1006));
  NOR2_X1   g0806(.A1(new_n645), .A2(new_n783), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n774), .A2(new_n281), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G159), .B2(new_n749), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(new_n259), .A3(new_n970), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n770), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n350), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n753), .A2(G50), .B1(new_n315), .B2(new_n804), .ZN(new_n1013));
  XOR2_X1   g0813(.A(KEYINPUT106), .B(G150), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n202), .B2(new_n741), .C1(new_n757), .C2(new_n1014), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n1010), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n753), .A2(G317), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G322), .A2(new_n749), .B1(new_n804), .B2(G311), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n767), .C2(new_n800), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT48), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(KEYINPUT48), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n752), .A2(G294), .B1(G283), .B2(new_n761), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(KEYINPUT107), .B(KEYINPUT49), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n259), .B1(new_n758), .B2(G326), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n776), .B2(new_n460), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1016), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1006), .B(new_n1007), .C1(new_n734), .C2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n949), .B2(new_n717), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n712), .A2(new_n949), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n664), .B1(new_n711), .B2(new_n948), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(G393));
  INV_X1    g0834(.A(KEYINPUT108), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n944), .A2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(new_n943), .Z(new_n1037));
  OR2_X1    g0837(.A1(new_n934), .A2(new_n783), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n735), .B1(new_n505), .B2(new_n212), .C1(new_n726), .C2(new_n241), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n718), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT51), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n968), .A2(new_n810), .B1(new_n748), .B2(new_n319), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n807), .A2(new_n315), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n744), .A2(new_n278), .B1(new_n757), .B2(new_n978), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G68), .B2(new_n752), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n770), .A2(G77), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n259), .A4(new_n799), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n753), .A2(G311), .B1(new_n749), .B2(G317), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n752), .A2(G283), .B1(G322), .B2(new_n758), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n740), .A2(G294), .B1(new_n804), .B2(G303), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n259), .B1(new_n755), .B2(G107), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n761), .A2(new_n527), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1044), .A2(new_n1048), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1040), .B1(new_n1056), .B2(new_n734), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1037), .A2(new_n717), .B1(new_n1038), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n711), .A2(new_n948), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n665), .B1(new_n945), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1037), .B2(new_n1059), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1058), .A2(new_n1061), .ZN(G390));
  NOR3_X1   g0862(.A1(new_n866), .A2(new_n873), .A3(KEYINPUT99), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n875), .B1(new_n851), .B2(new_n878), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n914), .A2(new_n834), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n867), .B1(new_n1066), .B2(new_n851), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT100), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n862), .A2(new_n880), .A3(new_n881), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n832), .B1(new_n885), .B2(new_n890), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n851), .A2(new_n909), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n832), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n676), .A2(new_n643), .A3(new_n916), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n917), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n890), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n710), .A2(new_n890), .A3(new_n918), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1071), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n882), .A2(new_n883), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1077), .B1(new_n1082), .B2(new_n1070), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n906), .A2(G330), .ZN(new_n1084));
  OAI211_X1 g0884(.A(KEYINPUT109), .B(new_n1081), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1071), .A2(new_n1078), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT109), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1084), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1082), .A2(new_n731), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n795), .A2(new_n315), .ZN(new_n1092));
  INV_X1    g0892(.A(G283), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n776), .A2(new_n202), .B1(new_n1093), .B2(new_n748), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n259), .B(new_n1094), .C1(G87), .C2(new_n752), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n807), .A2(G97), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n968), .A2(new_n523), .B1(new_n757), .B2(new_n971), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G107), .B2(new_n804), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1095), .A2(new_n1047), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n755), .A2(G50), .B1(G125), .B2(new_n758), .ZN(new_n1100));
  INV_X1    g0900(.A(G132), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1100), .B1(new_n983), .B2(new_n744), .C1(new_n1101), .C2(new_n968), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n328), .B(new_n1102), .C1(G128), .C2(new_n749), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n774), .A2(new_n1014), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  XOR2_X1   g0906(.A(KEYINPUT54), .B(G143), .Z(new_n1107));
  NAND2_X1  g0907(.A1(new_n807), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1103), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1011), .A2(new_n810), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1099), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n719), .B(new_n1092), .C1(new_n1111), .C2(new_n734), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1090), .A2(new_n717), .B1(new_n1091), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT111), .ZN(new_n1114));
  AOI211_X1 g0914(.A(KEYINPUT109), .B(new_n1084), .C1(new_n1071), .C2(new_n1078), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1087), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n1081), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n427), .A2(G330), .A3(new_n912), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n894), .A2(new_n634), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n890), .B1(new_n710), .B2(new_n918), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT110), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n1084), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n885), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n912), .A2(G330), .A3(new_n790), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n890), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1124), .A2(new_n1125), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1119), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1114), .B(new_n664), .C1(new_n1117), .C2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1130), .B(KEYINPUT112), .Z(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1090), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1131), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1135));
  OAI21_X1  g0935(.A(KEYINPUT111), .B1(new_n1135), .B2(new_n665), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1113), .B1(new_n1134), .B2(new_n1137), .ZN(G378));
  XNOR2_X1  g0938(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n323), .A2(new_n640), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n343), .A2(new_n345), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n343), .B2(new_n345), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1145), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n1143), .A3(new_n1139), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT115), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1146), .A2(new_n1148), .A3(KEYINPUT115), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n911), .A2(G330), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1149), .ZN(new_n1155));
  INV_X1    g0955(.A(G330), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n925), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n832), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n892), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1154), .B(new_n1157), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1149), .B1(new_n911), .B2(G330), .ZN(new_n1161));
  AND4_X1   g0961(.A1(G330), .A2(new_n923), .A3(new_n924), .A4(new_n1153), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n884), .B(new_n892), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n717), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n753), .A2(G128), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1101), .B2(new_n744), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G125), .B2(new_n749), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n752), .A2(new_n1107), .B1(new_n740), .B2(G137), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(new_n319), .C2(new_n1011), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n755), .A2(G159), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G33), .B(G41), .C1(new_n758), .C2(G124), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n278), .B1(new_n326), .B2(G41), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT114), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n968), .A2(new_n457), .B1(new_n776), .B2(new_n201), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n741), .A2(new_n350), .B1(new_n757), .B2(new_n1093), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1008), .A2(G41), .A3(new_n259), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G116), .A2(new_n749), .B1(new_n804), .B2(G97), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n981), .A4(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT58), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1178), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1176), .B(new_n1186), .C1(new_n1185), .C2(new_n1184), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n734), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n719), .B1(new_n278), .B2(new_n794), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n1153), .C2(new_n732), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1166), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1119), .B1(new_n1090), .B2(new_n1130), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1165), .A2(KEYINPUT57), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n664), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1119), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1117), .B2(new_n1131), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1197), .B2(new_n1165), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1192), .B1(new_n1195), .B2(new_n1198), .ZN(G375));
  OAI22_X1  g0999(.A1(new_n505), .A2(new_n774), .B1(new_n968), .B2(new_n1093), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n259), .B(new_n1200), .C1(G77), .C2(new_n755), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n748), .A2(new_n971), .B1(new_n757), .B2(new_n800), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n527), .B2(new_n804), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n457), .C2(new_n767), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1011), .A2(new_n278), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n328), .B1(new_n755), .B2(G58), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT116), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n740), .A2(G150), .B1(new_n804), .B2(new_n1107), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n752), .A2(G159), .B1(new_n749), .B2(G132), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n753), .A2(G137), .B1(G128), .B2(new_n758), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n1204), .A2(new_n1012), .B1(new_n1205), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n734), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n719), .B1(new_n796), .B2(new_n202), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n1076), .C2(new_n732), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1129), .B2(new_n716), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1119), .A2(new_n1129), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n951), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1217), .B1(new_n1133), .B2(new_n1220), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT117), .Z(G381));
  OR2_X1    g1022(.A1(G375), .A2(G378), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1058), .A2(new_n1061), .A3(new_n820), .A4(new_n1224), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1223), .A2(G387), .A3(G381), .A4(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT118), .ZN(G407));
  NAND2_X1  g1027(.A1(new_n641), .A2(G213), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1223), .A2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT119), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(G407), .A2(G213), .A3(new_n1230), .ZN(G409));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G375), .A2(G378), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT121), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1164), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1160), .A2(new_n1163), .A3(KEYINPUT121), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n717), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1190), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1219), .B(new_n1165), .C1(new_n1135), .C2(new_n1119), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT120), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1136), .B(new_n1132), .C1(new_n1090), .C2(new_n1133), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1197), .A2(KEYINPUT120), .A3(new_n1219), .A4(new_n1165), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1113), .A4(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1233), .A2(new_n1228), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1228), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(G2897), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1119), .A2(new_n1129), .A3(KEYINPUT60), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n664), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT60), .B1(new_n1119), .B2(new_n1129), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1218), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1249), .B1(new_n1251), .B2(KEYINPUT122), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT122), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n1253), .A3(new_n1218), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n820), .B(new_n1216), .C1(new_n1252), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(KEYINPUT122), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1249), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1254), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1258), .B2(new_n1217), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1246), .A2(KEYINPUT123), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1247), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1246), .A2(KEYINPUT123), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1246), .A2(G2897), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1255), .A2(new_n1259), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT61), .B1(new_n1245), .B2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1233), .A2(new_n1228), .A3(new_n1244), .A4(new_n1260), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT124), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(KEYINPUT62), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1269), .A2(KEYINPUT62), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1269), .A2(KEYINPUT62), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1268), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1232), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1275));
  OR3_X1    g1075(.A1(new_n1268), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1276), .A2(KEYINPUT125), .A3(new_n1267), .A4(new_n1270), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  AND2_X1   g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(new_n1224), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G390), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1058), .B(new_n1061), .C1(new_n1224), .C2(new_n1279), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n996), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n996), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1278), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(G387), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(KEYINPUT126), .A3(new_n1283), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1275), .A2(new_n1277), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1268), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1293), .A2(KEYINPUT63), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(KEYINPUT63), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .A4(new_n1267), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1292), .A2(new_n1297), .ZN(G405));
  INV_X1    g1098(.A(new_n1260), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1299), .A2(KEYINPUT127), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1290), .B(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(KEYINPUT127), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1223), .A2(new_n1233), .A3(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1301), .B(new_n1303), .ZN(G402));
endmodule


