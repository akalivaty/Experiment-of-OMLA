

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595;

  NOR2_X1 U325 ( .A1(n372), .A2(n371), .ZN(n373) );
  XNOR2_X1 U326 ( .A(n522), .B(n521), .ZN(n551) );
  XNOR2_X1 U327 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n521) );
  XNOR2_X1 U328 ( .A(KEYINPUT38), .B(n454), .ZN(n484) );
  XNOR2_X1 U329 ( .A(n513), .B(KEYINPUT47), .ZN(n514) );
  INV_X1 U330 ( .A(KEYINPUT24), .ZN(n296) );
  XNOR2_X1 U331 ( .A(n515), .B(n514), .ZN(n520) );
  XNOR2_X1 U332 ( .A(n297), .B(n296), .ZN(n298) );
  INV_X1 U333 ( .A(KEYINPUT93), .ZN(n328) );
  NOR2_X1 U334 ( .A1(n555), .A2(n577), .ZN(n556) );
  XNOR2_X1 U335 ( .A(n299), .B(n298), .ZN(n303) );
  XNOR2_X1 U336 ( .A(n328), .B(KEYINPUT26), .ZN(n329) );
  XNOR2_X1 U337 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n458) );
  XNOR2_X1 U338 ( .A(n330), .B(n329), .ZN(n578) );
  XNOR2_X1 U339 ( .A(n459), .B(n458), .ZN(n508) );
  NAND2_X1 U340 ( .A1(n563), .A2(n562), .ZN(n573) );
  INV_X1 U341 ( .A(G50GAT), .ZN(n455) );
  XNOR2_X1 U342 ( .A(n455), .B(KEYINPUT100), .ZN(n456) );
  XNOR2_X1 U343 ( .A(n457), .B(n456), .ZN(G1331GAT) );
  XNOR2_X1 U344 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n293), .B(KEYINPUT2), .ZN(n349) );
  XOR2_X1 U346 ( .A(G50GAT), .B(G162GAT), .Z(n405) );
  XOR2_X1 U347 ( .A(n349), .B(n405), .Z(n295) );
  NAND2_X1 U348 ( .A1(G228GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U350 ( .A(G141GAT), .B(G22GAT), .Z(n432) );
  XNOR2_X1 U351 ( .A(n432), .B(KEYINPUT22), .ZN(n297) );
  XOR2_X1 U352 ( .A(KEYINPUT88), .B(KEYINPUT23), .Z(n301) );
  XNOR2_X1 U353 ( .A(KEYINPUT87), .B(G204GAT), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U355 ( .A(n303), .B(n302), .Z(n308) );
  XNOR2_X1 U356 ( .A(G106GAT), .B(G78GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n304), .B(G148GAT), .ZN(n441) );
  XOR2_X1 U358 ( .A(G211GAT), .B(KEYINPUT21), .Z(n306) );
  XNOR2_X1 U359 ( .A(G197GAT), .B(G218GAT), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n336) );
  XNOR2_X1 U361 ( .A(n441), .B(n336), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n555) );
  XOR2_X1 U363 ( .A(n555), .B(KEYINPUT28), .Z(n504) );
  XOR2_X1 U364 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n310) );
  XNOR2_X1 U365 ( .A(G134GAT), .B(G190GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U367 ( .A(n311), .B(G99GAT), .Z(n313) );
  XOR2_X1 U368 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(n437), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n318) );
  XNOR2_X1 U371 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n314), .B(KEYINPUT82), .ZN(n346) );
  XOR2_X1 U373 ( .A(G113GAT), .B(n346), .Z(n316) );
  NAND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U376 ( .A(n318), .B(n317), .Z(n327) );
  XNOR2_X1 U377 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n319), .B(G183GAT), .ZN(n320) );
  XOR2_X1 U379 ( .A(n320), .B(KEYINPUT84), .Z(n322) );
  XNOR2_X1 U380 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n340) );
  XOR2_X1 U382 ( .A(KEYINPUT86), .B(G176GAT), .Z(n324) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(G15GAT), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n340), .B(n325), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n562) );
  INV_X1 U387 ( .A(n562), .ZN(n501) );
  NAND2_X1 U388 ( .A1(n501), .A2(n555), .ZN(n330) );
  XOR2_X1 U389 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n332) );
  NAND2_X1 U390 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U392 ( .A(n333), .B(KEYINPUT91), .Z(n338) );
  XOR2_X1 U393 ( .A(G64GAT), .B(G92GAT), .Z(n335) );
  XNOR2_X1 U394 ( .A(G176GAT), .B(G204GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n442) );
  XNOR2_X1 U396 ( .A(n336), .B(n442), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U398 ( .A(G36GAT), .B(G190GAT), .Z(n397) );
  XOR2_X1 U399 ( .A(n339), .B(n397), .Z(n342) );
  XOR2_X1 U400 ( .A(G169GAT), .B(G8GAT), .Z(n419) );
  XNOR2_X1 U401 ( .A(n419), .B(n340), .ZN(n341) );
  XOR2_X1 U402 ( .A(n342), .B(n341), .Z(n549) );
  XNOR2_X1 U403 ( .A(n549), .B(KEYINPUT27), .ZN(n370) );
  XOR2_X1 U404 ( .A(KEYINPUT1), .B(KEYINPUT89), .Z(n348) );
  XOR2_X1 U405 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n344) );
  XNOR2_X1 U406 ( .A(G57GAT), .B(KEYINPUT5), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n360) );
  XOR2_X1 U410 ( .A(G134GAT), .B(KEYINPUT74), .Z(n404) );
  XOR2_X1 U411 ( .A(n404), .B(n349), .Z(n351) );
  NAND2_X1 U412 ( .A1(G225GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n358) );
  XOR2_X1 U414 ( .A(G85GAT), .B(G148GAT), .Z(n353) );
  XNOR2_X1 U415 ( .A(G141GAT), .B(G120GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U417 ( .A(n354), .B(G162GAT), .Z(n356) );
  XOR2_X1 U418 ( .A(G113GAT), .B(G1GAT), .Z(n421) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(n421), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U421 ( .A(n358), .B(n357), .Z(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n553) );
  INV_X1 U423 ( .A(n553), .ZN(n366) );
  OR2_X1 U424 ( .A1(n370), .A2(n366), .ZN(n361) );
  OR2_X1 U425 ( .A1(n578), .A2(n361), .ZN(n368) );
  NOR2_X1 U426 ( .A1(n501), .A2(n549), .ZN(n362) );
  NOR2_X1 U427 ( .A1(n555), .A2(n362), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n363), .B(KEYINPUT25), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n364), .B(KEYINPUT94), .ZN(n365) );
  OR2_X1 U430 ( .A1(n366), .A2(n365), .ZN(n367) );
  AND2_X1 U431 ( .A1(n368), .A2(n367), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n369), .B(KEYINPUT95), .ZN(n372) );
  NOR2_X1 U433 ( .A1(n370), .A2(n553), .ZN(n537) );
  NAND2_X1 U434 ( .A1(n537), .A2(n504), .ZN(n523) );
  NOR2_X1 U435 ( .A1(n523), .A2(n562), .ZN(n371) );
  XOR2_X1 U436 ( .A(KEYINPUT96), .B(n373), .Z(n467) );
  XOR2_X1 U437 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n375) );
  XNOR2_X1 U438 ( .A(G1GAT), .B(KEYINPUT78), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n394) );
  XOR2_X1 U440 ( .A(G155GAT), .B(G211GAT), .Z(n377) );
  XNOR2_X1 U441 ( .A(G22GAT), .B(G8GAT), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U443 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n379) );
  XNOR2_X1 U444 ( .A(G64GAT), .B(KEYINPUT77), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U446 ( .A(n381), .B(n380), .Z(n386) );
  XOR2_X1 U447 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n383) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U450 ( .A(KEYINPUT76), .B(n384), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U452 ( .A(G78GAT), .B(G71GAT), .Z(n388) );
  XNOR2_X1 U453 ( .A(G183GAT), .B(G127GAT), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U455 ( .A(n390), .B(n389), .Z(n392) );
  XOR2_X1 U456 ( .A(G15GAT), .B(KEYINPUT69), .Z(n425) );
  XOR2_X1 U457 ( .A(G57GAT), .B(KEYINPUT13), .Z(n447) );
  XNOR2_X1 U458 ( .A(n425), .B(n447), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U460 ( .A(n394), .B(n393), .ZN(n587) );
  XOR2_X1 U461 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n396) );
  XNOR2_X1 U462 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n395) );
  XNOR2_X1 U463 ( .A(n396), .B(n395), .ZN(n409) );
  XOR2_X1 U464 ( .A(KEYINPUT10), .B(n397), .Z(n399) );
  XOR2_X1 U465 ( .A(G99GAT), .B(G85GAT), .Z(n436) );
  XNOR2_X1 U466 ( .A(G218GAT), .B(n436), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U468 ( .A(KEYINPUT73), .B(G92GAT), .Z(n401) );
  NAND2_X1 U469 ( .A1(G232GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U470 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U471 ( .A(n403), .B(n402), .Z(n407) );
  XNOR2_X1 U472 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n414) );
  XOR2_X1 U475 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n411) );
  XNOR2_X1 U476 ( .A(G43GAT), .B(G29GAT), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U478 ( .A(KEYINPUT68), .B(n412), .Z(n422) );
  INV_X1 U479 ( .A(n422), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n572) );
  XNOR2_X1 U481 ( .A(KEYINPUT36), .B(n572), .ZN(n592) );
  NOR2_X1 U482 ( .A1(n587), .A2(n592), .ZN(n415) );
  NAND2_X1 U483 ( .A1(n467), .A2(n415), .ZN(n416) );
  XNOR2_X1 U484 ( .A(KEYINPUT37), .B(n416), .ZN(n461) );
  XOR2_X1 U485 ( .A(KEYINPUT30), .B(G197GAT), .Z(n418) );
  XNOR2_X1 U486 ( .A(G36GAT), .B(G50GAT), .ZN(n417) );
  XNOR2_X1 U487 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U488 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U489 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U490 ( .A(n424), .B(n423), .ZN(n429) );
  XOR2_X1 U491 ( .A(n425), .B(KEYINPUT29), .Z(n427) );
  NAND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U494 ( .A(n429), .B(n428), .Z(n435) );
  XOR2_X1 U495 ( .A(KEYINPUT70), .B(KEYINPUT65), .Z(n431) );
  XNOR2_X1 U496 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n564) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n451) );
  XOR2_X1 U501 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n439) );
  NAND2_X1 U502 ( .A1(G230GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U504 ( .A(n440), .B(KEYINPUT71), .Z(n444) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n446) );
  INV_X1 U507 ( .A(KEYINPUT33), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n447), .B(KEYINPUT31), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n450) );
  NAND2_X1 U511 ( .A1(n451), .A2(n450), .ZN(n453) );
  OR2_X1 U512 ( .A1(n451), .A2(n450), .ZN(n452) );
  NAND2_X1 U513 ( .A1(n453), .A2(n452), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n564), .A2(n459), .ZN(n470) );
  NAND2_X1 U515 ( .A1(n461), .A2(n470), .ZN(n454) );
  NOR2_X1 U516 ( .A1(n504), .A2(n484), .ZN(n457) );
  INV_X1 U517 ( .A(G92GAT), .ZN(n465) );
  INV_X1 U518 ( .A(n564), .ZN(n579) );
  XOR2_X1 U519 ( .A(n508), .B(KEYINPUT101), .Z(n566) );
  NOR2_X1 U520 ( .A1(n579), .A2(n566), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT102), .ZN(n487) );
  NAND2_X1 U522 ( .A1(n487), .A2(n461), .ZN(n462) );
  XOR2_X1 U523 ( .A(KEYINPUT107), .B(n462), .Z(n503) );
  NOR2_X1 U524 ( .A1(n549), .A2(n503), .ZN(n463) );
  XNOR2_X1 U525 ( .A(KEYINPUT108), .B(n463), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n465), .B(n464), .ZN(G1337GAT) );
  NAND2_X1 U527 ( .A1(n587), .A2(n572), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT16), .ZN(n469) );
  INV_X1 U529 ( .A(n467), .ZN(n468) );
  NOR2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n488) );
  NAND2_X1 U531 ( .A1(n470), .A2(n488), .ZN(n478) );
  NOR2_X1 U532 ( .A1(n553), .A2(n478), .ZN(n472) );
  XNOR2_X1 U533 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  NOR2_X1 U536 ( .A1(n549), .A2(n478), .ZN(n474) );
  XOR2_X1 U537 ( .A(G8GAT), .B(n474), .Z(G1325GAT) );
  NOR2_X1 U538 ( .A1(n501), .A2(n478), .ZN(n476) );
  XNOR2_X1 U539 ( .A(KEYINPUT35), .B(KEYINPUT98), .ZN(n475) );
  XNOR2_X1 U540 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(n477), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n504), .A2(n478), .ZN(n479) );
  XOR2_X1 U543 ( .A(G22GAT), .B(n479), .Z(G1327GAT) );
  NOR2_X1 U544 ( .A1(n484), .A2(n553), .ZN(n481) );
  XNOR2_X1 U545 ( .A(KEYINPUT99), .B(KEYINPUT39), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U547 ( .A(G29GAT), .B(n482), .Z(G1328GAT) );
  NOR2_X1 U548 ( .A1(n484), .A2(n549), .ZN(n483) );
  XOR2_X1 U549 ( .A(G36GAT), .B(n483), .Z(G1329GAT) );
  NOR2_X1 U550 ( .A1(n484), .A2(n501), .ZN(n485) );
  XOR2_X1 U551 ( .A(KEYINPUT40), .B(n485), .Z(n486) );
  XNOR2_X1 U552 ( .A(G43GAT), .B(n486), .ZN(G1330GAT) );
  NAND2_X1 U553 ( .A1(n488), .A2(n487), .ZN(n496) );
  NOR2_X1 U554 ( .A1(n553), .A2(n496), .ZN(n489) );
  XOR2_X1 U555 ( .A(G57GAT), .B(n489), .Z(n490) );
  XNOR2_X1 U556 ( .A(KEYINPUT42), .B(n490), .ZN(G1332GAT) );
  NOR2_X1 U557 ( .A1(n549), .A2(n496), .ZN(n492) );
  XNOR2_X1 U558 ( .A(G64GAT), .B(KEYINPUT103), .ZN(n491) );
  XNOR2_X1 U559 ( .A(n492), .B(n491), .ZN(G1333GAT) );
  NOR2_X1 U560 ( .A1(n501), .A2(n496), .ZN(n494) );
  XNOR2_X1 U561 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n493) );
  XNOR2_X1 U562 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U563 ( .A(G71GAT), .B(n495), .ZN(G1334GAT) );
  NOR2_X1 U564 ( .A1(n504), .A2(n496), .ZN(n498) );
  XNOR2_X1 U565 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n497) );
  XNOR2_X1 U566 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U567 ( .A(G78GAT), .B(n499), .ZN(G1335GAT) );
  NOR2_X1 U568 ( .A1(n553), .A2(n503), .ZN(n500) );
  XOR2_X1 U569 ( .A(G85GAT), .B(n500), .Z(G1336GAT) );
  NOR2_X1 U570 ( .A1(n501), .A2(n503), .ZN(n502) );
  XOR2_X1 U571 ( .A(G99GAT), .B(n502), .Z(G1338GAT) );
  NOR2_X1 U572 ( .A1(n504), .A2(n503), .ZN(n506) );
  XNOR2_X1 U573 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U575 ( .A(G106GAT), .B(n507), .ZN(G1339GAT) );
  OR2_X1 U576 ( .A1(n564), .A2(n508), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n509), .B(KEYINPUT46), .ZN(n512) );
  INV_X1 U578 ( .A(n572), .ZN(n510) );
  NOR2_X1 U579 ( .A1(n587), .A2(n510), .ZN(n511) );
  NAND2_X1 U580 ( .A1(n512), .A2(n511), .ZN(n515) );
  XOR2_X1 U581 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n513) );
  INV_X1 U582 ( .A(n587), .ZN(n570) );
  NOR2_X1 U583 ( .A1(n592), .A2(n570), .ZN(n516) );
  XNOR2_X1 U584 ( .A(KEYINPUT45), .B(n516), .ZN(n517) );
  NAND2_X1 U585 ( .A1(n517), .A2(n564), .ZN(n518) );
  NOR2_X1 U586 ( .A1(n518), .A2(n459), .ZN(n519) );
  NOR2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n522) );
  NOR2_X1 U588 ( .A1(n551), .A2(n523), .ZN(n524) );
  NAND2_X1 U589 ( .A1(n562), .A2(n524), .ZN(n532) );
  NOR2_X1 U590 ( .A1(n564), .A2(n532), .ZN(n525) );
  XOR2_X1 U591 ( .A(G113GAT), .B(n525), .Z(G1340GAT) );
  NOR2_X1 U592 ( .A1(n566), .A2(n532), .ZN(n527) );
  XNOR2_X1 U593 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U595 ( .A(G120GAT), .B(n528), .Z(G1341GAT) );
  NOR2_X1 U596 ( .A1(n570), .A2(n532), .ZN(n530) );
  XNOR2_X1 U597 ( .A(KEYINPUT114), .B(KEYINPUT50), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n531), .Z(G1342GAT) );
  NOR2_X1 U600 ( .A1(n572), .A2(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U603 ( .A(G134GAT), .B(n535), .Z(G1343GAT) );
  NOR2_X1 U604 ( .A1(n551), .A2(n578), .ZN(n536) );
  NAND2_X1 U605 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(KEYINPUT116), .B(n538), .ZN(n546) );
  NOR2_X1 U607 ( .A1(n564), .A2(n546), .ZN(n539) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n539), .Z(G1344GAT) );
  NOR2_X1 U609 ( .A1(n546), .A2(n508), .ZN(n543) );
  XOR2_X1 U610 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n541) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n540) );
  XNOR2_X1 U612 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n543), .B(n542), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n570), .A2(n546), .ZN(n544) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(n544), .Z(n545) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n545), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n546), .A2(n572), .ZN(n548) );
  XNOR2_X1 U618 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n547) );
  XNOR2_X1 U619 ( .A(n548), .B(n547), .ZN(G1347GAT) );
  XNOR2_X1 U620 ( .A(KEYINPUT120), .B(n549), .ZN(n550) );
  NOR2_X1 U621 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n552), .B(KEYINPUT54), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n577) );
  XNOR2_X1 U624 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n556), .A2(n557), .ZN(n561) );
  INV_X1 U626 ( .A(n556), .ZN(n559) );
  INV_X1 U627 ( .A(n557), .ZN(n558) );
  NAND2_X1 U628 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n563) );
  NOR2_X1 U630 ( .A1(n573), .A2(n564), .ZN(n565) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n565), .Z(G1348GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n573), .ZN(n568) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(n569), .ZN(G1349GAT) );
  NOR2_X1 U636 ( .A1(n570), .A2(n573), .ZN(n571) );
  XOR2_X1 U637 ( .A(G183GAT), .B(n571), .Z(G1350GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G190GAT), .B(n576), .Z(G1351GAT) );
  XOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT60), .Z(n581) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n590) );
  NAND2_X1 U644 ( .A1(n590), .A2(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n583) );
  XOR2_X1 U646 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n590), .A2(n459), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(n586), .ZN(G1353GAT) );
  XOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT125), .Z(n589) );
  NAND2_X1 U653 ( .A1(n590), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1354GAT) );
  INV_X1 U655 ( .A(n590), .ZN(n591) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n594) );
  XNOR2_X1 U657 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XOR2_X1 U659 ( .A(G218GAT), .B(n595), .Z(G1355GAT) );
endmodule

