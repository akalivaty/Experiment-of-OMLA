//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G235), .A3(G237), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G101), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n463), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n464), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  AND2_X1   g057(.A1(new_n467), .A2(new_n468), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n472), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n495), .B2(G114), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT68), .ZN(new_n498));
  OAI211_X1 g073(.A(G2104), .B(new_n494), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  XNOR2_X1  g074(.A(new_n499), .B(KEYINPUT69), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n467), .A2(new_n472), .A3(new_n468), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n476), .A2(new_n464), .A3(new_n472), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n502), .B1(new_n506), .B2(new_n503), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n501), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n500), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n515), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n511), .A2(new_n512), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT5), .B(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n522), .A2(G88), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n515), .A2(new_n517), .ZN(new_n528));
  INV_X1    g103(.A(G62), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(KEYINPUT71), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT71), .B1(new_n530), .B2(G651), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n514), .B(new_n526), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(G166));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n528), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n524), .A2(KEYINPUT72), .A3(G63), .A4(G651), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n538), .A2(new_n539), .B1(G51), .B2(new_n513), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n522), .A2(G89), .A3(new_n525), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  XOR2_X1   g120(.A(KEYINPUT73), .B(G90), .Z(new_n546));
  NAND3_X1  g121(.A1(new_n522), .A2(new_n525), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n528), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n513), .A2(G52), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n547), .A2(new_n551), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n528), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G651), .B1(G43), .B2(new_n513), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n522), .A2(new_n525), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n528), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n522), .A2(G91), .A3(new_n525), .ZN(new_n573));
  XNOR2_X1  g148(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n513), .A2(G53), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g150(.A(G53), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n576));
  OR2_X1    g151(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n575), .A2(KEYINPUT75), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT75), .B1(new_n575), .B2(new_n578), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n572), .B(new_n573), .C1(new_n579), .C2(new_n580), .ZN(G299));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n534), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n533), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(new_n531), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n585), .A2(KEYINPUT76), .A3(new_n514), .A4(new_n526), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(G303));
  AND2_X1   g162(.A1(new_n522), .A2(new_n525), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G87), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n524), .A2(G74), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n513), .B2(G49), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n588), .A2(G86), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n528), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G48), .B2(new_n513), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G651), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT78), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  INV_X1    g180(.A(new_n513), .ZN(new_n606));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  OAI221_X1 g182(.A(new_n604), .B1(new_n605), .B2(new_n606), .C1(new_n607), .C2(new_n560), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n522), .A2(G92), .A3(new_n525), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT10), .A4(G92), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n513), .A2(G54), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n524), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(new_n602), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n573), .A2(new_n572), .ZN(new_n623));
  INV_X1    g198(.A(new_n580), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n575), .A2(new_n578), .A3(KEYINPUT75), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n622), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n622), .B1(new_n626), .B2(G868), .ZN(G280));
  XOR2_X1   g203(.A(KEYINPUT79), .B(G559), .Z(new_n629));
  OAI21_X1  g204(.A(new_n619), .B1(G860), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT80), .Z(G148));
  NAND2_X1  g206(.A1(new_n619), .A2(new_n629), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g210(.A1(new_n506), .A2(new_n475), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n485), .A2(G123), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n488), .A2(G135), .ZN(new_n641));
  OR2_X1    g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n642), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n639), .A2(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT82), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2438), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT15), .B(G2435), .Z(new_n657));
  XOR2_X1   g232(.A(new_n656), .B(new_n657), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n654), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT83), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(KEYINPUT17), .B2(new_n667), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n664), .A2(new_n665), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n671), .B(new_n673), .C1(KEYINPUT17), .C2(new_n667), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n667), .B(KEYINPUT85), .Z(new_n675));
  OAI211_X1 g250(.A(new_n670), .B(new_n674), .C1(new_n673), .C2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT86), .B(G2096), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  OR3_X1    g267(.A1(new_n685), .A2(new_n688), .A3(new_n691), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1986), .B(G1996), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1981), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1991), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n696), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  NAND2_X1  g276(.A1(new_n485), .A2(G119), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n488), .A2(G131), .ZN(new_n703));
  NOR2_X1   g278(.A1(G95), .A2(G2105), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(new_n472), .B2(G107), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n702), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G25), .B(new_n706), .S(G29), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT35), .B(G1991), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(G288), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT33), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1976), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n598), .B(KEYINPUT77), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(new_n710), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G6), .B2(new_n710), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT32), .B(G1981), .Z(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n710), .A2(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n710), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n718), .A2(new_n719), .B1(G1971), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(G1971), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n715), .A2(new_n720), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n709), .B1(new_n725), .B2(KEYINPUT34), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n710), .A2(G24), .ZN(new_n727));
  INV_X1    g302(.A(G290), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n710), .ZN(new_n729));
  INV_X1    g304(.A(G1986), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n726), .B(new_n731), .C1(KEYINPUT34), .C2(new_n725), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT88), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n736), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT29), .Z(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n710), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n710), .ZN(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n562), .A2(new_n710), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n710), .B2(G19), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G2084), .ZN(new_n749));
  AND2_X1   g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  NOR2_X1   g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n736), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n753), .B(new_n754), .C1(new_n481), .C2(new_n736), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n748), .A2(G1341), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n741), .A2(new_n745), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n748), .A2(G1341), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n739), .A2(new_n740), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n483), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(G2105), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT26), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n485), .A2(KEYINPUT95), .A3(G129), .ZN(new_n766));
  AOI21_X1  g341(.A(KEYINPUT95), .B1(new_n485), .B2(G129), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n762), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  MUX2_X1   g343(.A(G32), .B(new_n768), .S(G29), .Z(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n755), .A2(new_n749), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT93), .Z(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n619), .A2(new_n710), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G4), .B2(new_n710), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n774), .ZN(new_n778));
  OR2_X1    g353(.A1(G29), .A2(G33), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT25), .Z(new_n781));
  AND2_X1   g356(.A1(new_n476), .A2(new_n464), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n782), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n783));
  INV_X1    g358(.A(G139), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n781), .B1(new_n472), .B2(new_n783), .C1(new_n487), .C2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n779), .B1(new_n785), .B2(new_n736), .ZN(new_n786));
  INV_X1    g361(.A(G2072), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT94), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n736), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n736), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT96), .B(G2078), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT97), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n791), .B(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n644), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G29), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n786), .A2(new_n787), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT31), .B(G11), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT30), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(G28), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(G28), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n800), .A2(new_n801), .A3(new_n736), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n778), .A2(new_n789), .A3(new_n794), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n760), .A2(new_n771), .A3(new_n777), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n710), .A2(G20), .ZN(new_n806));
  OAI211_X1 g381(.A(KEYINPUT23), .B(new_n806), .C1(new_n626), .C2(new_n710), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(KEYINPUT23), .B2(new_n806), .ZN(new_n808));
  INV_X1    g383(.A(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n736), .A2(G26), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT89), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n488), .A2(new_n813), .A3(G140), .ZN(new_n814));
  INV_X1    g389(.A(G140), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT89), .B1(new_n487), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(G104), .A2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n485), .A2(G128), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n821), .A2(KEYINPUT90), .A3(G29), .ZN(new_n822));
  AOI21_X1  g397(.A(KEYINPUT90), .B1(new_n821), .B2(G29), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n812), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT91), .B(G2067), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n805), .A2(new_n810), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n710), .A2(G5), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G171), .B2(new_n710), .ZN(new_n829));
  INV_X1    g404(.A(G1961), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n733), .A2(KEYINPUT88), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n732), .A2(new_n734), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n735), .A2(new_n827), .A3(new_n831), .A4(new_n833), .ZN(G150));
  INV_X1    g409(.A(G150), .ZN(G311));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  INV_X1    g411(.A(G80), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n528), .A2(new_n836), .B1(new_n837), .B2(new_n510), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT98), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n840));
  OAI221_X1 g415(.A(new_n840), .B1(new_n837), .B2(new_n510), .C1(new_n528), .C2(new_n836), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(G651), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n522), .A2(G93), .A3(new_n525), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n513), .A2(G55), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n843), .A2(KEYINPUT99), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT99), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n843), .A2(new_n844), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n843), .A2(KEYINPUT99), .A3(new_n844), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n561), .B1(new_n854), .B2(new_n842), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n561), .B(new_n842), .C1(new_n845), .C2(new_n846), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT39), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n619), .A2(G559), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT38), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n859), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n849), .B1(new_n862), .B2(G860), .ZN(G145));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT102), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(KEYINPUT102), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n865), .B(new_n866), .C1(G118), .C2(new_n472), .ZN(new_n867));
  INV_X1    g442(.A(G130), .ZN(new_n868));
  INV_X1    g443(.A(G142), .ZN(new_n869));
  OAI221_X1 g444(.A(new_n867), .B1(new_n484), .B2(new_n868), .C1(new_n869), .C2(new_n487), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n637), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n706), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n785), .A2(KEYINPUT101), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n821), .A2(G164), .ZN(new_n876));
  INV_X1    g451(.A(G164), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n817), .A2(new_n877), .A3(new_n819), .A4(new_n820), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n768), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n878), .A3(new_n768), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n785), .B(KEYINPUT101), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n883), .A2(new_n879), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n873), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n874), .B1(new_n883), .B2(new_n879), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n880), .A2(new_n884), .A3(new_n881), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n872), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(KEYINPUT103), .A3(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n492), .B(KEYINPUT100), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G160), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n492), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n481), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n644), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n897), .A3(new_n795), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n891), .A2(new_n892), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n872), .B1(new_n888), .B2(new_n889), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n890), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n899), .A2(new_n906), .A3(new_n900), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n899), .B2(new_n900), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT104), .A4(new_n872), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n902), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g489(.A1(new_n618), .A2(new_n626), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  NAND4_X1  g491(.A1(G299), .A2(new_n615), .A3(new_n614), .A4(new_n617), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n618), .A2(KEYINPUT106), .A3(new_n626), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n917), .ZN(new_n921));
  XNOR2_X1  g496(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n920), .A2(KEYINPUT41), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n858), .B(new_n632), .ZN(new_n925));
  MUX2_X1   g500(.A(new_n924), .B(new_n921), .S(new_n925), .Z(new_n926));
  XOR2_X1   g501(.A(new_n926), .B(KEYINPUT42), .Z(new_n927));
  NAND2_X1  g502(.A1(new_n716), .A2(new_n534), .ZN(new_n928));
  NAND2_X1  g503(.A1(G305), .A2(G166), .ZN(new_n929));
  XNOR2_X1  g504(.A(G288), .B(KEYINPUT108), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n928), .B2(new_n929), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n932), .A2(G290), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n929), .ZN(new_n935));
  INV_X1    g510(.A(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n728), .B1(new_n937), .B2(new_n931), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n927), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n927), .A2(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(G868), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G868), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n847), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(G295));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n944), .ZN(G331));
  NAND2_X1  g521(.A1(new_n920), .A2(KEYINPUT41), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n922), .B1(new_n915), .B2(new_n917), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  XNOR2_X1  g526(.A(G171), .B(G286), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(KEYINPUT109), .C1(new_n855), .C2(new_n857), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n952), .B1(new_n855), .B2(new_n857), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n847), .A2(new_n562), .ZN(new_n956));
  XNOR2_X1  g531(.A(G286), .B(G301), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n957), .A3(new_n856), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n950), .A2(new_n951), .A3(new_n953), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n953), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n948), .B1(new_n920), .B2(KEYINPUT41), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT110), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n954), .A2(new_n921), .A3(new_n958), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n966));
  OAI21_X1  g541(.A(G290), .B1(new_n932), .B2(new_n933), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n937), .A2(new_n728), .A3(new_n931), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n965), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n966), .B1(new_n965), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n954), .A2(new_n958), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n961), .A2(new_n921), .B1(new_n924), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G37), .B1(new_n939), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT43), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n924), .A2(new_n973), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n961), .A2(new_n921), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n969), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n977), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n984), .B(new_n975), .C1(new_n970), .C2(new_n971), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI211_X1 g564(.A(KEYINPUT112), .B(KEYINPUT44), .C1(new_n985), .C2(new_n986), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n982), .B1(new_n989), .B2(new_n990), .ZN(G397));
  AND3_X1   g566(.A1(new_n501), .A2(new_n505), .A3(new_n507), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT69), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n499), .B(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n500), .B2(new_n508), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT113), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT114), .B(G40), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n473), .A2(new_n480), .A3(new_n1003), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1005), .A2(G1996), .A3(new_n768), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1005), .B(KEYINPUT116), .Z(new_n1007));
  XNOR2_X1  g582(.A(new_n821), .B(G2067), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n768), .A2(G1996), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1006), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n706), .A2(new_n708), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n706), .A2(new_n708), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1007), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1005), .A2(G1986), .A3(G290), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1005), .A2(new_n730), .A3(new_n728), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT115), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT45), .B(new_n999), .C1(new_n500), .C2(new_n508), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1004), .B1(new_n998), .B2(new_n1000), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1021), .B1(new_n1026), .B2(G2078), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n473), .A2(new_n480), .A3(new_n1003), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n999), .C1(new_n500), .C2(new_n508), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n830), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1021), .A2(G2078), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1025), .A2(new_n1022), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1027), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G171), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1032), .A2(G2084), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1029), .B1(KEYINPUT45), .B2(new_n995), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1022), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n744), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G8), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G286), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1043), .B(new_n1044), .C1(new_n1045), .C2(KEYINPUT51), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT51), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1047));
  OAI211_X1 g622(.A(G8), .B(new_n1047), .C1(new_n1042), .C2(G286), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1046), .B(new_n1048), .C1(G168), .C2(new_n1043), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1037), .B1(new_n1049), .B2(KEYINPUT62), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1971), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1032), .A2(G2090), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(G303), .B2(G8), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  AOI211_X1 g631(.A(KEYINPUT55), .B(new_n1056), .C1(new_n583), .C2(new_n586), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(G8), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1004), .A2(new_n1000), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n1056), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n712), .A2(G1976), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT52), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n598), .A2(G1981), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n598), .A2(G1981), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1070), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(KEYINPUT49), .A3(new_n1068), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n1073), .A3(new_n1063), .ZN(new_n1074));
  INV_X1    g649(.A(G1976), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1063), .A2(new_n1064), .A3(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1066), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1059), .A2(new_n1061), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT125), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1059), .A2(new_n1061), .A3(new_n1081), .A4(new_n1078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1050), .B(new_n1083), .C1(KEYINPUT62), .C2(new_n1049), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1042), .A2(G8), .A3(G168), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1085), .A2(KEYINPUT63), .A3(new_n1078), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1078), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1074), .A2(new_n1075), .A3(new_n712), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1063), .B1(new_n1094), .B2(new_n1070), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT118), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1099), .B(new_n1096), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1084), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G40), .ZN(new_n1102));
  XOR2_X1   g677(.A(new_n479), .B(KEYINPUT123), .Z(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(G2105), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1002), .A2(new_n473), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1002), .A2(KEYINPUT124), .A3(new_n473), .A4(new_n1104), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1107), .A2(new_n1024), .A3(new_n1034), .A4(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(new_n1027), .A3(new_n1033), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G171), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(KEYINPUT54), .C1(G171), .C2(new_n1036), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1037), .B1(new_n1110), .B2(G171), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1112), .A2(new_n1083), .A3(new_n1115), .A4(new_n1049), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1032), .A2(new_n809), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1032), .A2(KEYINPUT119), .A3(new_n809), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1024), .A2(new_n1025), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n575), .A2(new_n578), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n573), .A2(new_n1125), .A3(new_n572), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT57), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n626), .B1(KEYINPUT120), .B2(new_n1126), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(KEYINPUT57), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1124), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1120), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT119), .B1(new_n1032), .B2(new_n809), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1123), .B(new_n1130), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(KEYINPUT61), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1135), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1130), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1062), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT58), .B(G1341), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1026), .B2(G1996), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n562), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT59), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1147), .A3(new_n562), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1136), .A2(new_n1140), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT121), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1136), .A2(new_n1140), .A3(new_n1149), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1032), .A2(new_n774), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(G2067), .B2(new_n1141), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1156), .B2(new_n618), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n618), .A2(new_n1156), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1151), .A2(new_n1153), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1138), .A2(new_n618), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1139), .B1(new_n1161), .B2(new_n1155), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1116), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1020), .B1(new_n1101), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1007), .B1(new_n768), .B2(new_n1008), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1005), .A2(G1996), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT46), .Z(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT47), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n821), .A2(G2067), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1007), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1016), .B(KEYINPUT48), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n1015), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1169), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1164), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g751(.A1(new_n913), .A2(new_n700), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n679), .A2(G319), .A3(new_n680), .ZN(new_n1179));
  XNOR2_X1  g753(.A(new_n1179), .B(KEYINPUT126), .ZN(new_n1180));
  NAND4_X1  g754(.A1(new_n1178), .A2(new_n661), .A3(new_n987), .A4(new_n1180), .ZN(G225));
  INV_X1    g755(.A(G225), .ZN(G308));
endmodule


