//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND3_X1   g0009(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n210));
  AOI21_X1  g0010(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n209), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT67), .Z(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n221), .A2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT69), .ZN(new_n241));
  XOR2_X1   g0041(.A(G58), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G169), .ZN(new_n248));
  OR2_X1    g0048(.A1(KEYINPUT71), .A2(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT71), .A2(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G45), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(G41), .A3(new_n250), .ZN(new_n252));
  AND2_X1   g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n251), .A2(new_n252), .A3(G238), .A4(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(new_n253), .B2(new_n254), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT70), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT70), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n258), .B(new_n259), .C1(new_n264), .C2(G45), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G226), .A2(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G232), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G1698), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n268), .A2(new_n271), .B1(G33), .B2(G97), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n254), .B1(new_n210), .B2(new_n211), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n256), .B(new_n265), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G97), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n267), .A2(G1698), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G226), .B2(G1698), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n276), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n273), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT13), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(new_n256), .A4(new_n265), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n248), .B1(new_n275), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT14), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n275), .A2(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(G179), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n288), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT78), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n287), .A2(KEYINPUT78), .A3(new_n288), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G1), .A2(G13), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT65), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G20), .A2(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G50), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT77), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n213), .A2(G33), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n306), .A2(new_n202), .B1(new_n213), .B2(G68), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n302), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT11), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT71), .A2(G1), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT71), .A2(G1), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n311), .A2(new_n312), .A3(new_n213), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n302), .B1(G13), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n313), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(G68), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n308), .A2(new_n309), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n249), .A2(G13), .A3(G20), .A4(new_n250), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n217), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT12), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n310), .A2(new_n316), .A3(new_n317), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n296), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n289), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G190), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n289), .A2(G200), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n331));
  INV_X1    g0131(.A(G226), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n265), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n271), .A2(G222), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n271), .A2(G1698), .ZN(new_n338));
  XOR2_X1   g0138(.A(KEYINPUT72), .B(G223), .Z(new_n339));
  OAI221_X1 g0139(.A(new_n337), .B1(new_n202), .B2(new_n271), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n283), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n335), .A2(KEYINPUT73), .A3(new_n290), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n303), .A2(G150), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT8), .B(G58), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n343), .B1(new_n201), .B2(new_n213), .C1(new_n344), .C2(new_n306), .ZN(new_n345));
  INV_X1    g0145(.A(G50), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n345), .A2(new_n302), .B1(new_n346), .B2(new_n319), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n314), .A2(G50), .A3(new_n315), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n342), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n334), .B1(new_n283), .B2(new_n340), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT73), .B1(new_n351), .B2(G169), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n290), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n344), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n213), .B2(new_n202), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT75), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT15), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(G87), .ZN(new_n362));
  INV_X1    g0162(.A(G87), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(KEYINPUT15), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n360), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(KEYINPUT15), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(G87), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT75), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n306), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n302), .B1(new_n359), .B2(new_n370), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n313), .A2(new_n302), .A3(new_n202), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n202), .B2(new_n319), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n271), .A2(G232), .A3(new_n336), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n281), .A2(G107), .ZN(new_n376));
  INV_X1    g0176(.A(G238), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n375), .B(new_n376), .C1(new_n338), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n283), .ZN(new_n379));
  INV_X1    g0179(.A(G244), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n331), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n265), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n374), .B1(new_n383), .B2(G190), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n378), .A2(new_n283), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n265), .B1(new_n331), .B2(new_n380), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n248), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n379), .A2(new_n290), .A3(new_n265), .A4(new_n381), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n374), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n341), .A2(G190), .A3(new_n265), .A4(new_n333), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n349), .A2(KEYINPUT9), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n349), .A2(KEYINPUT9), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n397), .A2(new_n398), .B1(new_n351), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT10), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n393), .B(KEYINPUT76), .ZN(new_n402));
  INV_X1    g0202(.A(new_n398), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n335), .A2(new_n341), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n403), .A2(new_n396), .B1(G200), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT10), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI211_X1 g0207(.A(new_n354), .B(new_n392), .C1(new_n401), .C2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G223), .A2(G1698), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n332), .B2(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n271), .ZN(new_n411));
  INV_X1    g0211(.A(G33), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n363), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n283), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n331), .A2(new_n267), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(new_n265), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n248), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n414), .A2(new_n415), .A3(new_n290), .A4(new_n265), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT7), .B1(new_n281), .B2(new_n213), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT7), .ZN(new_n421));
  NOR4_X1   g0221(.A1(new_n279), .A2(new_n280), .A3(new_n421), .A4(G20), .ZN(new_n422));
  OAI21_X1  g0222(.A(G68), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(G58), .B(G68), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(G20), .B1(G159), .B2(new_n303), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(KEYINPUT16), .A3(new_n425), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n302), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n315), .A2(new_n355), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n431), .A2(KEYINPUT79), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n318), .A2(new_n212), .A3(new_n301), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n431), .B2(KEYINPUT79), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n432), .A2(new_n434), .B1(new_n319), .B2(new_n344), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n419), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n438));
  INV_X1    g0238(.A(new_n436), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n416), .A2(G200), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n414), .A2(new_n415), .A3(G190), .A4(new_n265), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(KEYINPUT17), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n419), .A2(new_n436), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n430), .A2(new_n435), .A3(new_n440), .A4(new_n441), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT17), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n438), .A2(new_n443), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n419), .A2(new_n436), .A3(new_n444), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n444), .B1(new_n419), .B2(new_n436), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n446), .B(KEYINPUT17), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT80), .ZN(new_n456));
  AND4_X1   g0256(.A1(new_n330), .A2(new_n408), .A3(new_n451), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(G250), .A2(G1698), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(G257), .B2(new_n336), .ZN(new_n460));
  INV_X1    g0260(.A(G294), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n460), .A2(new_n281), .B1(new_n412), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n249), .A2(new_n463), .A3(G45), .A4(new_n250), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT5), .B1(new_n261), .B2(new_n263), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n283), .A2(new_n462), .B1(new_n466), .B2(new_n258), .ZN(new_n467));
  OAI211_X1 g0267(.A(G264), .B(new_n255), .C1(new_n464), .C2(new_n465), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT87), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  OAI211_X1 g0271(.A(G179), .B(new_n467), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT88), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n462), .A2(new_n283), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n262), .A2(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n260), .A2(KEYINPUT70), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G45), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n311), .A2(new_n312), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n478), .A2(new_n480), .A3(new_n258), .A4(new_n463), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n474), .A2(new_n468), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G169), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n472), .A2(new_n473), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n473), .B1(new_n472), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n318), .A2(G107), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n486), .A2(KEYINPUT25), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(KEYINPUT25), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n249), .A2(G33), .A3(new_n250), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n318), .A2(new_n212), .A3(new_n490), .A4(new_n301), .ZN(new_n491));
  INV_X1    g0291(.A(G107), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n213), .B(G87), .C1(new_n279), .C2(new_n280), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT22), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT22), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n271), .A2(new_n498), .A3(new_n213), .A4(G87), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G116), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n306), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n213), .B2(G107), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n492), .A2(KEYINPUT23), .A3(G20), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT24), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n500), .A2(new_n509), .A3(new_n506), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n495), .B1(new_n511), .B2(new_n302), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n484), .A2(new_n485), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G244), .B(new_n336), .C1(new_n279), .C2(new_n280), .ZN(new_n514));
  NOR2_X1   g0314(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n515), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n271), .A2(G244), .A3(new_n336), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n516), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n283), .ZN(new_n522));
  OAI211_X1 g0322(.A(G257), .B(new_n255), .C1(new_n464), .C2(new_n465), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n523), .A2(new_n481), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n248), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  AND2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G97), .A2(G107), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n492), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(G97), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT81), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT6), .A2(G97), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n303), .A2(G77), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n421), .B1(new_n271), .B2(G20), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n492), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n302), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n319), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n491), .B2(new_n543), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n522), .A2(new_n524), .A3(new_n290), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n526), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(G107), .B1(new_n420), .B2(new_n422), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(new_n536), .A3(new_n537), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n545), .B1(new_n551), .B2(new_n302), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n522), .A2(new_n524), .A3(G190), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n523), .A2(new_n481), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n283), .B2(new_n521), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n552), .B(new_n553), .C1(new_n399), .C2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n318), .B1(new_n365), .B2(new_n368), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n529), .A2(new_n363), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT19), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT83), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT83), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT19), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n276), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n558), .B1(new_n563), .B2(G20), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n271), .A2(new_n213), .A3(G68), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n560), .B(new_n562), .C1(new_n306), .C2(new_n543), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n557), .B1(new_n567), .B2(new_n302), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT75), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT75), .B1(new_n366), .B2(new_n367), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n314), .A2(new_n571), .A3(KEYINPUT84), .A4(new_n490), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT84), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n491), .B2(new_n369), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n480), .A2(new_n258), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n251), .A2(G250), .A3(new_n255), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G116), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n377), .A2(new_n336), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n380), .A2(G1698), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n582), .C1(new_n279), .C2(new_n280), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n273), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n290), .ZN(new_n586));
  NOR2_X1   g0386(.A1(G238), .A2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n380), .B2(G1698), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n271), .B1(G33), .B2(G116), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n578), .B(new_n577), .C1(new_n589), .C2(new_n273), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n248), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n576), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n585), .A2(G190), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(G200), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n314), .A2(G87), .A3(new_n490), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n593), .A2(new_n568), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n549), .A2(new_n556), .A3(new_n592), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n482), .A2(G190), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n399), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n500), .A2(new_n509), .A3(new_n506), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n509), .B1(new_n500), .B2(new_n506), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n302), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n493), .B1(new_n487), .B2(new_n488), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n513), .A2(new_n597), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(G257), .B(new_n336), .C1(new_n279), .C2(new_n280), .ZN(new_n609));
  OAI211_X1 g0409(.A(G264), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n269), .A2(G303), .A3(new_n270), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n283), .ZN(new_n613));
  OAI211_X1 g0413(.A(G270), .B(new_n255), .C1(new_n464), .C2(new_n465), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n614), .A2(KEYINPUT85), .A3(new_n481), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT85), .B1(new_n614), .B2(new_n481), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT86), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT86), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n619), .B(new_n613), .C1(new_n615), .C2(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G200), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n314), .A2(G116), .A3(new_n490), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n319), .A2(new_n501), .ZN(new_n624));
  AOI21_X1  g0424(.A(G20), .B1(G33), .B2(G283), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n412), .A2(G97), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n625), .A2(new_n626), .B1(G20), .B2(new_n501), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT20), .B1(new_n627), .B2(new_n302), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n627), .A2(new_n302), .A3(KEYINPUT20), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n623), .B(new_n624), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n618), .A2(G190), .A3(new_n620), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n622), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n248), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n614), .A2(new_n481), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT85), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n614), .A2(new_n481), .A3(KEYINPUT85), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n619), .B1(new_n639), .B2(new_n613), .ZN(new_n640));
  INV_X1    g0440(.A(new_n620), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n634), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT21), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n290), .B1(new_n612), .B2(new_n283), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n639), .A2(new_n630), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n630), .A2(KEYINPUT21), .A3(G169), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n621), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n633), .A2(new_n644), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n458), .A2(new_n608), .A3(new_n650), .ZN(G372));
  INV_X1    g0451(.A(new_n391), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n324), .B1(new_n328), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n455), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n454), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n401), .A2(new_n407), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n354), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n592), .A2(new_n596), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n658), .B2(new_n549), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT89), .B1(new_n590), .B2(new_n248), .ZN(new_n660));
  OAI211_X1 g0460(.A(KEYINPUT89), .B(new_n248), .C1(new_n579), .C2(new_n584), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n576), .B(new_n586), .C1(new_n660), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n576), .A2(new_n586), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n662), .A2(new_n660), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n596), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT90), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n663), .A2(new_n669), .A3(new_n596), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n549), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n664), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n549), .B(new_n556), .C1(new_n600), .C2(new_n605), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n668), .B2(new_n670), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n472), .A2(new_n483), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n605), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n644), .A2(new_n649), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n657), .B1(new_n458), .B2(new_n681), .ZN(G369));
  OAI21_X1  g0482(.A(new_n648), .B1(new_n640), .B2(new_n641), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n646), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT21), .B1(new_n621), .B2(new_n634), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n311), .A2(new_n312), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n213), .A2(G13), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(new_n691), .A3(new_n688), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n686), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n485), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n472), .A2(new_n473), .A3(new_n483), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n605), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n606), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n695), .B(KEYINPUT91), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n701), .B(new_n702), .C1(new_n512), .C2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n513), .A2(new_n697), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n704), .A2(KEYINPUT92), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT92), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n698), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(new_n605), .A3(new_n676), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n706), .A2(new_n707), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n703), .A2(new_n631), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n684), .B2(new_n685), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n650), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n710), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n207), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n264), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n558), .A2(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n219), .B2(new_n720), .ZN(new_n723));
  XOR2_X1   g0523(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n724));
  XNOR2_X1  g0524(.A(new_n723), .B(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n675), .A2(new_n678), .ZN(new_n726));
  INV_X1    g0526(.A(new_n549), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n663), .A2(new_n669), .A3(new_n596), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n669), .B1(new_n663), .B2(new_n596), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n727), .B(new_n672), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n663), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n552), .B1(new_n248), .B2(new_n525), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n592), .A3(new_n548), .A4(new_n596), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n731), .B1(new_n733), .B2(KEYINPUT26), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n703), .B1(new_n726), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n644), .A2(new_n701), .A3(new_n649), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n731), .B1(new_n675), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n727), .B(KEYINPUT26), .C1(new_n728), .C2(new_n729), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n733), .A2(new_n672), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(KEYINPUT95), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT95), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n733), .A2(new_n744), .A3(new_n672), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(KEYINPUT29), .A3(new_n703), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n738), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n585), .A2(new_n474), .A3(new_n645), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n468), .B(new_n469), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(new_n639), .A3(new_n751), .A4(new_n555), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT30), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n585), .A2(new_n474), .A3(new_n645), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n525), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n756), .A2(KEYINPUT30), .A3(new_n751), .A4(new_n639), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n599), .A2(new_n290), .A3(new_n525), .A4(new_n590), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n620), .B2(new_n618), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n697), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT31), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT94), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n607), .A2(new_n686), .A3(new_n633), .A4(new_n703), .ZN(new_n766));
  OAI211_X1 g0566(.A(KEYINPUT31), .B(new_n697), .C1(new_n758), .C2(new_n760), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n761), .A2(KEYINPUT94), .A3(new_n762), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n765), .A2(new_n766), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n769), .A2(G330), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n749), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT96), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n725), .B1(new_n772), .B2(G1), .ZN(G364));
  NOR2_X1   g0573(.A1(new_n714), .A2(G330), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT97), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n259), .B1(new_n688), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n719), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n775), .A2(new_n715), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n213), .B1(KEYINPUT99), .B2(new_n248), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(KEYINPUT99), .B2(new_n248), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n299), .A2(new_n300), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n213), .A2(G179), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G159), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT32), .ZN(new_n791));
  INV_X1    g0591(.A(G190), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n785), .A2(new_n792), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n213), .A2(new_n290), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n795), .A2(G190), .A3(new_n399), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n791), .B1(new_n492), .B2(new_n793), .C1(new_n217), .C2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n794), .A2(G190), .A3(G200), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n290), .A2(new_n399), .A3(G190), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n800), .A2(G50), .B1(G97), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n363), .B2(new_n804), .C1(KEYINPUT32), .C2(new_n790), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n794), .A2(new_n786), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n794), .A2(G190), .A3(new_n399), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n271), .B1(new_n806), .B2(new_n202), .C1(new_n216), .C2(new_n807), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n798), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n281), .B1(new_n806), .B2(new_n810), .C1(new_n811), .C2(new_n807), .ZN(new_n812));
  INV_X1    g0612(.A(new_n787), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n813), .A2(KEYINPUT101), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(KEYINPUT101), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n812), .B1(new_n817), .B2(G329), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n799), .B(KEYINPUT100), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G326), .ZN(new_n821));
  INV_X1    g0621(.A(new_n802), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n461), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  INV_X1    g0624(.A(G303), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n824), .A2(new_n793), .B1(new_n804), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT33), .B(G317), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n823), .B(new_n826), .C1(new_n796), .C2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n818), .A2(new_n821), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n809), .B1(KEYINPUT102), .B2(new_n829), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n829), .A2(KEYINPUT102), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n784), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n784), .ZN(new_n833));
  NOR2_X1   g0633(.A1(G13), .A2(G33), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(G20), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n271), .A2(new_n207), .ZN(new_n838));
  INV_X1    g0638(.A(G355), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n838), .A2(new_n839), .B1(G116), .B2(new_n207), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT98), .Z(new_n841));
  AND2_X1   g0641(.A1(new_n243), .A2(G45), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n718), .A2(new_n271), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(G45), .B2(new_n219), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n841), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n779), .B(new_n832), .C1(new_n837), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n836), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n714), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n780), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  AOI22_X1  g0650(.A1(new_n382), .A2(new_n248), .B1(new_n371), .B2(new_n373), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT104), .B1(new_n851), .B2(new_n390), .ZN(new_n852));
  AND4_X1   g0652(.A1(KEYINPUT104), .A2(new_n389), .A3(new_n374), .A4(new_n390), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n384), .A2(new_n385), .B1(new_n697), .B2(new_n374), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT105), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n652), .A2(new_n856), .A3(new_n697), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT105), .B1(new_n391), .B2(new_n703), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n854), .A2(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n703), .B(new_n860), .C1(new_n726), .C2(new_n735), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT106), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n680), .A2(KEYINPUT106), .A3(new_n703), .A4(new_n860), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n863), .A2(new_n864), .B1(new_n736), .B2(new_n859), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n779), .B1(new_n865), .B2(new_n770), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n770), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n859), .A2(new_n834), .ZN(new_n869));
  INV_X1    g0669(.A(new_n807), .ZN(new_n870));
  INV_X1    g0670(.A(new_n806), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n870), .A2(G143), .B1(new_n871), .B2(G159), .ZN(new_n872));
  INV_X1    g0672(.A(G137), .ZN(new_n873));
  INV_X1    g0673(.A(G150), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n872), .B1(new_n873), .B2(new_n799), .C1(new_n874), .C2(new_n797), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT34), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n817), .A2(G132), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n822), .A2(new_n216), .B1(new_n804), .B2(new_n346), .ZN(new_n880));
  INV_X1    g0680(.A(new_n793), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n281), .B(new_n880), .C1(G68), .C2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n817), .A2(G311), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n363), .A2(new_n793), .B1(new_n804), .B2(new_n492), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(G283), .B2(new_n796), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n281), .B1(new_n807), .B2(new_n461), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(G116), .B2(new_n871), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n800), .A2(G303), .B1(G97), .B2(new_n802), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n884), .A2(new_n886), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n784), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n833), .A2(new_n834), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT103), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n779), .B(new_n891), .C1(new_n202), .C2(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n867), .A2(new_n868), .B1(new_n869), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(G384));
  OR2_X1    g0697(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n898), .A2(G116), .A3(new_n214), .A4(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(KEYINPUT107), .B(KEYINPUT36), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n900), .B(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n219), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(G77), .C1(new_n216), .C2(new_n217), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n346), .A2(G68), .ZN(new_n905));
  AOI211_X1 g0705(.A(G13), .B(new_n687), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  INV_X1    g0709(.A(new_n693), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n436), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n454), .B2(new_n455), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n437), .A2(new_n911), .A3(new_n446), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n437), .A2(new_n911), .A3(KEYINPUT37), .A4(new_n446), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n909), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n911), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n449), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n920), .A2(KEYINPUT38), .A3(new_n916), .A4(new_n915), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n597), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n923), .A2(new_n701), .A3(new_n702), .A4(new_n703), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n763), .B(new_n767), .C1(new_n650), .C2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n291), .ZN(new_n926));
  INV_X1    g0726(.A(new_n295), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT78), .B1(new_n287), .B2(new_n288), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n322), .B(new_n697), .C1(new_n929), .C2(new_n329), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n697), .A2(new_n322), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n328), .B(new_n931), .C1(new_n296), .C2(new_n323), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n859), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n908), .B1(new_n922), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n918), .A2(new_n921), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n936), .A2(KEYINPUT40), .A3(new_n925), .A4(new_n933), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT110), .Z(new_n939));
  INV_X1    g0739(.A(new_n925), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n939), .A2(new_n458), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n939), .B1(new_n458), .B2(new_n940), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n941), .A2(G330), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n454), .A2(new_n910), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT109), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n946), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n936), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n918), .A2(new_n921), .A3(KEYINPUT109), .A4(KEYINPUT39), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n324), .A2(new_n703), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n944), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n854), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n703), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT108), .ZN(new_n958));
  INV_X1    g0758(.A(new_n864), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n697), .B1(new_n673), .B2(new_n679), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT106), .B1(new_n960), .B2(new_n860), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n958), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n930), .A2(new_n932), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n936), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n738), .A2(new_n457), .A3(new_n748), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n657), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n965), .B(new_n967), .Z(new_n968));
  OAI22_X1  g0768(.A1(new_n943), .A2(new_n968), .B1(new_n687), .B2(new_n688), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n943), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n907), .B1(new_n969), .B2(new_n970), .ZN(G367));
  NAND2_X1  g0771(.A1(new_n727), .A2(new_n697), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n549), .B(new_n556), .C1(new_n552), .C2(new_n703), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n716), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT112), .Z(new_n976));
  NAND2_X1  g0776(.A1(new_n568), .A2(new_n595), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n697), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n728), .B2(new_n729), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n731), .A2(new_n977), .A3(new_n697), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n976), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n976), .A2(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n974), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n708), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n549), .B1(new_n701), .B2(new_n973), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n991), .A2(KEYINPUT42), .B1(new_n703), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT113), .Z(new_n997));
  NOR2_X1   g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n989), .B(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n719), .B(KEYINPUT41), .Z(new_n1000));
  INV_X1    g0800(.A(new_n716), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n710), .A2(new_n990), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT44), .Z(new_n1003));
  NOR2_X1   g0803(.A1(new_n710), .A2(new_n990), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT45), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1001), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n711), .B1(new_n686), .B2(new_n697), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n708), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n715), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1003), .A2(new_n1005), .A3(new_n1001), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1007), .A2(new_n772), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1000), .B1(new_n1013), .B2(new_n772), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n776), .B(KEYINPUT114), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n999), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n837), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n238), .B2(new_n843), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n571), .A2(new_n718), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n779), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n807), .A2(new_n874), .B1(new_n787), .B2(new_n873), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n281), .B(new_n1022), .C1(G50), .C2(new_n871), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n820), .A2(G143), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n822), .A2(new_n217), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G159), .B2(new_n796), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n804), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1027), .A2(G58), .B1(new_n881), .B2(G77), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(G317), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n807), .A2(new_n825), .B1(new_n787), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n271), .B(new_n1031), .C1(G283), .C2(new_n871), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n796), .A2(G294), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n881), .A2(G97), .B1(new_n802), .B2(G107), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1027), .A2(G116), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT46), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT115), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1027), .A2(KEYINPUT115), .A3(KEYINPUT46), .A4(G116), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n819), .C2(new_n810), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1029), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT47), .Z(new_n1044));
  OAI221_X1 g0844(.A(new_n1021), .B1(new_n1044), .B2(new_n784), .C1(new_n981), .C2(new_n847), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1017), .A2(new_n1045), .ZN(G387));
  OAI22_X1  g0846(.A1(new_n838), .A2(new_n721), .B1(G107), .B2(new_n207), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n721), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n1048), .C1(G68), .C2(G77), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n344), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n718), .B(new_n271), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n235), .A2(G45), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1047), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n870), .A2(G50), .B1(new_n813), .B2(G150), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n271), .C1(new_n217), .C2(new_n806), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n797), .A2(new_n344), .B1(new_n788), .B2(new_n799), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n202), .A2(new_n804), .B1(new_n793), .B2(new_n543), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n369), .A2(new_n822), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n870), .A2(G317), .B1(new_n871), .B2(G303), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n797), .B2(new_n810), .C1(new_n819), .C2(new_n811), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1027), .A2(G294), .B1(new_n802), .B2(G283), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n271), .B1(new_n813), .B2(G326), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n501), .B2(new_n793), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1060), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n778), .B1(new_n1018), .B2(new_n1054), .C1(new_n1074), .C2(new_n784), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n711), .B2(new_n836), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT116), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n772), .A2(new_n1011), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n719), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n772), .A2(new_n1011), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(G393));
  INV_X1    g0882(.A(new_n1012), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1083), .A2(new_n1006), .A3(new_n1015), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n990), .A2(new_n836), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n837), .B1(new_n543), .B2(new_n207), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n246), .B2(new_n843), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(KEYINPUT117), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(KEYINPUT117), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n778), .A3(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n822), .A2(new_n202), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n797), .A2(new_n346), .B1(new_n793), .B2(new_n363), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G68), .C2(new_n1027), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n874), .A2(new_n799), .B1(new_n807), .B2(new_n788), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT51), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n871), .A2(new_n355), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n281), .B1(new_n813), .B2(G143), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n281), .B1(new_n787), .B2(new_n811), .C1(new_n492), .C2(new_n793), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G283), .B2(new_n1027), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT118), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n810), .A2(new_n807), .B1(new_n799), .B2(new_n1030), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n796), .A2(G303), .B1(G294), .B2(new_n871), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n501), .C2(new_n822), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1098), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT119), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1090), .B1(new_n1107), .B2(new_n833), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1084), .B1(new_n1085), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1079), .B1(new_n1083), .B2(new_n1006), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1013), .A2(new_n1110), .A3(new_n719), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(G390));
  NAND2_X1  g0912(.A1(new_n936), .A2(new_n953), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n957), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n697), .B1(new_n740), .B2(new_n746), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n860), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1113), .B1(new_n1117), .B2(new_n963), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n958), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n863), .B2(new_n864), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n963), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n953), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n950), .A2(new_n951), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n925), .A2(G330), .A3(new_n933), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n769), .A2(G330), .A3(new_n860), .A4(new_n963), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1129), .B(new_n1118), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1123), .A2(new_n834), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n778), .B1(new_n893), .B2(new_n355), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT54), .B(G143), .ZN(new_n1134));
  INV_X1    g0934(.A(G132), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n271), .B1(new_n806), .B2(new_n1134), .C1(new_n1135), .C2(new_n807), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n817), .B2(G125), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n804), .A2(new_n874), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n796), .A2(G137), .B1(new_n800), .B2(G128), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n881), .A2(G50), .B1(new_n802), .B2(G159), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1142), .A2(KEYINPUT122), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n816), .A2(new_n461), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n281), .B1(new_n806), .B2(new_n543), .C1(new_n501), .C2(new_n807), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n217), .A2(new_n793), .B1(new_n804), .B2(new_n363), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1091), .B1(G107), .B2(new_n796), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(new_n824), .C2(new_n799), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1142), .A2(KEYINPUT122), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1143), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1133), .B1(new_n1151), .B2(new_n833), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1131), .A2(new_n1016), .B1(new_n1132), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n457), .A2(G330), .A3(new_n925), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n966), .A2(new_n1154), .A3(new_n657), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT120), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n925), .A2(G330), .A3(new_n860), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1121), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1128), .A2(new_n1158), .A3(new_n1116), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n765), .A2(new_n768), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n767), .B1(new_n650), .B2(new_n924), .ZN(new_n1161));
  OAI211_X1 g0961(.A(G330), .B(new_n860), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1125), .B1(new_n1162), .B2(new_n1121), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1159), .B1(new_n1163), .B2(new_n1120), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT120), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n966), .A2(new_n1154), .A3(new_n1165), .A4(new_n657), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1156), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT121), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT121), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1156), .A2(new_n1164), .A3(new_n1169), .A4(new_n1166), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n719), .B1(new_n1131), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1118), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1128), .C1(new_n1174), .C2(new_n952), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1170), .B2(new_n1168), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1153), .B1(new_n1172), .B2(new_n1177), .ZN(G378));
  INV_X1    g0978(.A(KEYINPUT124), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1156), .A2(new_n1179), .A3(new_n1166), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n1156), .B2(new_n1166), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1184), .B2(new_n1176), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n935), .A2(G330), .A3(new_n937), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n349), .A2(new_n910), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n354), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n656), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n656), .A2(new_n1188), .A3(new_n1187), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1186), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1195), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1197), .A2(new_n935), .A3(G330), .A4(new_n937), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n965), .A2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n955), .A2(new_n1196), .A3(new_n964), .A4(new_n1198), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1182), .B1(new_n1131), .B2(new_n1171), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(KEYINPUT57), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n719), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1197), .A2(new_n835), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n271), .A2(new_n264), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n492), .B2(new_n807), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1025), .B(new_n1210), .C1(new_n817), .C2(G283), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n804), .A2(new_n202), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n799), .A2(new_n501), .B1(new_n793), .B2(new_n216), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G97), .C2(new_n796), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1211), .B(new_n1214), .C1(new_n369), .C2(new_n806), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT123), .Z(new_n1216));
  INV_X1    g1016(.A(KEYINPUT58), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(G33), .A2(G41), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1209), .A2(G50), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n800), .A2(G125), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n797), .B2(new_n1135), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G150), .B2(new_n802), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n870), .A2(G128), .B1(new_n871), .B2(G137), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n804), .C2(new_n1134), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  INV_X1    g1027(.A(G124), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1220), .B1(new_n787), .B2(new_n1228), .C1(new_n788), .C2(new_n793), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1226), .B2(KEYINPUT59), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1221), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1218), .A2(new_n1219), .A3(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n778), .B1(G50), .B2(new_n893), .C1(new_n1232), .C2(new_n784), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1208), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1202), .B2(new_n1016), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1207), .A2(new_n1235), .ZN(G375));
  NAND2_X1  g1036(.A1(new_n1121), .A2(new_n834), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n778), .B1(new_n893), .B2(G68), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n797), .A2(new_n1134), .B1(new_n804), .B2(new_n788), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G132), .B2(new_n800), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n817), .A2(G128), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n271), .B1(new_n806), .B2(new_n874), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G137), .B2(new_n870), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n881), .A2(G58), .B1(new_n802), .B2(G50), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1240), .A2(new_n1241), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n816), .A2(new_n825), .B1(new_n543), .B2(new_n804), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT125), .Z(new_n1247));
  OAI221_X1 g1047(.A(new_n281), .B1(new_n806), .B2(new_n492), .C1(new_n824), .C2(new_n807), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(new_n1059), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G294), .A2(new_n800), .B1(new_n881), .B2(G77), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n501), .C2(new_n797), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1245), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1238), .B1(new_n1252), .B2(new_n833), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1164), .A2(new_n1016), .B1(new_n1237), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1156), .A2(new_n1166), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1164), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1168), .A2(new_n1170), .A3(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1254), .B1(new_n1258), .B2(new_n1000), .ZN(G381));
  OR3_X1    g1059(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1260));
  NOR4_X1   g1060(.A1(G387), .A2(new_n1260), .A3(G390), .A4(G381), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1132), .A2(new_n1152), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1176), .B2(new_n1015), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n720), .B1(new_n1184), .B2(new_n1176), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1131), .A2(new_n1171), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1207), .A2(new_n1235), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1261), .A2(new_n1266), .A3(new_n1267), .ZN(G407));
  NAND2_X1  g1068(.A1(new_n694), .A2(G213), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1267), .A2(new_n1266), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G407), .A2(G213), .A3(new_n1271), .ZN(G409));
  XNOR2_X1  g1072(.A(G393), .B(new_n849), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1017), .A2(new_n1045), .A3(G390), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G390), .B1(new_n1017), .B2(new_n1045), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(G390), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1017), .A2(new_n1045), .A3(G390), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1273), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1235), .C1(new_n1203), .C2(new_n1206), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1201), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n964), .A2(new_n955), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1016), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1234), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1000), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1288), .B1(new_n1185), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT126), .B1(new_n1290), .B2(G378), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1289), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1235), .B1(new_n1204), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1266), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1283), .A2(new_n1291), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1258), .A2(KEYINPUT60), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1164), .B1(new_n1166), .B2(new_n1156), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n719), .B1(new_n1298), .B2(KEYINPUT60), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(G384), .A3(new_n1254), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1258), .B2(KEYINPUT60), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1254), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n896), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1296), .A2(new_n1269), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1296), .A2(new_n1309), .A3(new_n1269), .A4(new_n1306), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1290), .A2(G378), .A3(KEYINPUT126), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1294), .B1(new_n1266), .B2(new_n1293), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1270), .B1(new_n1315), .B2(new_n1283), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1270), .A2(G2897), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1306), .B2(KEYINPUT127), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT127), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1317), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1302), .A2(KEYINPUT127), .A3(new_n1305), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1318), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1312), .B1(new_n1316), .B2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1282), .B1(new_n1311), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1321), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1296), .A2(new_n1269), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT61), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  AND2_X1   g1131(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1316), .A2(KEYINPUT63), .A3(new_n1306), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1307), .A2(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1326), .A2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(G375), .A2(new_n1266), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1338), .A2(new_n1283), .A3(new_n1319), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1319), .B1(new_n1338), .B2(new_n1283), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1282), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1341), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1343), .A2(new_n1332), .A3(new_n1339), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1342), .A2(new_n1344), .ZN(G402));
endmodule


