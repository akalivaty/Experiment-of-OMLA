

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786;

  XNOR2_X1 U373 ( .A(n439), .B(G478), .ZN(n596) );
  XNOR2_X1 U374 ( .A(n516), .B(n515), .ZN(n542) );
  XNOR2_X1 U375 ( .A(n491), .B(G134), .ZN(n516) );
  XNOR2_X1 U376 ( .A(n573), .B(KEYINPUT111), .ZN(n422) );
  NOR2_X2 U377 ( .A1(n669), .A2(n757), .ZN(n670) );
  NOR2_X2 U378 ( .A1(n676), .A2(n757), .ZN(n677) );
  NOR2_X1 U379 ( .A1(G953), .A2(G237), .ZN(n402) );
  NOR2_X1 U380 ( .A1(n598), .A2(n596), .ZN(n508) );
  XNOR2_X1 U381 ( .A(n523), .B(n522), .ZN(n621) );
  AND2_X1 U382 ( .A1(n427), .A2(n704), .ZN(n424) );
  AND2_X1 U383 ( .A1(n420), .A2(n415), .ZN(n414) );
  XNOR2_X1 U384 ( .A(n641), .B(n640), .ZN(n392) );
  OR2_X1 U385 ( .A1(n784), .A2(n452), .ZN(n427) );
  NOR2_X1 U386 ( .A1(n735), .A2(n733), .ZN(n642) );
  AND2_X1 U387 ( .A1(n568), .A2(n616), .ZN(n403) );
  BUF_X1 U388 ( .A(n621), .Z(n555) );
  XNOR2_X1 U389 ( .A(n470), .B(n352), .ZN(n456) );
  XNOR2_X1 U390 ( .A(n506), .B(n437), .ZN(n598) );
  XNOR2_X1 U391 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U392 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U393 ( .A(n386), .B(n381), .ZN(n673) );
  XNOR2_X1 U394 ( .A(n383), .B(n382), .ZN(n381) );
  XNOR2_X1 U395 ( .A(n443), .B(n466), .ZN(n382) );
  XNOR2_X1 U396 ( .A(n464), .B(G146), .ZN(n495) );
  XNOR2_X2 U397 ( .A(KEYINPUT68), .B(G101), .ZN(n539) );
  XNOR2_X1 U398 ( .A(n759), .B(n519), .ZN(n386) );
  XNOR2_X1 U399 ( .A(n402), .B(n394), .ZN(n393) );
  INV_X1 U400 ( .A(KEYINPUT81), .ZN(n394) );
  AND2_X1 U401 ( .A1(n717), .A2(n411), .ZN(n592) );
  OR2_X1 U402 ( .A1(n349), .A2(n613), .ZN(n417) );
  NAND2_X1 U403 ( .A1(n419), .A2(KEYINPUT88), .ZN(n418) );
  INV_X1 U404 ( .A(n611), .ZN(n419) );
  XNOR2_X1 U405 ( .A(n580), .B(n579), .ZN(n429) );
  XNOR2_X1 U406 ( .A(n647), .B(n646), .ZN(n375) );
  AND2_X1 U407 ( .A1(n370), .A2(n653), .ZN(n369) );
  NAND2_X1 U408 ( .A1(n786), .A2(KEYINPUT90), .ZN(n370) );
  XNOR2_X1 U409 ( .A(n600), .B(n599), .ZN(n734) );
  INV_X1 U410 ( .A(G125), .ZN(n464) );
  XNOR2_X1 U411 ( .A(KEYINPUT15), .B(G902), .ZN(n657) );
  NAND2_X1 U412 ( .A1(n607), .A2(n608), .ZN(n610) );
  NAND2_X1 U413 ( .A1(n377), .A2(n588), .ZN(n608) );
  INV_X1 U414 ( .A(n617), .ZN(n632) );
  XNOR2_X1 U415 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n566) );
  BUF_X1 U416 ( .A(n551), .Z(n722) );
  NOR2_X1 U417 ( .A1(G902), .A2(n681), .ZN(n523) );
  NAND2_X1 U418 ( .A1(n393), .A2(G210), .ZN(n410) );
  XNOR2_X1 U419 ( .A(KEYINPUT4), .B(G131), .ZN(n515) );
  XNOR2_X1 U420 ( .A(n406), .B(n405), .ZN(n758) );
  INV_X1 U421 ( .A(G110), .ZN(n405) );
  XNOR2_X1 U422 ( .A(G107), .B(G104), .ZN(n406) );
  AND2_X1 U423 ( .A1(n393), .A2(G214), .ZN(n500) );
  XNOR2_X1 U424 ( .A(G131), .B(G140), .ZN(n501) );
  XNOR2_X1 U425 ( .A(n495), .B(n494), .ZN(n773) );
  INV_X1 U426 ( .A(KEYINPUT10), .ZN(n494) );
  XNOR2_X1 U427 ( .A(n758), .B(n387), .ZN(n519) );
  XNOR2_X1 U428 ( .A(n539), .B(KEYINPUT72), .ZN(n387) );
  NAND2_X1 U429 ( .A1(n592), .A2(n634), .ZN(n583) );
  BUF_X1 U430 ( .A(n456), .Z(n404) );
  XNOR2_X1 U431 ( .A(n507), .B(n438), .ZN(n437) );
  NOR2_X1 U432 ( .A1(G902), .A2(n665), .ZN(n506) );
  INV_X1 U433 ( .A(G475), .ZN(n438) );
  NAND2_X1 U434 ( .A1(n440), .A2(n544), .ZN(n439) );
  INV_X1 U435 ( .A(KEYINPUT64), .ZN(n442) );
  NAND2_X1 U436 ( .A1(n418), .A2(n416), .ZN(n415) );
  NAND2_X1 U437 ( .A1(n611), .A2(n417), .ZN(n416) );
  NAND2_X1 U438 ( .A1(n413), .A2(n351), .ZN(n412) );
  INV_X1 U439 ( .A(KEYINPUT46), .ZN(n452) );
  AND2_X1 U440 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U441 ( .A1(G234), .A2(G237), .ZN(n475) );
  NAND2_X1 U442 ( .A1(n530), .A2(G221), .ZN(n509) );
  XNOR2_X1 U443 ( .A(n376), .B(KEYINPUT20), .ZN(n530) );
  NAND2_X1 U444 ( .A1(n657), .A2(G234), .ZN(n376) );
  XNOR2_X1 U445 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n484) );
  NAND2_X1 U446 ( .A1(n374), .A2(n372), .ZN(n709) );
  NAND2_X1 U447 ( .A1(n373), .A2(KEYINPUT90), .ZN(n372) );
  NAND2_X1 U448 ( .A1(n615), .A2(n428), .ZN(n617) );
  AND2_X1 U449 ( .A1(n616), .A2(n614), .ZN(n428) );
  XNOR2_X1 U450 ( .A(n773), .B(n455), .ZN(n454) );
  XNOR2_X1 U451 ( .A(KEYINPUT99), .B(KEYINPUT97), .ZN(n455) );
  XNOR2_X1 U452 ( .A(G128), .B(KEYINPUT24), .ZN(n459) );
  XNOR2_X1 U453 ( .A(n461), .B(KEYINPUT98), .ZN(n460) );
  INV_X1 U454 ( .A(KEYINPUT23), .ZN(n461) );
  XNOR2_X1 U455 ( .A(G116), .B(G107), .ZN(n487) );
  XNOR2_X1 U456 ( .A(n385), .B(n384), .ZN(n383) );
  XNOR2_X1 U457 ( .A(n491), .B(KEYINPUT4), .ZN(n384) );
  XNOR2_X1 U458 ( .A(n463), .B(n495), .ZN(n385) );
  XOR2_X1 U459 ( .A(KEYINPUT17), .B(KEYINPUT86), .Z(n463) );
  INV_X1 U460 ( .A(n657), .ZN(n395) );
  INV_X1 U461 ( .A(n648), .ZN(n449) );
  NOR2_X1 U462 ( .A1(n576), .A2(KEYINPUT32), .ZN(n447) );
  XNOR2_X1 U463 ( .A(n474), .B(n473), .ZN(n623) );
  XNOR2_X1 U464 ( .A(n400), .B(n458), .ZN(n457) );
  INV_X1 U465 ( .A(KEYINPUT82), .ZN(n458) );
  NAND2_X1 U466 ( .A1(n403), .A2(n364), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n514), .B(n513), .ZN(n577) );
  XNOR2_X1 U468 ( .A(n410), .B(n536), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n536), .B(n465), .ZN(n759) );
  XNOR2_X1 U470 ( .A(KEYINPUT16), .B(G122), .ZN(n465) );
  XNOR2_X1 U471 ( .A(n504), .B(n505), .ZN(n665) );
  BUF_X1 U472 ( .A(n679), .Z(n753) );
  XNOR2_X1 U473 ( .A(n518), .B(n356), .ZN(n520) );
  NOR2_X1 U474 ( .A1(n749), .A2(G953), .ZN(n391) );
  NAND2_X1 U475 ( .A1(n462), .A2(n450), .ZN(n650) );
  NAND2_X1 U476 ( .A1(n445), .A2(n444), .ZN(n678) );
  AND2_X1 U477 ( .A1(n446), .A2(n448), .ZN(n445) );
  NAND2_X1 U478 ( .A1(n550), .A2(n447), .ZN(n444) );
  NAND2_X1 U479 ( .A1(n576), .A2(KEYINPUT32), .ZN(n448) );
  INV_X1 U480 ( .A(n726), .ZN(n441) );
  NAND2_X1 U481 ( .A1(n598), .A2(n597), .ZN(n698) );
  XNOR2_X1 U482 ( .A(n390), .B(n388), .ZN(G75) );
  XNOR2_X1 U483 ( .A(n389), .B(KEYINPUT53), .ZN(n388) );
  NAND2_X1 U484 ( .A1(n716), .A2(n391), .ZN(n390) );
  INV_X1 U485 ( .A(KEYINPUT120), .ZN(n389) );
  AND2_X1 U486 ( .A1(n598), .A2(n596), .ZN(n349) );
  XOR2_X1 U487 ( .A(n456), .B(KEYINPUT38), .Z(n350) );
  AND2_X1 U488 ( .A1(n611), .A2(KEYINPUT88), .ZN(n351) );
  XOR2_X1 U489 ( .A(n469), .B(n468), .Z(n352) );
  XOR2_X1 U490 ( .A(n545), .B(G472), .Z(n353) );
  XOR2_X1 U491 ( .A(G122), .B(G104), .Z(n354) );
  AND2_X1 U492 ( .A1(n651), .A2(n652), .ZN(n355) );
  XNOR2_X1 U493 ( .A(G146), .B(KEYINPUT84), .ZN(n356) );
  AND2_X1 U494 ( .A1(n621), .A2(KEYINPUT100), .ZN(n357) );
  AND2_X1 U495 ( .A1(n709), .A2(n706), .ZN(n358) );
  INV_X1 U496 ( .A(G210), .ZN(n535) );
  XOR2_X1 U497 ( .A(n502), .B(n501), .Z(n359) );
  XOR2_X1 U498 ( .A(n460), .B(n459), .Z(n360) );
  XOR2_X1 U499 ( .A(n482), .B(KEYINPUT0), .Z(n361) );
  XOR2_X1 U500 ( .A(n585), .B(KEYINPUT73), .Z(n362) );
  INV_X1 U501 ( .A(G953), .ZN(n763) );
  INV_X1 U502 ( .A(n577), .ZN(n550) );
  AND2_X2 U503 ( .A1(n367), .A2(n395), .ZN(n679) );
  NAND2_X1 U504 ( .A1(n363), .A2(n587), .ZN(n590) );
  INV_X1 U505 ( .A(n782), .ZN(n363) );
  XNOR2_X2 U506 ( .A(n430), .B(KEYINPUT35), .ZN(n782) );
  NAND2_X1 U507 ( .A1(n368), .A2(n396), .ZN(n367) );
  AND2_X1 U508 ( .A1(n364), .A2(n552), .ZN(n595) );
  NAND2_X1 U509 ( .A1(n558), .A2(n559), .ZN(n364) );
  NAND2_X1 U510 ( .A1(n366), .A2(n365), .ZN(n368) );
  NAND2_X1 U511 ( .A1(n398), .A2(n397), .ZN(n365) );
  NAND2_X1 U512 ( .A1(n399), .A2(n358), .ZN(n366) );
  AND2_X1 U513 ( .A1(n371), .A2(n369), .ZN(n374) );
  NAND2_X1 U514 ( .A1(n375), .A2(n355), .ZN(n371) );
  INV_X1 U515 ( .A(n375), .ZN(n373) );
  NAND2_X1 U516 ( .A1(n378), .A2(n586), .ZN(n377) );
  NAND2_X1 U517 ( .A1(n379), .A2(n589), .ZN(n378) );
  INV_X1 U518 ( .A(n429), .ZN(n379) );
  NAND2_X1 U519 ( .A1(n511), .A2(n380), .ZN(n514) );
  NAND2_X1 U520 ( .A1(n441), .A2(n380), .ZN(n594) );
  NAND2_X1 U521 ( .A1(n380), .A2(n595), .ZN(n686) );
  NAND2_X1 U522 ( .A1(n584), .A2(n380), .ZN(n432) );
  XNOR2_X2 U523 ( .A(n483), .B(n361), .ZN(n380) );
  XNOR2_X2 U524 ( .A(n409), .B(n408), .ZN(n536) );
  NAND2_X1 U525 ( .A1(n392), .A2(n426), .ZN(n425) );
  NOR2_X1 U526 ( .A1(n392), .A2(n452), .ZN(n451) );
  XNOR2_X1 U527 ( .A(n392), .B(G131), .ZN(G33) );
  INV_X1 U528 ( .A(n707), .ZN(n764) );
  NAND2_X1 U529 ( .A1(n707), .A2(KEYINPUT2), .ZN(n396) );
  INV_X1 U530 ( .A(n709), .ZN(n397) );
  INV_X1 U531 ( .A(n656), .ZN(n398) );
  INV_X1 U532 ( .A(n654), .ZN(n399) );
  NAND2_X1 U533 ( .A1(n639), .A2(n695), .ZN(n641) );
  XNOR2_X2 U534 ( .A(n571), .B(n570), .ZN(n639) );
  NOR2_X1 U535 ( .A1(n707), .A2(KEYINPUT80), .ZN(n654) );
  XNOR2_X1 U536 ( .A(n432), .B(n362), .ZN(n431) );
  NOR2_X2 U537 ( .A1(n615), .A2(n719), .ZN(n411) );
  NAND2_X1 U538 ( .A1(n555), .A2(n411), .ZN(n557) );
  XNOR2_X1 U539 ( .A(n401), .B(n453), .ZN(n754) );
  XNOR2_X1 U540 ( .A(n454), .B(n529), .ZN(n401) );
  NAND2_X1 U541 ( .A1(n525), .A2(G217), .ZN(n490) );
  XNOR2_X1 U542 ( .A(n486), .B(n485), .ZN(n525) );
  XNOR2_X1 U543 ( .A(n434), .B(n631), .ZN(n433) );
  XNOR2_X1 U544 ( .A(n407), .B(n541), .ZN(n543) );
  XNOR2_X2 U545 ( .A(KEYINPUT3), .B(G119), .ZN(n408) );
  XNOR2_X2 U546 ( .A(G116), .B(G113), .ZN(n409) );
  NAND2_X1 U547 ( .A1(n357), .A2(n411), .ZN(n559) );
  NAND2_X1 U548 ( .A1(n422), .A2(n349), .ZN(n612) );
  NAND2_X1 U549 ( .A1(n414), .A2(n412), .ZN(n435) );
  INV_X1 U550 ( .A(n422), .ZN(n413) );
  NAND2_X1 U551 ( .A1(n422), .A2(n421), .ZN(n420) );
  AND2_X1 U552 ( .A1(n349), .A2(n613), .ZN(n421) );
  NOR2_X1 U553 ( .A1(n423), .A2(n451), .ZN(n436) );
  NAND2_X1 U554 ( .A1(n425), .A2(n424), .ZN(n423) );
  AND2_X1 U555 ( .A1(n784), .A2(n452), .ZN(n426) );
  XNOR2_X2 U556 ( .A(n534), .B(n533), .ZN(n615) );
  NAND2_X1 U557 ( .A1(n591), .A2(n429), .ZN(n606) );
  NAND2_X1 U558 ( .A1(n431), .A2(n349), .ZN(n430) );
  NAND2_X1 U559 ( .A1(n436), .A2(n433), .ZN(n647) );
  NAND2_X1 U560 ( .A1(n435), .A2(n630), .ZN(n434) );
  INV_X1 U561 ( .A(n750), .ZN(n440) );
  INV_X1 U562 ( .A(n717), .ZN(n581) );
  XNOR2_X2 U563 ( .A(n621), .B(n524), .ZN(n717) );
  XNOR2_X1 U564 ( .A(n503), .B(n359), .ZN(n504) );
  XNOR2_X2 U565 ( .A(n583), .B(n582), .ZN(n744) );
  XNOR2_X2 U566 ( .A(n442), .B(G953), .ZN(n517) );
  NAND2_X1 U567 ( .A1(n517), .A2(G224), .ZN(n443) );
  NAND2_X1 U568 ( .A1(n577), .A2(KEYINPUT32), .ZN(n446) );
  NAND2_X1 U569 ( .A1(n678), .A2(n578), .ZN(n580) );
  NAND2_X1 U570 ( .A1(n456), .A2(n730), .ZN(n474) );
  NAND2_X1 U571 ( .A1(n449), .A2(n404), .ZN(n637) );
  INV_X1 U572 ( .A(n404), .ZN(n450) );
  NOR2_X1 U573 ( .A1(n754), .A2(G902), .ZN(n534) );
  XNOR2_X1 U574 ( .A(n360), .B(n528), .ZN(n453) );
  NAND2_X1 U575 ( .A1(n457), .A2(n404), .ZN(n573) );
  NAND2_X1 U576 ( .A1(n457), .A2(n350), .ZN(n571) );
  XOR2_X1 U577 ( .A(n649), .B(KEYINPUT43), .Z(n462) );
  XNOR2_X1 U578 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n524) );
  OR2_X1 U579 ( .A1(n517), .A2(G952), .ZN(n668) );
  XNOR2_X2 U580 ( .A(G143), .B(G128), .ZN(n491) );
  XOR2_X1 U581 ( .A(KEYINPUT85), .B(KEYINPUT18), .Z(n466) );
  NAND2_X1 U582 ( .A1(n673), .A2(n657), .ZN(n470) );
  NOR2_X1 U583 ( .A1(G237), .A2(G902), .ZN(n467) );
  XNOR2_X1 U584 ( .A(n467), .B(KEYINPUT78), .ZN(n471) );
  OR2_X1 U585 ( .A1(n471), .A2(n535), .ZN(n469) );
  INV_X1 U586 ( .A(KEYINPUT95), .ZN(n468) );
  INV_X1 U587 ( .A(G214), .ZN(n497) );
  OR2_X1 U588 ( .A1(n471), .A2(n497), .ZN(n730) );
  INV_X1 U589 ( .A(n730), .ZN(n565) );
  INV_X1 U590 ( .A(KEYINPUT83), .ZN(n472) );
  XNOR2_X1 U591 ( .A(n472), .B(KEYINPUT19), .ZN(n473) );
  XOR2_X1 U592 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n476) );
  XNOR2_X1 U593 ( .A(n476), .B(n475), .ZN(n479) );
  NAND2_X1 U594 ( .A1(G902), .A2(n479), .ZN(n560) );
  INV_X1 U595 ( .A(n560), .ZN(n477) );
  NOR2_X1 U596 ( .A1(G898), .A2(n763), .ZN(n761) );
  NAND2_X1 U597 ( .A1(n477), .A2(n761), .ZN(n478) );
  XNOR2_X1 U598 ( .A(n478), .B(KEYINPUT96), .ZN(n480) );
  NAND2_X1 U599 ( .A1(G952), .A2(n479), .ZN(n743) );
  OR2_X1 U600 ( .A1(n743), .A2(G953), .ZN(n563) );
  NAND2_X1 U601 ( .A1(n480), .A2(n563), .ZN(n481) );
  NAND2_X1 U602 ( .A1(n623), .A2(n481), .ZN(n483) );
  INV_X1 U603 ( .A(KEYINPUT67), .ZN(n482) );
  NAND2_X1 U604 ( .A1(G234), .A2(n517), .ZN(n486) );
  XNOR2_X1 U605 ( .A(n484), .B(KEYINPUT70), .ZN(n485) );
  XNOR2_X1 U606 ( .A(n487), .B(KEYINPUT9), .ZN(n488) );
  XOR2_X1 U607 ( .A(n488), .B(KEYINPUT7), .Z(n489) );
  XNOR2_X1 U608 ( .A(n490), .B(n489), .ZN(n493) );
  XOR2_X1 U609 ( .A(n516), .B(G122), .Z(n492) );
  XNOR2_X1 U610 ( .A(n493), .B(n492), .ZN(n750) );
  XNOR2_X1 U611 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n496) );
  XNOR2_X1 U612 ( .A(n496), .B(n773), .ZN(n505) );
  XNOR2_X1 U613 ( .A(G143), .B(G113), .ZN(n498) );
  XNOR2_X1 U614 ( .A(n354), .B(n498), .ZN(n499) );
  XNOR2_X1 U615 ( .A(n500), .B(n499), .ZN(n503) );
  XOR2_X1 U616 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n502) );
  INV_X1 U617 ( .A(KEYINPUT13), .ZN(n507) );
  XNOR2_X1 U618 ( .A(n508), .B(KEYINPUT105), .ZN(n733) );
  XOR2_X1 U619 ( .A(n509), .B(KEYINPUT21), .Z(n614) );
  INV_X1 U620 ( .A(n614), .ZN(n719) );
  NOR2_X1 U621 ( .A1(n733), .A2(n719), .ZN(n510) );
  XNOR2_X1 U622 ( .A(n510), .B(KEYINPUT106), .ZN(n511) );
  INV_X1 U623 ( .A(KEYINPUT75), .ZN(n512) );
  XNOR2_X1 U624 ( .A(n512), .B(KEYINPUT22), .ZN(n513) );
  XNOR2_X1 U625 ( .A(G137), .B(G140), .ZN(n526) );
  XNOR2_X1 U626 ( .A(n542), .B(n526), .ZN(n772) );
  NAND2_X1 U627 ( .A1(G227), .A2(n517), .ZN(n518) );
  XNOR2_X1 U628 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U629 ( .A(n772), .B(n521), .ZN(n681) );
  XNOR2_X1 U630 ( .A(KEYINPUT71), .B(G469), .ZN(n522) );
  NAND2_X1 U631 ( .A1(n525), .A2(G221), .ZN(n529) );
  XNOR2_X1 U632 ( .A(G119), .B(G110), .ZN(n527) );
  XNOR2_X1 U633 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U634 ( .A1(G217), .A2(n530), .ZN(n532) );
  INV_X1 U635 ( .A(KEYINPUT25), .ZN(n531) );
  XNOR2_X1 U636 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U637 ( .A1(n581), .A2(n615), .ZN(n548) );
  XNOR2_X1 U638 ( .A(G146), .B(G137), .ZN(n538) );
  XNOR2_X1 U639 ( .A(KEYINPUT79), .B(KEYINPUT5), .ZN(n537) );
  XNOR2_X1 U640 ( .A(n538), .B(n537), .ZN(n540) );
  XNOR2_X1 U641 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U642 ( .A(n542), .B(n543), .ZN(n658) );
  INV_X1 U643 ( .A(G902), .ZN(n544) );
  NAND2_X1 U644 ( .A1(n658), .A2(n544), .ZN(n546) );
  INV_X1 U645 ( .A(KEYINPUT74), .ZN(n545) );
  XNOR2_X2 U646 ( .A(n546), .B(n353), .ZN(n551) );
  XNOR2_X2 U647 ( .A(n551), .B(KEYINPUT107), .ZN(n618) );
  INV_X1 U648 ( .A(n618), .ZN(n547) );
  NOR2_X1 U649 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U650 ( .A1(n550), .A2(n549), .ZN(n578) );
  XNOR2_X1 U651 ( .A(n578), .B(G110), .ZN(G12) );
  NOR2_X1 U652 ( .A1(n615), .A2(n717), .ZN(n553) );
  INV_X1 U653 ( .A(n722), .ZN(n552) );
  XNOR2_X1 U654 ( .A(n552), .B(KEYINPUT6), .ZN(n634) );
  INV_X1 U655 ( .A(n634), .ZN(n574) );
  NAND2_X1 U656 ( .A1(n553), .A2(n574), .ZN(n554) );
  OR2_X1 U657 ( .A1(n577), .A2(n554), .ZN(n604) );
  XNOR2_X1 U658 ( .A(n604), .B(G101), .ZN(G3) );
  INV_X1 U659 ( .A(KEYINPUT100), .ZN(n556) );
  NAND2_X1 U660 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U661 ( .A1(n517), .A2(n560), .ZN(n561) );
  XOR2_X1 U662 ( .A(KEYINPUT108), .B(n561), .Z(n562) );
  OR2_X1 U663 ( .A1(n562), .A2(G900), .ZN(n564) );
  NAND2_X1 U664 ( .A1(n564), .A2(n563), .ZN(n616) );
  NOR2_X2 U665 ( .A1(n618), .A2(n565), .ZN(n567) );
  XNOR2_X1 U666 ( .A(n567), .B(n566), .ZN(n568) );
  INV_X1 U667 ( .A(KEYINPUT91), .ZN(n569) );
  XNOR2_X1 U668 ( .A(n569), .B(KEYINPUT39), .ZN(n570) );
  INV_X1 U669 ( .A(n598), .ZN(n572) );
  NAND2_X1 U670 ( .A1(n572), .A2(n596), .ZN(n701) );
  INV_X1 U671 ( .A(n701), .ZN(n690) );
  NAND2_X1 U672 ( .A1(n639), .A2(n690), .ZN(n653) );
  XNOR2_X1 U673 ( .A(n653), .B(G134), .ZN(G36) );
  XNOR2_X1 U674 ( .A(n612), .B(G143), .ZN(G45) );
  AND2_X1 U675 ( .A1(n615), .A2(n717), .ZN(n575) );
  NAND2_X1 U676 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U677 ( .A(KEYINPUT92), .ZN(n579) );
  INV_X1 U678 ( .A(KEYINPUT33), .ZN(n582) );
  INV_X1 U679 ( .A(n744), .ZN(n584) );
  XNOR2_X1 U680 ( .A(KEYINPUT34), .B(KEYINPUT87), .ZN(n585) );
  INV_X1 U681 ( .A(KEYINPUT44), .ZN(n587) );
  NOR2_X1 U682 ( .A1(n782), .A2(n587), .ZN(n586) );
  INV_X1 U683 ( .A(KEYINPUT65), .ZN(n589) );
  NAND2_X1 U684 ( .A1(n589), .A2(n587), .ZN(n588) );
  NAND2_X1 U685 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U686 ( .A1(n592), .A2(n722), .ZN(n726) );
  XNOR2_X1 U687 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n593) );
  XNOR2_X1 U688 ( .A(n594), .B(n593), .ZN(n700) );
  NAND2_X1 U689 ( .A1(n700), .A2(n686), .ZN(n602) );
  INV_X1 U690 ( .A(n596), .ZN(n597) );
  NAND2_X1 U691 ( .A1(n701), .A2(n698), .ZN(n600) );
  INV_X1 U692 ( .A(KEYINPUT104), .ZN(n599) );
  INV_X1 U693 ( .A(n734), .ZN(n601) );
  NAND2_X1 U694 ( .A1(n602), .A2(n601), .ZN(n603) );
  AND2_X1 U695 ( .A1(n604), .A2(n603), .ZN(n605) );
  INV_X1 U696 ( .A(KEYINPUT45), .ZN(n609) );
  XNOR2_X2 U697 ( .A(n610), .B(n609), .ZN(n707) );
  NAND2_X1 U698 ( .A1(n734), .A2(KEYINPUT47), .ZN(n611) );
  INV_X1 U699 ( .A(KEYINPUT88), .ZN(n613) );
  OR2_X1 U700 ( .A1(n734), .A2(KEYINPUT47), .ZN(n625) );
  OR2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n620) );
  INV_X1 U702 ( .A(KEYINPUT28), .ZN(n619) );
  XNOR2_X1 U703 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n622), .A2(n555), .ZN(n643) );
  INV_X1 U705 ( .A(n623), .ZN(n624) );
  NOR2_X1 U706 ( .A1(n643), .A2(n624), .ZN(n696) );
  NAND2_X1 U707 ( .A1(n625), .A2(n696), .ZN(n629) );
  INV_X1 U708 ( .A(n696), .ZN(n627) );
  INV_X1 U709 ( .A(KEYINPUT47), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n630) );
  INV_X1 U712 ( .A(KEYINPUT76), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n730), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n698), .A2(n633), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n648) );
  INV_X1 U716 ( .A(KEYINPUT36), .ZN(n636) );
  XNOR2_X1 U717 ( .A(n637), .B(n636), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n638), .A2(n717), .ZN(n704) );
  INV_X1 U719 ( .A(n698), .ZN(n695) );
  XNOR2_X1 U720 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n350), .A2(n730), .ZN(n735) );
  XNOR2_X1 U722 ( .A(n642), .B(KEYINPUT41), .ZN(n745) );
  NOR2_X1 U723 ( .A1(n745), .A2(n643), .ZN(n645) );
  XNOR2_X1 U724 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n644) );
  XNOR2_X1 U725 ( .A(n645), .B(n644), .ZN(n784) );
  INV_X1 U726 ( .A(KEYINPUT48), .ZN(n646) );
  NOR2_X1 U727 ( .A1(n717), .A2(n648), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n650), .B(KEYINPUT109), .ZN(n786) );
  INV_X1 U729 ( .A(n786), .ZN(n651) );
  INV_X1 U730 ( .A(KEYINPUT90), .ZN(n652) );
  INV_X1 U731 ( .A(KEYINPUT2), .ZN(n706) );
  NAND2_X1 U732 ( .A1(n706), .A2(KEYINPUT80), .ZN(n655) );
  NOR2_X1 U733 ( .A1(n707), .A2(n655), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n679), .A2(G472), .ZN(n661) );
  XNOR2_X1 U735 ( .A(KEYINPUT94), .B(KEYINPUT62), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n658), .B(n659), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U738 ( .A1(n662), .A2(n668), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U740 ( .A1(n679), .A2(G475), .ZN(n667) );
  XNOR2_X1 U741 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n664) );
  XNOR2_X1 U742 ( .A(n667), .B(n666), .ZN(n669) );
  INV_X1 U743 ( .A(n668), .ZN(n757) );
  XNOR2_X1 U744 ( .A(n670), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U745 ( .A1(n679), .A2(G210), .ZN(n675) );
  XOR2_X1 U746 ( .A(KEYINPUT93), .B(KEYINPUT54), .Z(n671) );
  XNOR2_X1 U747 ( .A(n671), .B(KEYINPUT55), .ZN(n672) );
  XNOR2_X1 U748 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U749 ( .A(n677), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U750 ( .A(n678), .B(G119), .ZN(G21) );
  NAND2_X1 U751 ( .A1(n753), .A2(G469), .ZN(n683) );
  XOR2_X1 U752 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n680) );
  XNOR2_X1 U753 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U755 ( .A1(n684), .A2(n757), .ZN(G54) );
  NOR2_X1 U756 ( .A1(n686), .A2(n698), .ZN(n685) );
  XOR2_X1 U757 ( .A(G104), .B(n685), .Z(G6) );
  NOR2_X1 U758 ( .A1(n686), .A2(n701), .ZN(n688) );
  XNOR2_X1 U759 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U761 ( .A(G107), .B(n689), .ZN(G9) );
  XOR2_X1 U762 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n692) );
  NAND2_X1 U763 ( .A1(n690), .A2(n696), .ZN(n691) );
  XNOR2_X1 U764 ( .A(n692), .B(n691), .ZN(n694) );
  XOR2_X1 U765 ( .A(G128), .B(KEYINPUT114), .Z(n693) );
  XNOR2_X1 U766 ( .A(n694), .B(n693), .ZN(G30) );
  NAND2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U768 ( .A(n697), .B(G146), .ZN(G48) );
  NOR2_X1 U769 ( .A1(n698), .A2(n700), .ZN(n699) );
  XOR2_X1 U770 ( .A(G113), .B(n699), .Z(G15) );
  NOR2_X1 U771 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U772 ( .A(G116), .B(n702), .Z(G18) );
  XOR2_X1 U773 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n703) );
  XNOR2_X1 U774 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U775 ( .A(G125), .B(n705), .ZN(G27) );
  NAND2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U777 ( .A(KEYINPUT89), .B(n708), .Z(n715) );
  BUF_X1 U778 ( .A(n709), .Z(n710) );
  NAND2_X1 U779 ( .A1(n764), .A2(KEYINPUT2), .ZN(n711) );
  NAND2_X1 U780 ( .A1(n397), .A2(n711), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n710), .A2(KEYINPUT2), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U784 ( .A1(n717), .A2(n411), .ZN(n718) );
  XOR2_X1 U785 ( .A(KEYINPUT50), .B(n718), .Z(n725) );
  XOR2_X1 U786 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n721) );
  NAND2_X1 U787 ( .A1(n615), .A2(n719), .ZN(n720) );
  XNOR2_X1 U788 ( .A(n721), .B(n720), .ZN(n723) );
  NOR2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n727) );
  AND2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U792 ( .A(KEYINPUT51), .B(n728), .Z(n729) );
  NOR2_X1 U793 ( .A1(n745), .A2(n729), .ZN(n740) );
  NOR2_X1 U794 ( .A1(n350), .A2(n730), .ZN(n731) );
  XNOR2_X1 U795 ( .A(n731), .B(KEYINPUT118), .ZN(n732) );
  NOR2_X1 U796 ( .A1(n733), .A2(n732), .ZN(n737) );
  NOR2_X1 U797 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U798 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U799 ( .A1(n738), .A2(n744), .ZN(n739) );
  NOR2_X1 U800 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U801 ( .A(n741), .B(KEYINPUT52), .ZN(n742) );
  NOR2_X1 U802 ( .A1(n743), .A2(n742), .ZN(n747) );
  NOR2_X1 U803 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U804 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U805 ( .A(n748), .B(KEYINPUT119), .ZN(n749) );
  NAND2_X1 U806 ( .A1(n753), .A2(G478), .ZN(n751) );
  XNOR2_X1 U807 ( .A(n750), .B(n751), .ZN(n752) );
  NOR2_X1 U808 ( .A1(n757), .A2(n752), .ZN(G63) );
  NAND2_X1 U809 ( .A1(n753), .A2(G217), .ZN(n755) );
  XNOR2_X1 U810 ( .A(n755), .B(n754), .ZN(n756) );
  NOR2_X1 U811 ( .A1(n757), .A2(n756), .ZN(G66) );
  XNOR2_X1 U812 ( .A(n758), .B(G101), .ZN(n760) );
  XOR2_X1 U813 ( .A(n760), .B(n759), .Z(n762) );
  NOR2_X1 U814 ( .A1(n762), .A2(n761), .ZN(n771) );
  NAND2_X1 U815 ( .A1(n764), .A2(n763), .ZN(n768) );
  NAND2_X1 U816 ( .A1(G953), .A2(G224), .ZN(n765) );
  XNOR2_X1 U817 ( .A(KEYINPUT61), .B(n765), .ZN(n766) );
  NAND2_X1 U818 ( .A1(n766), .A2(G898), .ZN(n767) );
  NAND2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U820 ( .A(n769), .B(KEYINPUT122), .ZN(n770) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(G69) );
  XOR2_X1 U822 ( .A(n772), .B(n773), .Z(n777) );
  XNOR2_X1 U823 ( .A(G227), .B(n777), .ZN(n774) );
  NAND2_X1 U824 ( .A1(n774), .A2(G900), .ZN(n775) );
  XNOR2_X1 U825 ( .A(n775), .B(KEYINPUT124), .ZN(n776) );
  NAND2_X1 U826 ( .A1(n776), .A2(G953), .ZN(n781) );
  XOR2_X1 U827 ( .A(KEYINPUT123), .B(n777), .Z(n778) );
  XNOR2_X1 U828 ( .A(n710), .B(n778), .ZN(n779) );
  NAND2_X1 U829 ( .A1(n779), .A2(n517), .ZN(n780) );
  NAND2_X1 U830 ( .A1(n781), .A2(n780), .ZN(G72) );
  XNOR2_X1 U831 ( .A(n782), .B(G122), .ZN(n783) );
  XNOR2_X1 U832 ( .A(n783), .B(KEYINPUT125), .ZN(G24) );
  XNOR2_X1 U833 ( .A(G137), .B(n784), .ZN(n785) );
  XNOR2_X1 U834 ( .A(n785), .B(KEYINPUT126), .ZN(G39) );
  XOR2_X1 U835 ( .A(G140), .B(n786), .Z(G42) );
endmodule

