//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1207,
    new_n1208, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  NOR2_X1   g0016(.A1(G58), .A2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n219), .A2(G50), .A3(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  INV_X1    g0029(.A(G238), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n228), .B1(new_n202), .B2(new_n229), .C1(new_n203), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n210), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n213), .B1(new_n216), .B2(new_n221), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n229), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(new_n203), .A2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n208), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n251), .B1(new_n252), .B2(new_n223), .C1(new_n254), .C2(new_n201), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n214), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT11), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n208), .A3(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n207), .A2(KEYINPUT12), .A3(G13), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n260), .B1(KEYINPUT12), .B2(new_n262), .C1(new_n251), .C2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n259), .A2(KEYINPUT11), .ZN(new_n265));
  INV_X1    g0065(.A(new_n257), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G1), .B2(new_n208), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n203), .B1(new_n267), .B2(KEYINPUT12), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n264), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n214), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n229), .A2(G1698), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n277), .B(new_n278), .C1(G226), .C2(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G97), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n272), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n270), .B2(new_n271), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  AOI21_X1  g0085(.A(G1), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n286), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n272), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n287), .B1(new_n289), .B2(new_n230), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT13), .B1(new_n281), .B2(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n291), .A2(KEYINPUT73), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n281), .A2(new_n290), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT13), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(KEYINPUT73), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n292), .A2(G190), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n269), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n291), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(G200), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  AOI211_X1 g0103(.A(KEYINPUT72), .B(new_n303), .C1(new_n295), .C2(new_n291), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n299), .A2(new_n306), .A3(KEYINPUT74), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT74), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n298), .B2(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G238), .A2(G1698), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n277), .B(new_n311), .C1(new_n229), .C2(G1698), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(G107), .C2(new_n277), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n287), .C1(new_n224), .C2(new_n289), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G200), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n315), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n319), .A2(new_n252), .B1(new_n208), .B2(new_n223), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(new_n254), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n257), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT69), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n262), .A2(new_n223), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n324), .B(new_n325), .C1(new_n223), .C2(new_n267), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n315), .A2(G179), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n315), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n326), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT70), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n301), .A2(G169), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n292), .A2(G179), .A3(new_n295), .A4(new_n296), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n269), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G222), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G223), .A2(G1698), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n277), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(new_n313), .C1(G77), .C2(new_n277), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n272), .A2(G226), .A3(new_n288), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n287), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(G179), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n329), .B2(new_n347), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n253), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT67), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n321), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n202), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n350), .B1(new_n354), .B2(new_n252), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n257), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n201), .B1(new_n207), .B2(G20), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT68), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n262), .A2(new_n257), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n358), .A2(new_n359), .B1(new_n201), .B2(new_n262), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n349), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AND4_X1   g0163(.A1(new_n310), .A2(new_n333), .A3(new_n340), .A4(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(G223), .A2(G1698), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n277), .B(new_n365), .C1(G226), .C2(new_n341), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G33), .A2(G87), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n272), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n287), .B1(new_n289), .B2(new_n229), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n368), .A2(new_n369), .A3(new_n317), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n368), .A2(new_n369), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n370), .B1(G200), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  AND2_X1   g0173(.A1(KEYINPUT3), .A2(G33), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT3), .A2(G33), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NOR4_X1   g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(G20), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n277), .B2(G20), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n203), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n202), .A2(new_n203), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(new_n217), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G20), .B1(G159), .B2(new_n253), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n373), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT75), .B1(new_n374), .B2(new_n375), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT75), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n275), .A2(new_n387), .A3(new_n276), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n388), .A3(new_n208), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n377), .B1(new_n389), .B2(new_n376), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT16), .B(new_n383), .C1(new_n390), .C2(new_n203), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n385), .A2(new_n391), .A3(new_n257), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n354), .A2(new_n267), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n262), .B2(new_n354), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n372), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT76), .B1(new_n395), .B2(KEYINPUT17), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n395), .A2(KEYINPUT76), .A3(KEYINPUT17), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n372), .A2(new_n392), .A3(new_n398), .A4(new_n394), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT77), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n399), .A2(new_n400), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n396), .A2(new_n397), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n392), .A2(new_n394), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n371), .A2(G169), .ZN(new_n405));
  INV_X1    g0205(.A(G179), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n371), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g0208(.A(new_n408), .B(KEYINPUT18), .Z(new_n409));
  NAND2_X1  g0209(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n361), .A2(KEYINPUT9), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT9), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n356), .A2(new_n413), .A3(new_n360), .ZN(new_n414));
  INV_X1    g0214(.A(new_n347), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n412), .A2(new_n414), .B1(G190), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n347), .A2(G200), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT10), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n412), .A2(new_n414), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(G190), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(KEYINPUT71), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n416), .B(new_n417), .C1(KEYINPUT71), .C2(KEYINPUT10), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n364), .A2(new_n411), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n207), .A2(G45), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT79), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G41), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n428), .B1(new_n430), .B2(KEYINPUT5), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT5), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n429), .B2(G41), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n283), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n313), .B1(new_n431), .B2(new_n433), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G257), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .A4(new_n341), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G283), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n277), .A2(G250), .A3(G1698), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n277), .A2(G244), .A3(new_n341), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT4), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT78), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT78), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n441), .A2(new_n445), .A3(new_n442), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n440), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n434), .B(new_n436), .C1(new_n447), .C2(new_n272), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G200), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n207), .A2(G33), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n359), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G97), .ZN(new_n453));
  INV_X1    g0253(.A(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n262), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(KEYINPUT6), .A3(G97), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n454), .A2(new_n457), .ZN(new_n459));
  NOR2_X1   g0259(.A1(G97), .A2(G107), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n458), .B1(new_n461), .B2(KEYINPUT6), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n462), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n378), .A2(new_n379), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(new_n457), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n456), .B1(new_n465), .B2(new_n257), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n449), .B(new_n466), .C1(new_n317), .C2(new_n448), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n436), .A2(new_n434), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n444), .A2(new_n446), .ZN(new_n469));
  INV_X1    g0269(.A(new_n440), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n313), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n406), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n448), .A2(new_n329), .ZN(new_n474));
  INV_X1    g0274(.A(new_n466), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n467), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n208), .B(G87), .C1(new_n374), .C2(new_n375), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT85), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT85), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n277), .A2(new_n480), .A3(new_n208), .A4(G87), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT22), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(KEYINPUT85), .A3(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n208), .A2(KEYINPUT23), .A3(G107), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT86), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n485), .A2(new_n486), .B1(KEYINPUT23), .B2(G107), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n274), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n457), .A3(G20), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n208), .B1(new_n491), .B2(KEYINPUT86), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n484), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT24), .B1(new_n482), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT22), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n492), .A2(new_n487), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n484), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n266), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n262), .A2(new_n457), .ZN(new_n500));
  XOR2_X1   g0300(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n501));
  XNOR2_X1  g0301(.A(new_n500), .B(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n457), .B2(new_n451), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(G250), .B(new_n341), .C1(new_n374), .C2(new_n375), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G294), .ZN(new_n506));
  AND2_X1   g0306(.A1(G257), .A2(G1698), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n374), .B2(new_n375), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n435), .A2(G264), .B1(new_n509), .B2(new_n313), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n317), .A3(new_n434), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT88), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n434), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(G200), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n511), .A2(new_n512), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n504), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(G169), .B1(new_n510), .B2(new_n434), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n509), .A2(new_n313), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n285), .A2(G1), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n284), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n433), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G264), .A3(new_n272), .ZN(new_n524));
  AND4_X1   g0324(.A1(new_n406), .A2(new_n520), .A3(new_n434), .A4(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n499), .B2(new_n503), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n477), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n341), .A2(G257), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G264), .A2(G1698), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n275), .A2(new_n276), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G303), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n374), .A2(new_n375), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT82), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT82), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n275), .A2(G303), .A3(new_n276), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n530), .A2(new_n531), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n374), .A2(new_n375), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n540), .A3(new_n313), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n523), .A2(G270), .A3(new_n272), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n434), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT83), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n541), .A2(new_n543), .A3(KEYINPUT83), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n303), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n262), .A2(new_n489), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n359), .A2(G116), .A3(new_n450), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n256), .A2(new_n214), .B1(G20), .B2(new_n489), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n438), .B(new_n208), .C1(G33), .C2(new_n454), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT20), .B1(new_n552), .B2(new_n553), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n550), .B(new_n551), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n317), .B1(new_n546), .B2(new_n547), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n549), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n551), .A2(new_n550), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n554), .B(new_n555), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n329), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n546), .A2(new_n563), .A3(new_n547), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n541), .A2(new_n543), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT84), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(G179), .A4(new_n558), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n558), .A2(new_n543), .A3(new_n541), .A4(G179), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT84), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n546), .A2(new_n563), .A3(KEYINPUT21), .A4(new_n547), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n560), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n319), .ZN(new_n576));
  INV_X1    g0376(.A(new_n262), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n452), .A2(G87), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n277), .A2(new_n208), .A3(G68), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT80), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n280), .B2(new_n208), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n225), .A2(new_n454), .A3(new_n457), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n585), .A2(new_n586), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n579), .B(new_n580), .C1(new_n589), .C2(new_n266), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n224), .A2(G1698), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(G238), .B2(G1698), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n592), .A2(new_n539), .B1(new_n274), .B2(new_n489), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n313), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n521), .A2(new_n282), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n428), .A2(new_n226), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n272), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G190), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n303), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n266), .B1(new_n583), .B2(new_n588), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n451), .A2(new_n319), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n602), .A2(new_n578), .A3(new_n603), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n604), .A2(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n598), .A2(new_n406), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G169), .B2(new_n598), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n604), .B2(KEYINPUT81), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n529), .A2(new_n575), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n427), .A2(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n409), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n299), .A2(new_n306), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n340), .B1(new_n614), .B2(new_n331), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n615), .B2(new_n403), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n423), .A2(KEYINPUT90), .A3(new_n424), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT90), .B1(new_n423), .B2(new_n424), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n362), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n604), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n597), .A2(KEYINPUT89), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n597), .A2(KEYINPUT89), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n594), .A3(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n329), .A2(new_n625), .B1(new_n598), .B2(new_n406), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n566), .A2(new_n527), .A3(new_n572), .A4(new_n573), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n518), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n625), .A2(G200), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n599), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n590), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n467), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n629), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n609), .A2(KEYINPUT26), .A3(new_n630), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n628), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n621), .B1(new_n427), .B2(new_n639), .ZN(G369));
  NAND3_X1  g0440(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n558), .A2(new_n646), .ZN(new_n647));
  MUX2_X1   g0447(.A(new_n575), .B(new_n574), .S(new_n647), .Z(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n528), .ZN(new_n651));
  INV_X1    g0451(.A(new_n646), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n504), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n527), .B2(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n574), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n651), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n655), .B(new_n657), .C1(new_n527), .C2(new_n646), .ZN(G399));
  INV_X1    g0458(.A(new_n211), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n586), .A2(G116), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G1), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n221), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT28), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n631), .A2(new_n518), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n636), .B1(new_n666), .B2(new_n476), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n638), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n646), .B1(new_n668), .B2(new_n627), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n630), .A2(new_n635), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n628), .B1(new_n672), .B2(KEYINPUT26), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n609), .A2(new_n629), .A3(new_n630), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n635), .A2(new_n627), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n477), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n673), .B(new_n674), .C1(new_n666), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n652), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT29), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n544), .A2(new_n406), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n598), .A2(new_n510), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n472), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT30), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n472), .A2(new_n681), .A3(KEYINPUT30), .A4(new_n680), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n448), .A2(new_n406), .A3(new_n514), .A4(new_n625), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n684), .B(new_n685), .C1(new_n548), .C2(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n687), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT31), .B1(new_n687), .B2(new_n646), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n529), .A2(new_n575), .A3(new_n609), .A4(new_n652), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n671), .A2(new_n679), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n665), .B1(new_n694), .B2(G1), .ZN(G364));
  NOR2_X1   g0495(.A1(new_n261), .A2(G20), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G45), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n661), .A2(G1), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n650), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(G330), .B2(new_n648), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n214), .B1(G20), .B2(new_n329), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n208), .A2(new_n406), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT92), .Z(new_n704));
  NOR2_X1   g0504(.A1(G190), .A2(G200), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G311), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n208), .A2(G179), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(new_n317), .A3(G200), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G283), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n706), .A2(new_n707), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n317), .A2(G200), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n406), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G294), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n317), .A2(new_n303), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n703), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n277), .B(new_n721), .C1(G326), .C2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n703), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n726), .A2(new_n303), .A3(G190), .ZN(new_n727));
  XNOR2_X1  g0527(.A(KEYINPUT33), .B(G317), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n708), .A2(new_n705), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n727), .A2(new_n728), .B1(G329), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(new_n708), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n725), .B(new_n731), .C1(new_n533), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n704), .A2(new_n716), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n715), .B(new_n733), .C1(G322), .C2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n713), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G107), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(new_n202), .B2(new_n734), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n539), .B1(new_n727), .B2(G68), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n732), .A2(new_n225), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(G50), .B2(new_n724), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n740), .B(new_n742), .C1(new_n706), .C2(new_n223), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n719), .A2(new_n454), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n730), .A2(G159), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT32), .ZN(new_n746));
  NOR4_X1   g0546(.A1(new_n739), .A2(new_n743), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n702), .B1(new_n736), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n659), .A2(new_n539), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n749), .A2(G355), .B1(new_n489), .B2(new_n659), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n386), .A2(new_n388), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n659), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G45), .B2(new_n221), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n246), .A2(new_n285), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT91), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n702), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n755), .A2(KEYINPUT91), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n756), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n748), .A2(new_n762), .A3(new_n699), .ZN(new_n763));
  INV_X1    g0563(.A(new_n759), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n648), .B2(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n701), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(G396));
  XNOR2_X1  g0567(.A(new_n331), .B(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n327), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n638), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n666), .A2(new_n476), .ZN(new_n772));
  INV_X1    g0572(.A(new_n636), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(new_n774), .B2(new_n629), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n652), .B(new_n770), .C1(new_n775), .C2(new_n628), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n326), .A2(new_n646), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n769), .A2(new_n777), .B1(new_n331), .B2(new_n652), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n776), .B1(new_n669), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n699), .B1(new_n779), .B2(new_n693), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n693), .B2(new_n779), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n702), .A2(new_n757), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n698), .B1(new_n223), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n702), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n706), .A2(new_n489), .B1(new_n533), .B2(new_n723), .ZN(new_n785));
  INV_X1    g0585(.A(new_n727), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n785), .B1(new_n790), .B2(G283), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n734), .A2(new_n720), .B1(new_n713), .B2(new_n225), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n539), .B1(new_n729), .B2(new_n707), .C1(new_n732), .C2(new_n457), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n793), .A2(new_n744), .A3(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n727), .A2(G150), .B1(new_n724), .B2(G137), .ZN(new_n796));
  INV_X1    g0596(.A(G143), .ZN(new_n797));
  INV_X1    g0597(.A(G159), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n734), .B2(new_n797), .C1(new_n798), .C2(new_n706), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT34), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n713), .A2(new_n203), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n732), .A2(new_n201), .B1(new_n729), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n751), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(G58), .C2(new_n718), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n792), .A2(new_n795), .B1(new_n800), .B2(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n783), .B1(new_n784), .B2(new_n808), .C1(new_n778), .C2(new_n758), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n781), .A2(new_n809), .ZN(G384));
  NOR2_X1   g0610(.A1(new_n696), .A2(new_n207), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n612), .A2(new_n644), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT38), .ZN(new_n813));
  INV_X1    g0613(.A(new_n644), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n391), .A2(new_n257), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n383), .B1(new_n390), .B2(new_n203), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT16), .B1(new_n816), .B2(KEYINPUT100), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT100), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n818), .B(new_n383), .C1(new_n390), .C2(new_n203), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n815), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n394), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n814), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n407), .B1(new_n820), .B2(new_n821), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(new_n823), .A3(new_n395), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n824), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT101), .B1(new_n824), .B2(KEYINPUT37), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n404), .A2(new_n814), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n408), .A2(new_n827), .A3(new_n395), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(KEYINPUT37), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n825), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n822), .B1(new_n403), .B2(new_n409), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n813), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n826), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n824), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n828), .A2(KEYINPUT37), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n822), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n410), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n838), .A3(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n269), .A2(new_n652), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n340), .A2(new_n613), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n338), .B1(new_n307), .B2(new_n309), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(new_n842), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT98), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n639), .A2(new_n646), .A3(new_n769), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n768), .A2(new_n646), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n849), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n776), .A2(KEYINPUT98), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n846), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT99), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n840), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n847), .B(new_n849), .C1(new_n669), .C2(new_n770), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT98), .B1(new_n776), .B2(new_n851), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(KEYINPUT99), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n812), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n340), .A2(new_n646), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n828), .A2(KEYINPUT37), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n835), .A2(KEYINPUT103), .A3(new_n864), .ZN(new_n865));
  OR3_X1    g0665(.A1(new_n828), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n827), .B1(new_n403), .B2(new_n409), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n813), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT39), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n839), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n832), .B2(new_n839), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(KEYINPUT102), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n874), .B(new_n870), .C1(new_n832), .C2(new_n839), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n863), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n830), .A2(new_n813), .A3(new_n831), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n836), .B2(new_n838), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT39), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n874), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(KEYINPUT102), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT104), .A4(new_n871), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n862), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n860), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT105), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n427), .B1(new_n671), .B2(new_n679), .ZN(new_n886));
  INV_X1    g0686(.A(new_n621), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n885), .B(new_n888), .Z(new_n889));
  AND3_X1   g0689(.A1(new_n692), .A2(new_n845), .A3(new_n778), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n840), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n692), .A2(new_n845), .A3(new_n778), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n839), .A2(new_n869), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n891), .A2(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n364), .A2(new_n692), .A3(new_n411), .A4(new_n426), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(G330), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n898), .B2(new_n897), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n811), .B1(new_n889), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n889), .B2(new_n902), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n906));
  NOR4_X1   g0706(.A1(new_n905), .A2(new_n906), .A3(new_n216), .A4(new_n489), .ZN(new_n907));
  XOR2_X1   g0707(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n908));
  XOR2_X1   g0708(.A(new_n907), .B(new_n908), .Z(new_n909));
  OR3_X1    g0709(.A1(new_n221), .A2(new_n223), .A3(new_n381), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n201), .A2(G68), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(G1), .A3(new_n261), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n904), .A2(new_n909), .A3(new_n913), .ZN(G367));
  INV_X1    g0714(.A(new_n752), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n760), .B1(new_n211), .B2(new_n319), .C1(new_n915), .C2(new_n241), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n699), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT108), .Z(new_n918));
  NAND2_X1  g0718(.A1(new_n590), .A2(new_n646), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n635), .A2(new_n627), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n627), .B2(new_n919), .ZN(new_n921));
  INV_X1    g0721(.A(new_n706), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n790), .A2(G159), .B1(G50), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n737), .A2(G77), .ZN(new_n924));
  INV_X1    g0724(.A(G150), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n734), .ZN(new_n926));
  INV_X1    g0726(.A(new_n732), .ZN(new_n927));
  AOI22_X1  g0727(.A1(G143), .A2(new_n724), .B1(new_n927), .B2(G58), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n539), .B1(new_n730), .B2(G137), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n928), .B(new_n929), .C1(new_n203), .C2(new_n719), .ZN(new_n930));
  AOI22_X1  g0730(.A1(G283), .A2(new_n922), .B1(new_n735), .B2(G303), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n720), .B2(new_n789), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n737), .A2(G97), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n732), .A2(new_n489), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n934), .A2(KEYINPUT46), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n934), .A2(KEYINPUT46), .B1(new_n718), .B2(G107), .ZN(new_n936));
  INV_X1    g0736(.A(G317), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n723), .A2(new_n707), .B1(new_n729), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(new_n751), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n933), .A2(new_n935), .A3(new_n936), .A4(new_n939), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n926), .A2(new_n930), .B1(new_n932), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT47), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n702), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n941), .A2(new_n942), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n918), .B1(new_n764), .B2(new_n921), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n697), .A2(G1), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n476), .A2(new_n652), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT106), .Z(new_n949));
  AOI21_X1  g0749(.A(new_n477), .B1(new_n475), .B2(new_n646), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n657), .B1(new_n527), .B2(new_n646), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT44), .Z(new_n954));
  NOR2_X1   g0754(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT45), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT107), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n655), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n657), .B1(new_n654), .B2(new_n656), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n650), .B(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n694), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n694), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n660), .B(KEYINPUT41), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n947), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n951), .A2(new_n657), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT42), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n476), .B1(new_n951), .B2(new_n527), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n652), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n966), .A2(new_n968), .B1(KEYINPUT43), .B2(new_n921), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n655), .A2(new_n951), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n946), .B1(new_n964), .B2(new_n973), .ZN(G387));
  NAND2_X1  g0774(.A1(new_n960), .A2(new_n947), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n654), .A2(new_n764), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n732), .A2(new_n223), .B1(new_n729), .B2(new_n925), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n751), .B1(new_n719), .B2(new_n319), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(G159), .C2(new_n724), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n922), .A2(G68), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n786), .A2(new_n354), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n735), .B2(G50), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n979), .A2(new_n933), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n751), .B1(G326), .B2(new_n730), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n719), .A2(new_n714), .B1(new_n732), .B2(new_n720), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G303), .A2(new_n922), .B1(new_n735), .B2(G317), .ZN(new_n986));
  INV_X1    g0786(.A(G322), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n986), .B1(new_n707), .B2(new_n789), .C1(new_n987), .C2(new_n723), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT48), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n989), .B2(new_n988), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT49), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n984), .B1(new_n489), .B2(new_n713), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n983), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT110), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n784), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n996), .B2(new_n995), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n238), .A2(G45), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n662), .B(new_n285), .C1(new_n203), .C2(new_n223), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT109), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n321), .A2(G50), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT50), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(KEYINPUT109), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n999), .B(new_n752), .C1(new_n1001), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n749), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(G107), .B2(new_n211), .C1(new_n662), .C2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n698), .B1(new_n1008), .B2(new_n760), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n998), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n694), .A2(new_n960), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n660), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n694), .A2(new_n960), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n975), .B1(new_n976), .B2(new_n1010), .C1(new_n1012), .C2(new_n1013), .ZN(G393));
  NAND2_X1  g0814(.A1(new_n954), .A2(new_n956), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(new_n655), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n1011), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n961), .A2(new_n1017), .A3(new_n660), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n951), .A2(new_n759), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n790), .A2(G303), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n539), .B1(new_n729), .B2(new_n987), .C1(new_n732), .C2(new_n714), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G116), .B2(new_n718), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n922), .A2(G294), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n738), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n734), .A2(new_n707), .B1(new_n937), .B2(new_n723), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT52), .Z(new_n1026));
  OAI22_X1  g0826(.A1(new_n734), .A2(new_n798), .B1(new_n925), .B2(new_n723), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT51), .Z(new_n1028));
  INV_X1    g0828(.A(new_n321), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n922), .A2(new_n1029), .B1(new_n737), .B2(G87), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n719), .A2(new_n223), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n732), .A2(new_n203), .B1(new_n729), .B2(new_n797), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1031), .A2(new_n805), .A3(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1030), .B(new_n1033), .C1(new_n201), .C2(new_n789), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n1024), .A2(new_n1026), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n702), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n760), .B1(new_n454), .B2(new_n211), .C1(new_n915), .C2(new_n249), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1019), .A2(new_n699), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n947), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1018), .B(new_n1038), .C1(new_n1039), .C2(new_n1016), .ZN(G390));
  OAI21_X1  g0840(.A(new_n888), .B1(new_n427), .B2(new_n693), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n890), .A2(G330), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n692), .A2(G330), .A3(new_n778), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1043), .B1(new_n845), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n850), .A2(new_n852), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n851), .B1(new_n678), .B2(new_n769), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1042), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n858), .A2(new_n862), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n876), .A2(new_n1051), .A3(new_n882), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1048), .A2(new_n845), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n861), .B(KEYINPUT111), .Z(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n895), .A3(new_n1054), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1052), .A2(new_n1055), .A3(new_n1043), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1043), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1050), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1043), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1052), .A2(new_n1055), .A3(new_n1043), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(new_n1041), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1058), .A2(new_n1065), .A3(new_n660), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT112), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT112), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1058), .A2(new_n1065), .A3(new_n1068), .A4(new_n660), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1061), .A2(new_n947), .A3(new_n1062), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n698), .B1(new_n354), .B2(new_n782), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n790), .A2(G107), .B1(G116), .B2(new_n735), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n723), .A2(new_n714), .B1(new_n729), .B2(new_n720), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n1031), .A2(new_n1073), .A3(new_n741), .A4(new_n277), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n801), .B1(new_n922), .B2(G97), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n790), .A2(G137), .B1(G132), .B2(new_n735), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n927), .A2(G150), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT53), .ZN(new_n1079));
  INV_X1    g0879(.A(G128), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n719), .A2(new_n798), .B1(new_n723), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT54), .B(G143), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1077), .B(new_n1082), .C1(new_n706), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n539), .B1(new_n730), .B2(G125), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n713), .B2(new_n201), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT113), .Z(new_n1087));
  OAI21_X1  g0887(.A(new_n1076), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n702), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n876), .A2(new_n882), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1071), .B1(new_n1089), .B2(new_n1091), .C1(new_n1092), .C2(new_n758), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1070), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT115), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1070), .A2(KEYINPUT115), .A3(new_n1093), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1067), .A2(new_n1069), .A3(new_n1096), .A4(new_n1097), .ZN(G378));
  INV_X1    g0898(.A(KEYINPUT57), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1092), .A2(new_n861), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n890), .A2(new_n895), .A3(KEYINPUT40), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n893), .B1(new_n839), .B2(new_n832), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(G330), .C1(new_n1102), .C2(KEYINPUT40), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n361), .A2(new_n814), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT118), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n620), .B2(new_n363), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1107), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n618), .A2(new_n619), .A3(new_n362), .A4(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1105), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n619), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n423), .A2(KEYINPUT90), .A3(new_n424), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1112), .A2(new_n363), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1109), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n620), .A2(new_n363), .A3(new_n1107), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n1116), .A3(new_n1104), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1103), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1111), .A2(KEYINPUT119), .A3(new_n1117), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT119), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1119), .B1(new_n1103), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n840), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n858), .B2(KEYINPUT99), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(KEYINPUT99), .B2(new_n858), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1100), .A2(new_n1123), .A3(new_n1126), .A4(new_n812), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n896), .A2(G330), .B1(new_n1117), .B2(new_n1111), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1103), .A2(new_n1122), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n860), .B2(new_n883), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1099), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1056), .A2(new_n1057), .A3(new_n1050), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n1041), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n660), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT120), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1065), .A2(new_n1042), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n661), .B1(new_n1138), .B2(new_n1132), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT120), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1065), .A2(new_n1042), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(KEYINPUT57), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1144), .A2(new_n1039), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n757), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n732), .A2(new_n223), .B1(new_n729), .B2(new_n714), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n786), .A2(new_n454), .B1(new_n723), .B2(new_n489), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(G68), .C2(new_n718), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G107), .A2(new_n735), .B1(new_n922), .B2(new_n576), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n751), .A2(G41), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n737), .A2(G58), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT58), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1151), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G50), .B1(new_n274), .B2(new_n284), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1153), .A2(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT116), .Z(new_n1158));
  OAI22_X1  g0958(.A1(new_n786), .A2(new_n803), .B1(new_n732), .B2(new_n1083), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n735), .B2(G128), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G125), .A2(new_n724), .B1(new_n718), .B2(G150), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT117), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n922), .A2(G137), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1160), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n730), .C2(G124), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(new_n798), .C2(new_n713), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1167), .A2(new_n1168), .B1(new_n1154), .B2(new_n1153), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n702), .B1(new_n1158), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n698), .B1(new_n201), .B2(new_n782), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1146), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1145), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1143), .A2(new_n1173), .ZN(G375));
  NAND2_X1  g0974(.A1(new_n1063), .A2(new_n1041), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1050), .A2(new_n1175), .A3(new_n963), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n947), .B(KEYINPUT121), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT122), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n782), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n699), .B1(G68), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n846), .A2(new_n757), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT123), .Z(new_n1185));
  AOI22_X1  g0985(.A1(G294), .A2(new_n724), .B1(new_n927), .B2(G97), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n277), .B1(new_n730), .B2(G303), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n319), .C2(new_n719), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n790), .A2(G116), .B1(G283), .B2(new_n735), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1189), .B(new_n924), .C1(new_n457), .C2(new_n706), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1083), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n790), .A2(new_n1191), .B1(G137), .B2(new_n735), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n1152), .C1(new_n925), .C2(new_n706), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n805), .B1(G50), .B2(new_n718), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G132), .A2(new_n724), .B1(new_n927), .B2(G159), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n1080), .C2(new_n729), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1188), .A2(new_n1190), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1183), .B(new_n1185), .C1(new_n702), .C2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1176), .A2(new_n1181), .A3(new_n1199), .ZN(G381));
  INV_X1    g1000(.A(G375), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1096), .A2(new_n1066), .A3(new_n1097), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(G387), .A2(G390), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(G407));
  NAND2_X1  g1006(.A1(new_n645), .A2(G213), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1201), .A2(new_n1203), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(G407), .A2(G213), .A3(new_n1209), .ZN(G409));
  INV_X1    g1010(.A(KEYINPUT60), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1050), .B(new_n660), .C1(new_n1175), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1211), .B2(new_n1175), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1199), .A2(new_n1181), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1215), .A2(G384), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(G384), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT125), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1139), .A2(KEYINPUT120), .B1(KEYINPUT57), .B2(new_n1141), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1136), .B(new_n661), .C1(new_n1138), .C2(new_n1132), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G378), .B(new_n1173), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT124), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT124), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1143), .A2(new_n1225), .A3(G378), .A4(new_n1173), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1178), .B1(new_n1138), .B2(new_n963), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(new_n1144), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1202), .B1(new_n1229), .B2(new_n1172), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1220), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  AOI211_X1 g1032(.A(KEYINPUT125), .B(new_n1230), .C1(new_n1224), .C2(new_n1226), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1207), .B(new_n1219), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT62), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1208), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1218), .A2(new_n1235), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1236), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1208), .A2(G2897), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1218), .B(new_n1242), .Z(new_n1243));
  NOR2_X1   g1043(.A1(new_n1237), .A2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(KEYINPUT61), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1241), .A2(KEYINPUT126), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT126), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1239), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1245), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  XOR2_X1   g1050(.A(G387), .B(G390), .Z(new_n1251));
  XNOR2_X1  g1051(.A(G393), .B(new_n766), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT127), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1246), .A2(new_n1250), .A3(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1237), .A2(KEYINPUT63), .A3(new_n1219), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1255), .A2(KEYINPUT61), .A3(new_n1256), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(new_n1208), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1234), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1262), .B1(new_n1264), .B2(new_n1243), .C1(KEYINPUT63), .C2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1259), .A2(new_n1266), .ZN(G405));
  OAI21_X1  g1067(.A(new_n1227), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(new_n1219), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1258), .B(new_n1269), .ZN(G402));
endmodule


