//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT68), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT70), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n460), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n475), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  INV_X1    g057(.A(new_n476), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n463), .A2(new_n469), .A3(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n475), .A2(KEYINPUT71), .A3(G126), .A4(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n494), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT74), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(KEYINPUT73), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n510), .B(G543), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT72), .B1(new_n513), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(new_n508), .A3(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n509), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G62), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n506), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT6), .B(G651), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(G50), .A2(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G166));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT6), .B(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT75), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(G543), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n509), .A2(new_n515), .A3(new_n519), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n524), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n536), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n535), .A2(G52), .B1(G90), .B2(new_n538), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n506), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n535), .A2(G43), .B1(G81), .B2(new_n538), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n537), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n553), .A2(KEYINPUT78), .A3(G651), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(G651), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n550), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND4_X1  g139(.A1(new_n530), .A2(G53), .A3(G543), .A4(new_n532), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT79), .Z(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n537), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(new_n538), .B2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n546), .A2(new_n548), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  NAND2_X1  g150(.A1(new_n513), .A2(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n508), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(new_n510), .B1(new_n516), .B2(new_n518), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n579), .A2(G87), .A3(new_n509), .A4(new_n531), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n530), .A2(G49), .A3(G543), .A4(new_n532), .ZN(new_n581));
  AOI21_X1  g156(.A(G74), .B1(new_n579), .B2(new_n509), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n506), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT80), .ZN(new_n584));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n515), .A2(new_n519), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n578), .A2(new_n510), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n589), .A2(new_n590), .A3(new_n580), .A4(new_n581), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n584), .A2(new_n591), .ZN(G288));
  NAND4_X1  g167(.A1(new_n509), .A2(G86), .A3(new_n515), .A4(new_n519), .ZN(new_n593));
  NAND2_X1  g168(.A1(G48), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n524), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n509), .A2(G61), .A3(new_n515), .A4(new_n519), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT81), .Z(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n596), .A2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n535), .A2(G47), .B1(G85), .B2(new_n538), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(new_n506), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n538), .A2(G92), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT10), .Z(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n537), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n535), .A2(G54), .B1(G651), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n607), .B1(new_n615), .B2(G868), .ZN(G321));
  XOR2_X1   g191(.A(G321), .B(KEYINPUT82), .Z(G284));
  MUX2_X1   g192(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g193(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n615), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g200(.A1(new_n463), .A2(new_n469), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n473), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT83), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n481), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n460), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n483), .A2(KEYINPUT84), .A3(G135), .ZN(new_n636));
  AOI21_X1  g211(.A(KEYINPUT84), .B1(new_n483), .B2(G135), .ZN(new_n637));
  OAI221_X1 g212(.A(new_n633), .B1(new_n634), .B2(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n629), .B2(new_n630), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n632), .A2(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n645), .B(new_n651), .Z(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  AND3_X1   g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(KEYINPUT17), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n661), .B1(new_n662), .B2(new_n659), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n662), .A2(new_n659), .A3(new_n658), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n672), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  MUX2_X1   g263(.A(G6), .B(G305), .S(G16), .Z(new_n689));
  XOR2_X1   g264(.A(KEYINPUT32), .B(G1981), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT87), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n692), .A2(new_n693), .ZN(new_n700));
  MUX2_X1   g275(.A(G23), .B(new_n583), .S(G16), .Z(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT33), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n694), .A2(new_n699), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n706));
  MUX2_X1   g281(.A(G24), .B(G290), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G1986), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n481), .A2(G119), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n483), .A2(G131), .ZN(new_n710));
  OR2_X1    g285(.A1(G95), .A2(G2105), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n711), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT86), .Z(new_n714));
  MUX2_X1   g289(.A(G25), .B(new_n714), .S(G29), .Z(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n705), .A2(new_n706), .A3(new_n708), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT89), .B(KEYINPUT36), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(G168), .A2(G16), .ZN(new_n721));
  NOR2_X1   g296(.A1(G16), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(KEYINPUT94), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(KEYINPUT94), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1966), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n695), .A2(G4), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n615), .B2(new_n695), .ZN(new_n727));
  INV_X1    g302(.A(G1348), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n695), .A2(G20), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT23), .Z(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G299), .B2(G16), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1956), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n725), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n695), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n559), .B2(new_n695), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1341), .ZN(new_n737));
  NOR2_X1   g312(.A1(G171), .A2(new_n695), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G5), .B2(new_n695), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  NOR2_X1   g315(.A1(G29), .A2(G33), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT25), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G139), .B2(new_n483), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n626), .A2(G127), .ZN(new_n745));
  NAND2_X1  g320(.A1(G115), .A2(G2104), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n460), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n748), .B2(new_n747), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n741), .B1(new_n750), .B2(G29), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n739), .A2(new_n740), .B1(G2072), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n740), .B2(new_n739), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G32), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n473), .ZN(new_n756));
  INV_X1    g331(.A(G129), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n480), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT93), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT92), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n758), .B1(new_n761), .B2(KEYINPUT26), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(KEYINPUT26), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n755), .B1(new_n765), .B2(new_n754), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n754), .A2(G35), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT95), .Z(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n754), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT29), .B(G2090), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT30), .B(G28), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n754), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n638), .B2(new_n754), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n754), .A2(G26), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT28), .ZN(new_n780));
  INV_X1    g355(.A(G128), .ZN(new_n781));
  INV_X1    g356(.A(G140), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n781), .A2(new_n480), .B1(new_n476), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G104), .A2(G2105), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT90), .ZN(new_n785));
  INV_X1    g360(.A(G116), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n465), .B1(new_n786), .B2(G2105), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n783), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n780), .B1(new_n788), .B2(new_n754), .ZN(new_n789));
  INV_X1    g364(.A(G2067), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n771), .A2(new_n772), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n778), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT24), .ZN(new_n794));
  INV_X1    g369(.A(G34), .ZN(new_n795));
  AOI21_X1  g370(.A(G29), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G160), .B2(new_n754), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2084), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n754), .A2(G27), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n754), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2078), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n793), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n768), .B(new_n803), .C1(G2072), .C2(new_n751), .ZN(new_n804));
  OR4_X1    g379(.A1(new_n734), .A2(new_n737), .A3(new_n753), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n720), .A2(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  NAND2_X1  g382(.A1(new_n535), .A2(G55), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n538), .A2(G93), .ZN(new_n809));
  NAND2_X1  g384(.A1(G80), .A2(G543), .ZN(new_n810));
  INV_X1    g385(.A(G67), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n537), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n812), .A2(G651), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n808), .B(new_n809), .C1(KEYINPUT96), .C2(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n813), .A2(KEYINPUT96), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT98), .B(G860), .Z(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT37), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n615), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n816), .A2(new_n559), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n558), .B1(new_n814), .B2(new_n815), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n821), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT99), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n826), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n825), .A2(KEYINPUT97), .A3(new_n826), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n831), .A2(new_n817), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n819), .B1(new_n828), .B2(new_n833), .ZN(G145));
  AOI21_X1  g409(.A(new_n502), .B1(new_n497), .B2(new_n498), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT100), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT100), .B1(new_n491), .B2(new_n493), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n788), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n764), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n750), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n481), .A2(G130), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n483), .A2(G142), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n460), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n628), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n713), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT101), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n850), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n841), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G160), .B(new_n487), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(new_n638), .Z(new_n858));
  AOI21_X1  g433(.A(G37), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n852), .B(new_n860), .C1(new_n842), .C2(new_n850), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT102), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n859), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n863), .A2(KEYINPUT40), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT40), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(G395));
  XNOR2_X1  g443(.A(new_n824), .B(new_n622), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n615), .B(G299), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT41), .ZN(new_n872));
  XNOR2_X1  g447(.A(G299), .B(new_n614), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(new_n873), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT42), .ZN(new_n880));
  XNOR2_X1  g455(.A(G290), .B(G305), .ZN(new_n881));
  XNOR2_X1  g456(.A(G166), .B(new_n583), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n884), .A3(new_n878), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n880), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n880), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(G868), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(G868), .B2(new_n816), .ZN(G295));
  OAI21_X1  g464(.A(new_n888), .B1(G868), .B2(new_n816), .ZN(G331));
  XOR2_X1   g465(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n891));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  XNOR2_X1  g467(.A(G171), .B(G168), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n824), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n824), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n875), .A3(new_n872), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n824), .A2(new_n893), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(new_n873), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(KEYINPUT104), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n824), .A2(new_n893), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n883), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n897), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n883), .B(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n897), .A2(new_n903), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n892), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n900), .A2(new_n894), .A3(new_n902), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n875), .A3(new_n872), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n899), .A2(new_n895), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n907), .A2(new_n918), .A3(KEYINPUT43), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n891), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n908), .A2(new_n892), .A3(new_n913), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n907), .B2(new_n918), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT44), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(G397));
  INV_X1    g499(.A(G1384), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT106), .B1(new_n838), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(KEYINPUT45), .ZN(new_n927));
  INV_X1    g502(.A(G40), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n472), .A2(new_n928), .A3(new_n478), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n838), .A2(KEYINPUT106), .A3(new_n925), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OR3_X1    g506(.A1(new_n931), .A2(G1986), .A3(G290), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(G1986), .A3(G290), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n935), .B(KEYINPUT107), .Z(new_n936));
  XNOR2_X1  g511(.A(new_n788), .B(new_n790), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n764), .B2(G1996), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n931), .A2(G1996), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT108), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n941), .B2(new_n765), .ZN(new_n942));
  INV_X1    g517(.A(new_n716), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n713), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n933), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n936), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT109), .Z(new_n948));
  INV_X1    g523(.A(KEYINPUT49), .ZN(new_n949));
  INV_X1    g524(.A(G1981), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n596), .B2(new_n601), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n506), .B1(new_n597), .B2(new_n599), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n595), .A2(new_n952), .A3(G1981), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n838), .A2(new_n929), .A3(new_n925), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n955), .A2(G8), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n596), .A2(new_n601), .A3(new_n950), .ZN(new_n957));
  OAI21_X1  g532(.A(G1981), .B1(new_n595), .B2(new_n952), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT49), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n589), .A2(G1976), .A3(new_n580), .A4(new_n581), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n955), .A2(new_n961), .A3(G8), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n963));
  INV_X1    g538(.A(G1976), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n584), .A2(new_n964), .A3(new_n591), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n955), .A2(new_n961), .A3(G8), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT52), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n960), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(G8), .B1(new_n523), .B2(new_n527), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT55), .B(G8), .C1(new_n523), .C2(new_n527), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n838), .A2(KEYINPUT45), .A3(new_n925), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n504), .A2(new_n925), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n835), .B2(new_n494), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT110), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n975), .A2(new_n979), .A3(new_n929), .A4(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n982), .A2(new_n698), .ZN(new_n983));
  INV_X1    g558(.A(new_n478), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n470), .A2(new_n471), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(G40), .B(new_n984), .C1(new_n986), .C2(new_n460), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(KEYINPUT50), .B2(new_n976), .ZN(new_n988));
  INV_X1    g563(.A(G2090), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n838), .A2(new_n990), .A3(new_n925), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(G8), .B(new_n974), .C1(new_n983), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n499), .A2(new_n503), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT100), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n494), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT100), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT50), .B1(new_n1000), .B2(G1384), .ZN(new_n1001));
  AOI211_X1 g576(.A(KEYINPUT50), .B(G1384), .C1(new_n835), .C2(new_n494), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(new_n987), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n990), .B1(new_n838), .B2(new_n925), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n504), .A2(new_n990), .A3(new_n925), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n929), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT111), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1005), .A2(new_n1009), .A3(new_n989), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n982), .A2(new_n698), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n995), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n969), .B(new_n994), .C1(new_n974), .C2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT58), .B(G1341), .Z(new_n1014));
  NAND2_X1  g589(.A1(new_n955), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT120), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n982), .A2(G1996), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n559), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT59), .ZN(new_n1019));
  INV_X1    g594(.A(G1956), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT116), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT57), .B1(new_n571), .B2(new_n566), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n566), .A2(KEYINPUT79), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n566), .A2(KEYINPUT79), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1026), .A2(KEYINPUT57), .A3(new_n571), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT56), .B(G2072), .Z(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT118), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n982), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1022), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT61), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1022), .A2(new_n1030), .A3(KEYINPUT61), .A4(new_n1033), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n955), .A2(G2067), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n988), .A2(new_n991), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(new_n728), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(new_n614), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n614), .A2(KEYINPUT60), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1042), .A2(KEYINPUT60), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1019), .A2(new_n1038), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1030), .B1(new_n1022), .B2(new_n1033), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1041), .A2(new_n614), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT119), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1046), .B1(new_n1048), .B2(new_n1034), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1013), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n982), .B2(G2078), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1040), .A2(new_n740), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT45), .B1(new_n838), .B2(new_n925), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n925), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n929), .ZN(new_n1058));
  OR4_X1    g633(.A1(new_n1052), .A2(new_n1056), .A3(new_n1058), .A4(G2078), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1051), .B1(new_n1060), .B2(G301), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n927), .A2(new_n930), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n986), .A2(KEYINPUT122), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n986), .A2(KEYINPUT122), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(G2105), .A3(new_n1064), .ZN(new_n1065));
  NOR4_X1   g640(.A1(new_n478), .A2(new_n1052), .A3(new_n928), .A4(G2078), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1062), .A2(new_n975), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1055), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT123), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G171), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1068), .A2(KEYINPUT123), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1061), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1060), .A2(G171), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n1051), .C1(G171), .C2(new_n1068), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n1076));
  INV_X1    g651(.A(G1966), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G2084), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n988), .A2(new_n1081), .A3(new_n991), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT112), .B(new_n1077), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(G168), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1084), .A2(G8), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1083), .A2(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1080), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G286), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1076), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1084), .A2(G8), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(KEYINPUT51), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT121), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(G168), .B1(new_n1086), .B2(new_n1080), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT51), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1094), .B(new_n1095), .C1(KEYINPUT51), .C2(new_n1090), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1050), .A2(new_n1075), .A3(new_n1092), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1087), .A2(G8), .A3(G168), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1013), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n960), .A2(new_n966), .A3(new_n968), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n995), .B1(new_n1011), .B2(new_n992), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n974), .ZN(new_n1104));
  INV_X1    g679(.A(new_n974), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n995), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n995), .B(G286), .C1(new_n1086), .C2(new_n1080), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1104), .A2(new_n1107), .A3(KEYINPUT113), .A4(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1100), .A2(new_n1101), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(G8), .B1(new_n983), .B2(new_n993), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n974), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1112), .B2(new_n1111), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(KEYINPUT63), .A3(new_n1104), .A4(new_n1108), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G288), .A2(G1976), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n954), .A2(new_n959), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n953), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n956), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n994), .A2(new_n1102), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT115), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1124), .B(new_n1121), .C1(new_n1110), .C2(new_n1115), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1097), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1073), .A2(new_n1013), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1092), .A2(KEYINPUT124), .A3(new_n1096), .A4(KEYINPUT62), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n948), .B1(new_n1126), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n714), .A2(new_n943), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n942), .A2(new_n1136), .B1(new_n790), .B2(new_n788), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n932), .B(KEYINPUT48), .Z(new_n1138));
  OAI22_X1  g713(.A1(new_n1137), .A2(new_n931), .B1(new_n946), .B2(new_n1138), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n941), .A2(KEYINPUT46), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n933), .B1(new_n764), .B2(new_n937), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT125), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n941), .A2(KEYINPUT46), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1144), .A2(KEYINPUT126), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(KEYINPUT126), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT47), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT47), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n1149), .A3(new_n1146), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1139), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1135), .A2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g727(.A1(new_n914), .A2(new_n919), .ZN(new_n1154));
  INV_X1    g728(.A(new_n458), .ZN(new_n1155));
  NOR2_X1   g729(.A1(G227), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g730(.A(new_n1156), .B(KEYINPUT127), .ZN(new_n1157));
  NOR3_X1   g731(.A1(G229), .A2(G401), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g732(.A(new_n865), .ZN(new_n1159));
  AOI21_X1  g733(.A(new_n864), .B1(new_n859), .B2(new_n861), .ZN(new_n1160));
  OAI21_X1  g734(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g735(.A1(new_n1154), .A2(new_n1161), .ZN(G308));
  OAI221_X1 g736(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .C1(new_n914), .C2(new_n919), .ZN(G225));
endmodule


