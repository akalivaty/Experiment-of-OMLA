//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G107), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n191), .B1(KEYINPUT74), .B2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(KEYINPUT75), .A3(G104), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n195), .B2(new_n196), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n194), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G101), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n202), .B(new_n194), .C1(new_n198), .C2(new_n199), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT64), .B1(new_n205), .B2(G146), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n212), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n211), .A2(new_n214), .B1(new_n212), .B2(new_n216), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n200), .A2(new_n223), .A3(G101), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n204), .A2(new_n220), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT11), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G137), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT65), .A2(G134), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT65), .A2(G134), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G137), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT11), .A3(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(G137), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(G131), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n229), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(KEYINPUT11), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT65), .A2(G134), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n232), .A4(new_n233), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n235), .A2(KEYINPUT66), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(G131), .C1(new_n230), .C2(new_n234), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n216), .A2(new_n246), .A3(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n205), .A2(G146), .ZN(new_n248));
  OAI21_X1  g062(.A(G128), .B1(new_n248), .B2(new_n246), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n250), .B2(new_n216), .ZN(new_n251));
  OAI21_X1  g065(.A(G101), .B1(new_n193), .B2(new_n191), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n203), .A3(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n203), .A2(new_n252), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n211), .A2(new_n249), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n247), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(KEYINPUT10), .A3(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n225), .A2(new_n245), .A3(new_n255), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT77), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n203), .A2(new_n252), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n257), .A2(new_n247), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT10), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n224), .A2(new_n220), .A3(new_n222), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n204), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n245), .A4(new_n255), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n245), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n258), .B1(new_n203), .B2(new_n252), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT78), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n253), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n262), .A2(new_n273), .A3(new_n263), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT12), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT12), .B(new_n271), .C1(new_n274), .C2(new_n275), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n270), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(G110), .B(G140), .ZN(new_n282));
  INV_X1    g096(.A(G227), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G953), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n282), .B(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n261), .B2(new_n269), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n225), .A2(new_n255), .A3(new_n259), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT79), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n225), .A2(KEYINPUT79), .A3(new_n255), .A4(new_n259), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n271), .A3(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n281), .A2(new_n285), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G469), .B1(new_n292), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT80), .B(G469), .Z(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n285), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n270), .A2(new_n280), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n270), .B2(new_n291), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n294), .B(new_n296), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n189), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G478), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(KEYINPUT15), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G217), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n187), .A2(new_n305), .A3(G953), .ZN(new_n306));
  INV_X1    g120(.A(G122), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT87), .B1(new_n307), .B2(G116), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n309));
  INV_X1    g123(.A(G116), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G122), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(G116), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G107), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n190), .A3(new_n313), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT88), .ZN(new_n317));
  INV_X1    g131(.A(G128), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G143), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n205), .A2(KEYINPUT88), .A3(G128), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(G143), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n228), .A2(new_n229), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n315), .A2(new_n316), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT13), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n205), .A2(KEYINPUT88), .A3(G128), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT88), .B1(new_n205), .B2(G128), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n319), .A2(KEYINPUT13), .A3(new_n320), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n322), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n332), .A2(new_n333), .A3(G134), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n332), .B2(G134), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n326), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT90), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n338), .B(new_n326), .C1(new_n334), .C2(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n190), .B1(new_n313), .B2(KEYINPUT14), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n314), .B(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n324), .A2(new_n325), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n325), .B1(new_n321), .B2(new_n322), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(KEYINPUT91), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT91), .ZN(new_n347));
  INV_X1    g161(.A(new_n325), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n323), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n349), .B2(new_n344), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n342), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n306), .B1(new_n340), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n306), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n351), .B(new_n354), .C1(new_n337), .C2(new_n339), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n294), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT92), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n332), .A2(G134), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT89), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n332), .A2(new_n333), .A3(G134), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n338), .B1(new_n361), .B2(new_n326), .ZN(new_n362));
  INV_X1    g176(.A(new_n339), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n352), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n354), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n340), .A2(new_n352), .A3(new_n306), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT92), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(new_n294), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n304), .B1(new_n357), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G475), .A2(G902), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G113), .B(G122), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(new_n192), .ZN(new_n374));
  NOR2_X1   g188(.A1(G237), .A2(G953), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(G143), .A3(G214), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(G143), .B1(new_n375), .B2(G214), .ZN(new_n378));
  OAI211_X1 g192(.A(KEYINPUT18), .B(G131), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n378), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT18), .A2(G131), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G125), .ZN(new_n384));
  INV_X1    g198(.A(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G140), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G146), .ZN(new_n388));
  XNOR2_X1  g202(.A(G125), .B(G140), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(new_n208), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n379), .B(new_n382), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n385), .A2(KEYINPUT16), .A3(G140), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT16), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n208), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n389), .B2(KEYINPUT16), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G146), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT71), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n395), .A2(KEYINPUT71), .A3(new_n208), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT17), .ZN(new_n403));
  OAI21_X1  g217(.A(G131), .B1(new_n377), .B2(new_n378), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n380), .A2(new_n240), .A3(new_n376), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n406), .A3(new_n403), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT85), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n374), .B(new_n391), .C1(new_n405), .C2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT19), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n389), .B1(KEYINPUT84), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n389), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n398), .B1(new_n413), .B2(G146), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n404), .A2(new_n406), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n391), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n374), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n372), .B1(new_n409), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n391), .B1(new_n405), .B2(new_n408), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n417), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n423), .B2(new_n409), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT86), .B(G475), .Z(new_n425));
  OR2_X1    g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n303), .B1(new_n356), .B2(KEYINPUT92), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n370), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(G234), .A2(G237), .ZN(new_n430));
  INV_X1    g244(.A(G953), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n430), .A2(G952), .A3(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n430), .A2(G902), .A3(G953), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(G898), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G214), .B1(G237), .B2(G902), .ZN(new_n437));
  INV_X1    g251(.A(G119), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G116), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n310), .A2(G119), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT5), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n439), .A2(KEYINPUT5), .ZN(new_n443));
  INV_X1    g257(.A(G113), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT2), .B(G113), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n441), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n262), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n201), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n448), .A2(new_n441), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n449), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n224), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n451), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G122), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n451), .B(new_n457), .C1(new_n452), .C2(new_n455), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(KEYINPUT6), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n257), .A2(new_n462), .A3(new_n385), .A4(new_n247), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n257), .A2(new_n385), .A3(new_n247), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n221), .A2(new_n385), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G224), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n467), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n456), .A2(new_n472), .A3(new_n458), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n461), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n457), .B(KEYINPUT8), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n256), .B2(new_n450), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n442), .A2(KEYINPUT82), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT82), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n441), .A2(new_n478), .A3(KEYINPUT5), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n479), .A3(new_n445), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n262), .B1(new_n449), .B2(new_n480), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n476), .A2(new_n481), .B1(new_n467), .B2(KEYINPUT7), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT7), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n470), .B1(new_n467), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n262), .A2(new_n450), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n224), .A2(new_n454), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n488), .B2(new_n204), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n464), .B(KEYINPUT81), .C1(new_n385), .C2(new_n221), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n469), .B1(new_n490), .B2(new_n463), .ZN(new_n491));
  AND2_X1   g305(.A1(KEYINPUT83), .A2(KEYINPUT7), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n489), .A2(new_n457), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G210), .B1(G237), .B2(G902), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n474), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n474), .B2(new_n494), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n436), .B(new_n437), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n301), .A2(new_n429), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G472), .A2(G902), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT26), .B(G101), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n375), .A2(G210), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n220), .A2(new_n242), .A3(new_n222), .A4(new_n244), .ZN(new_n508));
  INV_X1    g322(.A(new_n454), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n240), .B1(G134), .B2(G137), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n348), .B2(G137), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n258), .A2(new_n241), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT28), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n242), .A2(new_n221), .A3(new_n244), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n509), .B1(new_n518), .B2(new_n512), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT28), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n512), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n454), .ZN(new_n524));
  AOI211_X1 g338(.A(new_n521), .B(new_n514), .C1(new_n524), .C2(new_n513), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n507), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n508), .A2(KEYINPUT30), .A3(new_n512), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n454), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n507), .A3(new_n513), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT31), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT31), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n531), .A2(new_n534), .A3(new_n507), .A4(new_n513), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n502), .B1(new_n527), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT32), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n508), .A2(new_n512), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n454), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n513), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n516), .B1(new_n542), .B2(KEYINPUT28), .ZN(new_n543));
  INV_X1    g357(.A(new_n507), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n514), .B1(new_n524), .B2(new_n513), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n515), .B1(new_n548), .B2(KEYINPUT69), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n549), .A2(new_n544), .A3(new_n525), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n531), .A2(new_n513), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n544), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n545), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n547), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G472), .ZN(new_n555));
  OAI211_X1 g369(.A(KEYINPUT32), .B(new_n502), .C1(new_n527), .C2(new_n536), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n539), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT70), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n539), .A2(new_n555), .A3(new_n559), .A4(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n438), .A2(G128), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n318), .A2(G119), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT24), .B(G110), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n318), .A2(KEYINPUT23), .A3(G119), .ZN(new_n566));
  INV_X1    g380(.A(new_n562), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n561), .B(new_n566), .C1(new_n567), .C2(KEYINPUT23), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n565), .B1(G110), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n400), .A2(new_n401), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n388), .B1(new_n397), .B2(G146), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n564), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n568), .B2(G110), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n571), .A2(new_n573), .A3(KEYINPUT72), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT72), .B1(new_n571), .B2(new_n573), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n570), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT22), .B(G137), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n431), .A2(G221), .A3(G234), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n570), .B(new_n579), .C1(new_n574), .C2(new_n575), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n294), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT25), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT25), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n581), .A2(new_n585), .A3(new_n294), .A4(new_n582), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n305), .B1(G234), .B2(new_n294), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(G902), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n581), .A2(new_n582), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT73), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n501), .A2(new_n558), .A3(new_n560), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  INV_X1    g408(.A(KEYINPUT93), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n281), .A2(new_n285), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n286), .A2(new_n291), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(G469), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n300), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n188), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n294), .B1(new_n527), .B2(new_n536), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(new_n537), .A3(new_n592), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n595), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n527), .A2(new_n536), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n606), .A2(new_n502), .B1(new_n602), .B2(G472), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n301), .A2(new_n607), .A3(KEYINPUT93), .A4(new_n592), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n427), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n367), .A2(KEYINPUT33), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n365), .A2(new_n612), .A3(new_n366), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(G478), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n302), .A2(new_n294), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n365), .B2(new_n366), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n302), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n499), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(KEYINPUT94), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT95), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n626));
  INV_X1    g440(.A(new_n419), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT20), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT96), .B1(new_n419), .B2(new_n420), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n627), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n426), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n616), .A2(new_n368), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n356), .A2(KEYINPUT92), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n303), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n428), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n626), .B1(new_n637), .B2(new_n499), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n370), .A2(new_n428), .ZN(new_n639));
  NOR4_X1   g453(.A1(new_n639), .A2(new_n498), .A3(new_n632), .A4(KEYINPUT97), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n609), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT35), .B(G107), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND3_X1  g458(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n645));
  OR3_X1    g459(.A1(new_n576), .A2(KEYINPUT36), .A3(new_n580), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n576), .B1(KEYINPUT36), .B2(new_n580), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n589), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n607), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n500), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n558), .A2(new_n560), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n437), .B(new_n649), .C1(new_n496), .C2(new_n497), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n432), .ZN(new_n658));
  INV_X1    g472(.A(new_n433), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n658), .B1(new_n659), .B2(G900), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n301), .A2(new_n637), .A3(new_n657), .A4(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n654), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n600), .A2(new_n657), .A3(new_n188), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n630), .A2(new_n426), .A3(new_n631), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n664), .B(new_n660), .C1(new_n370), .C2(new_n428), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n666), .A2(KEYINPUT98), .A3(new_n558), .A4(new_n560), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  XOR2_X1   g483(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n660), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n601), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n551), .A2(new_n507), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n294), .B1(new_n542), .B2(new_n507), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n539), .A2(new_n556), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n497), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n474), .A2(new_n494), .A3(new_n495), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n649), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n639), .A2(new_n610), .ZN(new_n687));
  AND4_X1   g501(.A1(new_n437), .A2(new_n685), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n674), .A2(new_n675), .A3(new_n680), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  INV_X1    g504(.A(new_n655), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n427), .A2(new_n614), .A3(new_n617), .A4(new_n660), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n663), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NOR2_X1   g509(.A1(new_n298), .A2(new_n299), .ZN(new_n696));
  OAI21_X1  g510(.A(G469), .B1(new_n696), .B2(G902), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n697), .A2(new_n188), .A3(new_n300), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n558), .A2(new_n698), .A3(new_n560), .A4(new_n592), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n620), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT41), .B(G113), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NOR2_X1   g516(.A1(new_n641), .A2(new_n699), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n310), .ZN(G18));
  NOR2_X1   g518(.A1(new_n686), .A2(new_n435), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n429), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n437), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n681), .B2(new_n682), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n697), .A2(new_n708), .A3(new_n188), .A4(new_n300), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n706), .A2(new_n710), .A3(new_n558), .A4(new_n560), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NAND2_X1  g526(.A1(new_n592), .A2(KEYINPUT101), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT101), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n588), .B2(new_n591), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n543), .A2(new_n507), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n502), .B1(new_n536), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n603), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n683), .A2(new_n437), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n639), .A2(new_n722), .A3(new_n610), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n721), .A2(new_n723), .A3(new_n436), .A4(new_n698), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT102), .B(G122), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G24));
  NOR4_X1   g540(.A1(new_n709), .A2(new_n720), .A3(new_n686), .A4(new_n692), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n385), .ZN(G27));
  INV_X1    g542(.A(new_n692), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n681), .A2(new_n437), .A3(new_n682), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n301), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n557), .A2(new_n716), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT42), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n600), .A2(new_n188), .A3(new_n731), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n558), .A3(new_n560), .A4(new_n592), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n240), .ZN(G33));
  INV_X1    g553(.A(new_n736), .ZN(new_n740));
  INV_X1    g554(.A(new_n665), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NOR2_X1   g557(.A1(new_n607), .A2(new_n686), .ZN(new_n744));
  INV_X1    g558(.A(new_n618), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n610), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT43), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(KEYINPUT103), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(KEYINPUT103), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n730), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n292), .A2(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n292), .A2(KEYINPUT45), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(G469), .A2(G902), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n300), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n757), .A2(new_n758), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n188), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n671), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n752), .B(new_n763), .C1(new_n751), .C2(new_n750), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  XNOR2_X1  g579(.A(new_n762), .B(KEYINPUT47), .ZN(new_n766));
  INV_X1    g580(.A(new_n592), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n655), .A2(new_n767), .A3(new_n729), .A4(new_n731), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n685), .A2(new_n437), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n698), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT111), .Z(new_n774));
  NOR4_X1   g588(.A1(new_n747), .A2(new_n658), .A3(new_n720), .A4(new_n717), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT50), .Z(new_n777));
  AND2_X1   g591(.A1(new_n697), .A2(new_n300), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n188), .B1(new_n778), .B2(KEYINPUT110), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(KEYINPUT110), .B2(new_n778), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n766), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n731), .A3(new_n775), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n698), .A2(new_n731), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT112), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n658), .B1(new_n784), .B2(KEYINPUT112), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n747), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT113), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n720), .A2(new_n686), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n680), .A2(new_n767), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n610), .A2(new_n787), .A3(new_n618), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n771), .B(new_n783), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n797), .B2(new_n796), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n771), .B1(new_n796), .B2(new_n783), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n787), .A2(new_n619), .A3(new_n793), .ZN(new_n801));
  INV_X1    g615(.A(G952), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n802), .B(G953), .C1(new_n775), .C2(new_n710), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n733), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n790), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT115), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT48), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n799), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n727), .B1(new_n691), .B2(new_n693), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n686), .A2(new_n660), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n301), .A2(KEYINPUT107), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT107), .B1(new_n301), .B2(new_n811), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n680), .B(new_n723), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n668), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n668), .A2(new_n810), .A3(new_n817), .A4(new_n814), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n724), .B(new_n711), .C1(new_n620), .C2(new_n699), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n738), .A3(new_n703), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT106), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT105), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n635), .A2(new_n823), .A3(new_n636), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT105), .B1(new_n370), .B2(new_n428), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n427), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n499), .B1(new_n826), .B2(new_n619), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n609), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n558), .A2(new_n560), .A3(new_n592), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n500), .B1(new_n829), .B2(new_n650), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n822), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n823), .B1(new_n635), .B2(new_n636), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n370), .A2(KEYINPUT105), .A3(new_n428), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n610), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n619), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n499), .A3(new_n605), .A4(new_n608), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(KEYINPUT106), .A3(new_n593), .A4(new_n651), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n791), .A2(new_n729), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n832), .A2(new_n833), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n649), .A2(new_n426), .A3(new_n660), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n631), .A3(new_n630), .A4(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n843), .B2(new_n655), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n844), .A2(new_n735), .B1(new_n741), .B2(new_n740), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n821), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(KEYINPUT108), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n850), .A2(new_n846), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n849), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  AND4_X1   g668(.A1(KEYINPUT53), .A2(new_n816), .A3(new_n818), .A4(new_n820), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT109), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n839), .A2(new_n856), .A3(new_n845), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n846), .A2(KEYINPUT109), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n851), .B1(new_n850), .B2(new_n846), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n854), .A2(new_n862), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n809), .A2(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n717), .A2(new_n746), .A3(new_n189), .A4(new_n707), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT104), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n778), .B(KEYINPUT49), .Z(new_n867));
  OR4_X1    g681(.A1(new_n680), .A2(new_n866), .A3(new_n685), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n864), .A2(new_n868), .ZN(G75));
  NOR2_X1   g683(.A1(new_n431), .A2(G952), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n859), .A2(new_n861), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(G210), .A3(G902), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n461), .A2(new_n473), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(new_n471), .Z(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT55), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n870), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT56), .B1(new_n872), .B2(KEYINPUT116), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n871), .A2(new_n879), .A3(G210), .A4(G902), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n881), .A2(KEYINPUT117), .A3(new_n875), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT117), .B1(new_n881), .B2(new_n875), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n886), .B(new_n877), .C1(new_n882), .C2(new_n883), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n887), .ZN(G51));
  XOR2_X1   g702(.A(new_n755), .B(KEYINPUT122), .Z(new_n889));
  AOI211_X1 g703(.A(new_n294), .B(new_n889), .C1(new_n859), .C2(new_n861), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n839), .A2(new_n856), .A3(new_n845), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n818), .A4(new_n820), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n856), .B1(new_n839), .B2(new_n845), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT54), .B1(new_n894), .B2(new_n848), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n896), .A3(new_n862), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n871), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n756), .B(KEYINPUT57), .Z(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n897), .A2(new_n902), .A3(new_n898), .A4(new_n899), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n696), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n890), .B1(new_n906), .B2(KEYINPUT121), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n870), .B1(new_n907), .B2(new_n909), .ZN(G54));
  NAND4_X1  g724(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n409), .A2(new_n418), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n870), .ZN(G60));
  NAND2_X1  g730(.A1(new_n611), .A2(new_n613), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n615), .B(KEYINPUT59), .Z(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n863), .B2(new_n918), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n917), .A2(new_n897), .A3(new_n898), .A4(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n870), .A3(new_n920), .ZN(G63));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n859), .B2(new_n861), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n646), .A2(new_n647), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n870), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n581), .A2(new_n582), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n927), .B1(new_n931), .B2(new_n925), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n929), .B(new_n932), .Z(G66));
  OAI21_X1  g747(.A(G953), .B1(new_n434), .B2(new_n468), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n703), .B(new_n819), .C1(new_n831), .C2(new_n838), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(G953), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n873), .B1(G898), .B2(new_n431), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G69));
  INV_X1    g752(.A(G900), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n283), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n763), .A2(new_n723), .A3(new_n805), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n668), .A2(new_n810), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI211_X1 g758(.A(new_n738), .B(new_n944), .C1(new_n741), .C2(new_n740), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n764), .A2(new_n769), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(G953), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n529), .A2(new_n530), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT124), .Z(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(new_n413), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n939), .A2(G953), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT126), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n943), .A2(new_n689), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT62), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n671), .B1(new_n834), .B2(new_n835), .ZN(new_n959));
  AOI211_X1 g773(.A(new_n946), .B(new_n958), .C1(new_n740), .C2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n952), .A2(new_n431), .ZN(new_n961));
  OAI221_X1 g775(.A(new_n941), .B1(new_n948), .B2(new_n955), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n962), .B(new_n963), .Z(G72));
  NAND2_X1  g778(.A1(new_n960), .A2(new_n935), .ZN(new_n965));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  AOI21_X1  g781(.A(new_n676), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n552), .A2(new_n532), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n853), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n945), .A2(new_n935), .A3(new_n947), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n507), .B(new_n551), .C1(new_n971), .C2(new_n967), .ZN(new_n972));
  NOR4_X1   g786(.A1(new_n968), .A2(new_n970), .A3(new_n870), .A4(new_n972), .ZN(G57));
endmodule


