

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578;

  XOR2_X1 U320 ( .A(KEYINPUT47), .B(n404), .Z(n288) );
  XNOR2_X1 U321 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U322 ( .A(n368), .B(n367), .ZN(n372) );
  NOR2_X1 U323 ( .A1(n515), .A2(n426), .ZN(n559) );
  XNOR2_X1 U324 ( .A(n377), .B(n376), .ZN(n566) );
  XNOR2_X1 U325 ( .A(n447), .B(KEYINPUT58), .ZN(n448) );
  XNOR2_X1 U326 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XOR2_X1 U327 ( .A(KEYINPUT82), .B(G92GAT), .Z(n290) );
  NAND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U329 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U330 ( .A(KEYINPUT84), .B(n291), .Z(n306) );
  XOR2_X1 U331 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n293) );
  XNOR2_X1 U332 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n292) );
  XOR2_X1 U333 ( .A(n293), .B(n292), .Z(n297) );
  XOR2_X1 U334 ( .A(KEYINPUT81), .B(KEYINPUT66), .Z(n295) );
  XNOR2_X1 U335 ( .A(G106GAT), .B(KEYINPUT65), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n299) );
  XOR2_X1 U338 ( .A(G50GAT), .B(G162GAT), .Z(n307) );
  XOR2_X1 U339 ( .A(G134GAT), .B(KEYINPUT83), .Z(n333) );
  XOR2_X1 U340 ( .A(n307), .B(n333), .Z(n298) );
  XNOR2_X1 U341 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U342 ( .A(G99GAT), .B(G85GAT), .Z(n364) );
  XNOR2_X1 U343 ( .A(n300), .B(n364), .ZN(n304) );
  XOR2_X1 U344 ( .A(G29GAT), .B(G43GAT), .Z(n302) );
  XNOR2_X1 U345 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n302), .B(n301), .ZN(n356) );
  XOR2_X1 U347 ( .A(G36GAT), .B(G190GAT), .Z(n412) );
  XNOR2_X1 U348 ( .A(n356), .B(n412), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n544) );
  INV_X1 U351 ( .A(n544), .ZN(n446) );
  XOR2_X1 U352 ( .A(G22GAT), .B(G155GAT), .Z(n393) );
  XNOR2_X1 U353 ( .A(n307), .B(n393), .ZN(n322) );
  XOR2_X1 U354 ( .A(G78GAT), .B(G148GAT), .Z(n309) );
  XNOR2_X1 U355 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n359) );
  XOR2_X1 U357 ( .A(n359), .B(KEYINPUT23), .Z(n311) );
  NAND2_X1 U358 ( .A1(G228GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U360 ( .A(G204GAT), .B(KEYINPUT92), .Z(n313) );
  XNOR2_X1 U361 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U363 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U364 ( .A(G211GAT), .B(KEYINPUT21), .Z(n317) );
  XNOR2_X1 U365 ( .A(G197GAT), .B(G218GAT), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n416) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n318), .B(KEYINPUT2), .ZN(n335) );
  XNOR2_X1 U369 ( .A(n416), .B(n335), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n459) );
  XOR2_X1 U372 ( .A(KEYINPUT4), .B(KEYINPUT94), .Z(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT93), .B(KEYINPUT6), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n341) );
  XOR2_X1 U375 ( .A(KEYINPUT1), .B(G57GAT), .Z(n326) );
  NAND2_X1 U376 ( .A1(G225GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U378 ( .A(KEYINPUT5), .B(n327), .ZN(n339) );
  XOR2_X1 U379 ( .A(G148GAT), .B(G155GAT), .Z(n329) );
  XNOR2_X1 U380 ( .A(G120GAT), .B(G162GAT), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U382 ( .A(n330), .B(G85GAT), .Z(n332) );
  XOR2_X1 U383 ( .A(G113GAT), .B(G1GAT), .Z(n344) );
  XNOR2_X1 U384 ( .A(G29GAT), .B(n344), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U386 ( .A(n334), .B(n333), .Z(n337) );
  XOR2_X1 U387 ( .A(KEYINPUT0), .B(G127GAT), .Z(n441) );
  XNOR2_X1 U388 ( .A(n441), .B(n335), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n515) );
  XOR2_X1 U392 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n343) );
  XNOR2_X1 U393 ( .A(KEYINPUT72), .B(KEYINPUT30), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U395 ( .A(G50GAT), .B(G36GAT), .Z(n346) );
  XOR2_X1 U396 ( .A(G169GAT), .B(G8GAT), .Z(n420) );
  XNOR2_X1 U397 ( .A(n344), .B(n420), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U399 ( .A(n348), .B(n347), .Z(n350) );
  NAND2_X1 U400 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U402 ( .A(KEYINPUT69), .B(G141GAT), .Z(n352) );
  XNOR2_X1 U403 ( .A(G197GAT), .B(G22GAT), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U405 ( .A(n354), .B(n353), .Z(n358) );
  XNOR2_X1 U406 ( .A(G15GAT), .B(KEYINPUT71), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n355), .B(KEYINPUT70), .ZN(n381) );
  XNOR2_X1 U408 ( .A(n356), .B(n381), .ZN(n357) );
  XOR2_X1 U409 ( .A(n358), .B(n357), .Z(n534) );
  XNOR2_X1 U410 ( .A(n359), .B(KEYINPUT79), .ZN(n361) );
  AND2_X1 U411 ( .A1(G230GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n361), .B(n360), .ZN(n368) );
  XOR2_X1 U413 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n363) );
  XNOR2_X1 U414 ( .A(KEYINPUT75), .B(KEYINPUT80), .ZN(n362) );
  XOR2_X1 U415 ( .A(n363), .B(n362), .Z(n366) );
  XOR2_X1 U416 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XNOR2_X1 U417 ( .A(n442), .B(n364), .ZN(n365) );
  XOR2_X1 U418 ( .A(KEYINPUT77), .B(KEYINPUT74), .Z(n370) );
  XNOR2_X1 U419 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n369) );
  XOR2_X1 U420 ( .A(n370), .B(n369), .Z(n371) );
  XNOR2_X1 U421 ( .A(n372), .B(n371), .ZN(n377) );
  XNOR2_X1 U422 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n373) );
  XNOR2_X1 U423 ( .A(n373), .B(KEYINPUT73), .ZN(n380) );
  XOR2_X1 U424 ( .A(G64GAT), .B(G92GAT), .Z(n375) );
  XNOR2_X1 U425 ( .A(G176GAT), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n375), .B(n374), .ZN(n413) );
  XNOR2_X1 U427 ( .A(n380), .B(n413), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n566), .B(KEYINPUT64), .ZN(n378) );
  XNOR2_X1 U429 ( .A(KEYINPUT41), .B(n378), .ZN(n549) );
  AND2_X1 U430 ( .A1(n534), .A2(n549), .ZN(n379) );
  XNOR2_X1 U431 ( .A(n379), .B(KEYINPUT46), .ZN(n403) );
  XNOR2_X1 U432 ( .A(n381), .B(n380), .ZN(n401) );
  XOR2_X1 U433 ( .A(G64GAT), .B(G183GAT), .Z(n383) );
  XNOR2_X1 U434 ( .A(G1GAT), .B(G8GAT), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U436 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n385) );
  XNOR2_X1 U437 ( .A(KEYINPUT85), .B(KEYINPUT89), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U439 ( .A(n387), .B(n386), .Z(n399) );
  XOR2_X1 U440 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n389) );
  XNOR2_X1 U441 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n397) );
  XOR2_X1 U443 ( .A(G78GAT), .B(G211GAT), .Z(n391) );
  XNOR2_X1 U444 ( .A(G71GAT), .B(G127GAT), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U446 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U447 ( .A1(G231GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U450 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U451 ( .A(n401), .B(n400), .Z(n541) );
  INV_X1 U452 ( .A(n541), .ZN(n571) );
  NAND2_X1 U453 ( .A1(n446), .A2(n571), .ZN(n402) );
  NOR2_X1 U454 ( .A1(n403), .A2(n402), .ZN(n404) );
  XOR2_X1 U455 ( .A(n544), .B(KEYINPUT36), .Z(n575) );
  NOR2_X1 U456 ( .A1(n571), .A2(n575), .ZN(n405) );
  XNOR2_X1 U457 ( .A(KEYINPUT45), .B(n405), .ZN(n406) );
  NAND2_X1 U458 ( .A1(n406), .A2(n566), .ZN(n407) );
  XOR2_X1 U459 ( .A(KEYINPUT109), .B(n407), .Z(n408) );
  NOR2_X1 U460 ( .A1(n534), .A2(n408), .ZN(n409) );
  XNOR2_X1 U461 ( .A(KEYINPUT110), .B(n409), .ZN(n410) );
  NOR2_X1 U462 ( .A1(n288), .A2(n410), .ZN(n411) );
  XNOR2_X1 U463 ( .A(n411), .B(KEYINPUT48), .ZN(n518) );
  XOR2_X1 U464 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U465 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U466 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U467 ( .A(n417), .B(n416), .Z(n422) );
  XOR2_X1 U468 ( .A(G183GAT), .B(KEYINPUT19), .Z(n419) );
  XNOR2_X1 U469 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n419), .B(n418), .ZN(n439) );
  XNOR2_X1 U471 ( .A(n420), .B(n439), .ZN(n421) );
  XOR2_X1 U472 ( .A(n422), .B(n421), .Z(n509) );
  INV_X1 U473 ( .A(n509), .ZN(n423) );
  NOR2_X1 U474 ( .A1(n518), .A2(n423), .ZN(n425) );
  XNOR2_X1 U475 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n424) );
  XOR2_X1 U476 ( .A(n425), .B(n424), .Z(n426) );
  NAND2_X1 U477 ( .A1(n459), .A2(n559), .ZN(n427) );
  XNOR2_X1 U478 ( .A(n427), .B(KEYINPUT55), .ZN(n445) );
  XOR2_X1 U479 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n429) );
  NAND2_X1 U480 ( .A1(G227GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U482 ( .A(n430), .B(KEYINPUT90), .Z(n438) );
  XOR2_X1 U483 ( .A(G134GAT), .B(G99GAT), .Z(n432) );
  XNOR2_X1 U484 ( .A(G43GAT), .B(G190GAT), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U486 ( .A(G176GAT), .B(G113GAT), .Z(n434) );
  XNOR2_X1 U487 ( .A(G169GAT), .B(G15GAT), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U491 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U492 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U493 ( .A(n444), .B(n443), .ZN(n519) );
  NAND2_X1 U494 ( .A1(n445), .A2(n519), .ZN(n556) );
  NOR2_X1 U495 ( .A1(n446), .A2(n556), .ZN(n449) );
  INV_X1 U496 ( .A(G190GAT), .ZN(n447) );
  NAND2_X1 U497 ( .A1(n566), .A2(n534), .ZN(n480) );
  NOR2_X1 U498 ( .A1(n571), .A2(n544), .ZN(n450) );
  XNOR2_X1 U499 ( .A(n450), .B(KEYINPUT16), .ZN(n467) );
  XOR2_X1 U500 ( .A(n509), .B(KEYINPUT95), .Z(n451) );
  XNOR2_X1 U501 ( .A(n451), .B(KEYINPUT27), .ZN(n516) );
  XNOR2_X1 U502 ( .A(n459), .B(KEYINPUT67), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n452), .B(KEYINPUT28), .ZN(n522) );
  NOR2_X1 U504 ( .A1(n522), .A2(n519), .ZN(n453) );
  NAND2_X1 U505 ( .A1(n516), .A2(n453), .ZN(n454) );
  NAND2_X1 U506 ( .A1(n515), .A2(n454), .ZN(n465) );
  AND2_X1 U507 ( .A1(n509), .A2(n519), .ZN(n455) );
  XNOR2_X1 U508 ( .A(KEYINPUT97), .B(n455), .ZN(n456) );
  NAND2_X1 U509 ( .A1(n456), .A2(n459), .ZN(n457) );
  XNOR2_X1 U510 ( .A(KEYINPUT25), .B(n457), .ZN(n458) );
  NOR2_X1 U511 ( .A1(n515), .A2(n458), .ZN(n463) );
  XNOR2_X1 U512 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n461) );
  NOR2_X1 U513 ( .A1(n519), .A2(n459), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n461), .B(n460), .ZN(n560) );
  NAND2_X1 U515 ( .A1(n560), .A2(n516), .ZN(n462) );
  NAND2_X1 U516 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U517 ( .A1(n465), .A2(n464), .ZN(n466) );
  XOR2_X1 U518 ( .A(KEYINPUT98), .B(n466), .Z(n476) );
  NAND2_X1 U519 ( .A1(n467), .A2(n476), .ZN(n496) );
  NOR2_X1 U520 ( .A1(n480), .A2(n496), .ZN(n474) );
  NAND2_X1 U521 ( .A1(n515), .A2(n474), .ZN(n470) );
  XOR2_X1 U522 ( .A(G1GAT), .B(KEYINPUT34), .Z(n468) );
  XNOR2_X1 U523 ( .A(KEYINPUT99), .B(n468), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n470), .B(n469), .ZN(G1324GAT) );
  NAND2_X1 U525 ( .A1(n509), .A2(n474), .ZN(n471) );
  XNOR2_X1 U526 ( .A(n471), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U527 ( .A(G15GAT), .B(KEYINPUT35), .Z(n473) );
  NAND2_X1 U528 ( .A1(n474), .A2(n519), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n473), .B(n472), .ZN(G1326GAT) );
  NAND2_X1 U530 ( .A1(n474), .A2(n522), .ZN(n475) );
  XNOR2_X1 U531 ( .A(n475), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 U532 ( .A(n476), .ZN(n477) );
  NOR2_X1 U533 ( .A1(n477), .A2(n575), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n478), .A2(n571), .ZN(n479) );
  XOR2_X1 U535 ( .A(KEYINPUT37), .B(n479), .Z(n505) );
  NOR2_X1 U536 ( .A1(n480), .A2(n505), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(KEYINPUT38), .ZN(n491) );
  NAND2_X1 U538 ( .A1(n515), .A2(n491), .ZN(n483) );
  XOR2_X1 U539 ( .A(G29GAT), .B(KEYINPUT39), .Z(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(G1328GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n485) );
  NAND2_X1 U542 ( .A1(n491), .A2(n509), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U544 ( .A(G36GAT), .B(n486), .ZN(G1329GAT) );
  XNOR2_X1 U545 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n490) );
  XOR2_X1 U546 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n488) );
  NAND2_X1 U547 ( .A1(n519), .A2(n491), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(G1330GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n493) );
  NAND2_X1 U551 ( .A1(n522), .A2(n491), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  XNOR2_X1 U554 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n498) );
  INV_X1 U555 ( .A(n534), .ZN(n562) );
  NAND2_X1 U556 ( .A1(n549), .A2(n562), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(KEYINPUT106), .ZN(n506) );
  NOR2_X1 U558 ( .A1(n506), .A2(n496), .ZN(n502) );
  NAND2_X1 U559 ( .A1(n502), .A2(n515), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1332GAT) );
  NAND2_X1 U561 ( .A1(n509), .A2(n502), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U563 ( .A(G71GAT), .B(KEYINPUT107), .Z(n501) );
  NAND2_X1 U564 ( .A1(n502), .A2(n519), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1334GAT) );
  XOR2_X1 U566 ( .A(G78GAT), .B(KEYINPUT43), .Z(n504) );
  NAND2_X1 U567 ( .A1(n502), .A2(n522), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  NOR2_X1 U569 ( .A1(n506), .A2(n505), .ZN(n512) );
  NAND2_X1 U570 ( .A1(n512), .A2(n515), .ZN(n507) );
  XNOR2_X1 U571 ( .A(KEYINPUT108), .B(n507), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G85GAT), .B(n508), .ZN(G1336GAT) );
  NAND2_X1 U573 ( .A1(n509), .A2(n512), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n519), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n522), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT44), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G106GAT), .B(n514), .ZN(G1339GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n517) );
  NOR2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n519), .A2(n532), .ZN(n520) );
  XOR2_X1 U583 ( .A(KEYINPUT111), .B(n520), .Z(n521) );
  NOR2_X1 U584 ( .A1(n522), .A2(n521), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n534), .A2(n528), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U587 ( .A(G120GAT), .B(KEYINPUT49), .Z(n525) );
  NAND2_X1 U588 ( .A1(n528), .A2(n549), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  NAND2_X1 U590 ( .A1(n541), .A2(n528), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(KEYINPUT50), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G127GAT), .B(n527), .ZN(G1342GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT51), .B(KEYINPUT112), .Z(n530) );
  NAND2_X1 U594 ( .A1(n528), .A2(n544), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G134GAT), .B(n531), .ZN(G1343GAT) );
  NAND2_X1 U597 ( .A1(n532), .A2(n560), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(KEYINPUT113), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n545), .A2(n534), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G141GAT), .B(n535), .ZN(G1344GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n537) );
  XNOR2_X1 U602 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U604 ( .A(KEYINPUT114), .B(n538), .Z(n540) );
  NAND2_X1 U605 ( .A1(n545), .A2(n549), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1345GAT) );
  NAND2_X1 U607 ( .A1(n541), .A2(n545), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(KEYINPUT116), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G155GAT), .B(n543), .ZN(G1346GAT) );
  XOR2_X1 U610 ( .A(G162GAT), .B(KEYINPUT117), .Z(n547) );
  NAND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1347GAT) );
  NOR2_X1 U613 ( .A1(n562), .A2(n556), .ZN(n548) );
  XOR2_X1 U614 ( .A(G169GAT), .B(n548), .Z(G1348GAT) );
  INV_X1 U615 ( .A(n549), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n550), .A2(n556), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n552) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(KEYINPUT119), .B(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  NOR2_X1 U622 ( .A1(n571), .A2(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1350GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT122), .ZN(n576) );
  NOR2_X1 U627 ( .A1(n562), .A2(n576), .ZN(n565) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1352GAT) );
  NOR2_X1 U631 ( .A1(n576), .A2(n566), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n568) );
  XNOR2_X1 U633 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n576), .ZN(n572) );
  XOR2_X1 U637 ( .A(G211GAT), .B(n572), .Z(G1354GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT62), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U639 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n578) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(n578), .B(n577), .Z(G1355GAT) );
endmodule

