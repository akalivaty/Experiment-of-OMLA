

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758;

  XNOR2_X1 U373 ( .A(n599), .B(KEYINPUT32), .ZN(n377) );
  NAND2_X1 U374 ( .A1(n625), .A2(n376), .ZN(n670) );
  XNOR2_X2 U375 ( .A(n448), .B(n478), .ZN(n376) );
  XNOR2_X2 U376 ( .A(n574), .B(n573), .ZN(n590) );
  XNOR2_X1 U377 ( .A(n465), .B(n464), .ZN(n474) );
  NAND2_X1 U378 ( .A1(n418), .A2(n471), .ZN(n470) );
  INV_X1 U379 ( .A(G953), .ZN(n743) );
  INV_X1 U380 ( .A(n470), .ZN(n658) );
  XNOR2_X2 U381 ( .A(n500), .B(n363), .ZN(n677) );
  AND2_X2 U382 ( .A1(n670), .A2(n371), .ZN(n466) );
  OR2_X2 U383 ( .A1(n600), .A2(n456), .ZN(n455) );
  INV_X2 U384 ( .A(n489), .ZN(n491) );
  XNOR2_X2 U385 ( .A(G116), .B(G119), .ZN(n489) );
  XNOR2_X2 U386 ( .A(n564), .B(KEYINPUT1), .ZN(n602) );
  XNOR2_X2 U387 ( .A(n554), .B(G469), .ZN(n564) );
  XNOR2_X2 U388 ( .A(KEYINPUT3), .B(KEYINPUT67), .ZN(n490) );
  XNOR2_X2 U389 ( .A(n566), .B(n463), .ZN(n751) );
  NAND2_X2 U390 ( .A1(n426), .A2(n425), .ZN(n566) );
  XNOR2_X2 U391 ( .A(n596), .B(n436), .ZN(n757) );
  INV_X1 U392 ( .A(n673), .ZN(n429) );
  INV_X1 U393 ( .A(KEYINPUT89), .ZN(n353) );
  NOR2_X1 U394 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U395 ( .A1(n414), .A2(n440), .ZN(n465) );
  NAND2_X1 U396 ( .A1(n480), .A2(n479), .ZN(n596) );
  AND2_X1 U397 ( .A1(n391), .A2(n390), .ZN(n389) );
  AND2_X1 U398 ( .A1(n481), .A2(n364), .ZN(n480) );
  AND2_X1 U399 ( .A1(n606), .A2(n428), .ZN(n599) );
  NAND2_X1 U400 ( .A1(n609), .A2(n437), .ZN(n593) );
  XNOR2_X1 U401 ( .A(n430), .B(n560), .ZN(n701) );
  AND2_X1 U402 ( .A1(n592), .A2(n438), .ZN(n437) );
  XNOR2_X1 U403 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X2 U404 ( .A1(G902), .A2(n725), .ZN(n543) );
  XNOR2_X1 U405 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U406 ( .A(n352), .B(n395), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n492), .B(n353), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n400), .B(n356), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n501), .B(KEYINPUT16), .ZN(n354) );
  XNOR2_X2 U410 ( .A(n413), .B(n350), .ZN(n636) );
  XNOR2_X2 U411 ( .A(n375), .B(n351), .ZN(n350) );
  XNOR2_X2 U412 ( .A(n355), .B(n354), .ZN(n375) );
  INV_X1 U413 ( .A(n517), .ZN(n356) );
  XNOR2_X2 U414 ( .A(n497), .B(n488), .ZN(n413) );
  XNOR2_X2 U415 ( .A(n740), .B(n487), .ZN(n497) );
  XNOR2_X2 U416 ( .A(n417), .B(n486), .ZN(n740) );
  XNOR2_X1 U417 ( .A(n609), .B(KEYINPUT90), .ZN(n612) );
  XNOR2_X2 U418 ( .A(n591), .B(KEYINPUT0), .ZN(n609) );
  INV_X1 U419 ( .A(n387), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n383), .B(n370), .ZN(n752) );
  NOR2_X1 U421 ( .A1(n431), .A2(n429), .ZN(n428) );
  BUF_X1 U422 ( .A(n572), .Z(n358) );
  NOR2_X2 U423 ( .A1(n636), .A2(n628), .ZN(n372) );
  XNOR2_X2 U424 ( .A(n455), .B(n369), .ZN(n700) );
  OR2_X1 U425 ( .A1(n565), .A2(n564), .ZN(n575) );
  AND2_X1 U426 ( .A1(n394), .A2(n662), .ZN(n393) );
  NAND2_X1 U427 ( .A1(n389), .A2(n386), .ZN(n392) );
  XNOR2_X1 U428 ( .A(n385), .B(KEYINPUT71), .ZN(n394) );
  INV_X1 U429 ( .A(G101), .ZN(n487) );
  XNOR2_X1 U430 ( .A(G134), .B(G131), .ZN(n741) );
  XOR2_X1 U431 ( .A(G137), .B(G140), .Z(n550) );
  XNOR2_X1 U432 ( .A(n741), .B(G146), .ZN(n552) );
  INV_X1 U433 ( .A(KEYINPUT38), .ZN(n419) );
  XNOR2_X1 U434 ( .A(n520), .B(n362), .ZN(n567) );
  NOR2_X1 U435 ( .A1(G902), .A2(n715), .ZN(n520) );
  NAND2_X1 U436 ( .A1(n388), .A2(n387), .ZN(n386) );
  NOR2_X1 U437 ( .A1(n751), .A2(n416), .ZN(n388) );
  NOR2_X1 U438 ( .A1(G902), .A2(G237), .ZN(n485) );
  XOR2_X1 U439 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n539) );
  INV_X1 U440 ( .A(KEYINPUT85), .ZN(n450) );
  AND2_X1 U441 ( .A1(G227), .A2(n743), .ZN(n484) );
  XNOR2_X1 U442 ( .A(n424), .B(G146), .ZN(n516) );
  INV_X1 U443 ( .A(G125), .ZN(n424) );
  XNOR2_X1 U444 ( .A(KEYINPUT18), .B(KEYINPUT76), .ZN(n396) );
  XNOR2_X1 U445 ( .A(G110), .B(KEYINPUT68), .ZN(n488) );
  XNOR2_X1 U446 ( .A(n399), .B(n397), .ZN(n492) );
  XNOR2_X1 U447 ( .A(KEYINPUT17), .B(KEYINPUT77), .ZN(n399) );
  NOR2_X1 U448 ( .A1(n398), .A2(G953), .ZN(n397) );
  INV_X1 U449 ( .A(KEYINPUT84), .ZN(n464) );
  XNOR2_X1 U450 ( .A(n435), .B(n427), .ZN(n498) );
  XNOR2_X1 U451 ( .A(n552), .B(n496), .ZN(n427) );
  XNOR2_X1 U452 ( .A(n535), .B(n378), .ZN(n739) );
  INV_X1 U453 ( .A(n550), .ZN(n378) );
  XOR2_X1 U454 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n510) );
  XNOR2_X1 U455 ( .A(KEYINPUT12), .B(KEYINPUT96), .ZN(n509) );
  XNOR2_X1 U456 ( .A(n516), .B(n476), .ZN(n535) );
  INV_X1 U457 ( .A(KEYINPUT10), .ZN(n476) );
  XOR2_X1 U458 ( .A(G131), .B(G140), .Z(n513) );
  NOR2_X1 U459 ( .A1(n690), .A2(n461), .ZN(n460) );
  INV_X1 U460 ( .A(KEYINPUT34), .ZN(n420) );
  AND2_X1 U461 ( .A1(n402), .A2(n360), .ZN(n556) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n402) );
  INV_X1 U463 ( .A(KEYINPUT30), .ZN(n403) );
  AND2_X1 U464 ( .A1(n677), .A2(n561), .ZN(n563) );
  INV_X2 U465 ( .A(n602), .ZN(n457) );
  INV_X1 U466 ( .A(KEYINPUT80), .ZN(n412) );
  INV_X1 U467 ( .A(KEYINPUT46), .ZN(n416) );
  NAND2_X1 U468 ( .A1(n361), .A2(n580), .ZN(n385) );
  NAND2_X1 U469 ( .A1(n409), .A2(n407), .ZN(n615) );
  NAND2_X1 U470 ( .A1(n470), .A2(n408), .ZN(n407) );
  AND2_X1 U471 ( .A1(n411), .A2(n410), .ZN(n409) );
  AND2_X1 U472 ( .A1(n548), .A2(KEYINPUT80), .ZN(n408) );
  XNOR2_X1 U473 ( .A(G902), .B(KEYINPUT15), .ZN(n537) );
  INV_X1 U474 ( .A(G224), .ZN(n398) );
  INV_X1 U475 ( .A(KEYINPUT48), .ZN(n415) );
  XNOR2_X1 U476 ( .A(G113), .B(G137), .ZN(n495) );
  INV_X1 U477 ( .A(KEYINPUT4), .ZN(n486) );
  XNOR2_X1 U478 ( .A(n439), .B(G107), .ZN(n501) );
  INV_X1 U479 ( .A(G122), .ZN(n439) );
  NOR2_X1 U480 ( .A1(G953), .A2(G237), .ZN(n511) );
  INV_X1 U481 ( .A(n537), .ZN(n628) );
  XNOR2_X1 U482 ( .A(n608), .B(n380), .ZN(n600) );
  INV_X1 U483 ( .A(KEYINPUT6), .ZN(n380) );
  NAND2_X1 U484 ( .A1(G234), .A2(G237), .ZN(n521) );
  NAND2_X1 U485 ( .A1(n677), .A2(n687), .ZN(n404) );
  NOR2_X1 U486 ( .A1(n429), .A2(n434), .ZN(n561) );
  NAND2_X1 U487 ( .A1(n360), .A2(n438), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n567), .B(n472), .ZN(n471) );
  INV_X1 U489 ( .A(KEYINPUT99), .ZN(n472) );
  INV_X1 U490 ( .A(n471), .ZN(n406) );
  XNOR2_X1 U491 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n478) );
  XNOR2_X1 U492 ( .A(n530), .B(n529), .ZN(n531) );
  INV_X1 U493 ( .A(KEYINPUT92), .ZN(n529) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n533) );
  INV_X1 U495 ( .A(KEYINPUT8), .ZN(n432) );
  NAND2_X1 U496 ( .A1(n743), .A2(G234), .ZN(n433) );
  XNOR2_X1 U497 ( .A(KEYINPUT100), .B(KEYINPUT9), .ZN(n405) );
  XNOR2_X1 U498 ( .A(G134), .B(KEYINPUT101), .ZN(n503) );
  XNOR2_X1 U499 ( .A(n553), .B(n459), .ZN(n458) );
  XNOR2_X1 U500 ( .A(n551), .B(G104), .ZN(n459) );
  NOR2_X1 U501 ( .A1(n571), .A2(n557), .ZN(n559) );
  XNOR2_X1 U502 ( .A(KEYINPUT65), .B(KEYINPUT19), .ZN(n573) );
  NAND2_X1 U503 ( .A1(n406), .A2(n568), .ZN(n548) );
  NOR2_X1 U504 ( .A1(n564), .A2(n601), .ZN(n611) );
  XNOR2_X1 U505 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U506 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U507 ( .A(n446), .B(n444), .ZN(n721) );
  XNOR2_X1 U508 ( .A(n445), .B(n502), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n504), .B(n447), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n503), .B(n405), .ZN(n445) );
  XNOR2_X1 U511 ( .A(n475), .B(n535), .ZN(n518) );
  NOR2_X1 U512 ( .A1(G952), .A2(n743), .ZN(n727) );
  XNOR2_X1 U513 ( .A(n443), .B(n442), .ZN(n441) );
  XNOR2_X1 U514 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n442) );
  NAND2_X1 U515 ( .A1(n555), .A2(n431), .ZN(n443) );
  INV_X1 U516 ( .A(KEYINPUT42), .ZN(n463) );
  INV_X1 U517 ( .A(n575), .ZN(n425) );
  NAND2_X1 U518 ( .A1(n584), .A2(n457), .ZN(n662) );
  XNOR2_X1 U519 ( .A(n583), .B(n379), .ZN(n584) );
  XNOR2_X1 U520 ( .A(KEYINPUT86), .B(KEYINPUT36), .ZN(n379) );
  INV_X1 U521 ( .A(n603), .ZN(n422) );
  INV_X1 U522 ( .A(KEYINPUT106), .ZN(n436) );
  BUF_X1 U523 ( .A(n602), .Z(n431) );
  OR2_X1 U524 ( .A1(n457), .A2(n594), .ZN(n359) );
  OR2_X1 U525 ( .A1(n588), .A2(n526), .ZN(n360) );
  AND2_X1 U526 ( .A1(n579), .A2(n401), .ZN(n361) );
  XOR2_X1 U527 ( .A(n508), .B(n507), .Z(n362) );
  XOR2_X1 U528 ( .A(n499), .B(G472), .Z(n363) );
  XNOR2_X1 U529 ( .A(n506), .B(n505), .ZN(n568) );
  INV_X1 U530 ( .A(n568), .ZN(n418) );
  AND2_X1 U531 ( .A1(n482), .A2(n595), .ZN(n364) );
  NOR2_X2 U532 ( .A1(n672), .A2(n673), .ZN(n679) );
  XOR2_X1 U533 ( .A(G143), .B(G122), .Z(n365) );
  AND2_X1 U534 ( .A1(n511), .A2(G210), .ZN(n366) );
  AND2_X1 U535 ( .A1(n663), .A2(KEYINPUT2), .ZN(n367) );
  AND2_X1 U536 ( .A1(n568), .A2(n412), .ZN(n368) );
  INV_X1 U537 ( .A(n440), .ZN(n664) );
  NAND2_X1 U538 ( .A1(n441), .A2(n581), .ZN(n440) );
  XNOR2_X1 U539 ( .A(KEYINPUT33), .B(KEYINPUT69), .ZN(n369) );
  XOR2_X1 U540 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n370) );
  OR2_X1 U541 ( .A1(n628), .A2(n627), .ZN(n371) );
  XNOR2_X2 U542 ( .A(n372), .B(n493), .ZN(n572) );
  AND2_X1 U543 ( .A1(n466), .A2(n467), .ZN(n373) );
  AND2_X2 U544 ( .A1(n466), .A2(n467), .ZN(n723) );
  NAND2_X1 U545 ( .A1(n468), .A2(n624), .ZN(n467) );
  NAND2_X1 U546 ( .A1(n752), .A2(n416), .ZN(n391) );
  XNOR2_X1 U547 ( .A(n381), .B(n415), .ZN(n414) );
  XNOR2_X1 U548 ( .A(n572), .B(n419), .ZN(n688) );
  XNOR2_X1 U549 ( .A(n607), .B(KEYINPUT103), .ZN(n754) );
  NOR2_X2 U550 ( .A1(n755), .A2(KEYINPUT44), .ZN(n604) );
  XNOR2_X1 U551 ( .A(n375), .B(n374), .ZN(n733) );
  INV_X1 U552 ( .A(KEYINPUT124), .ZN(n374) );
  NAND2_X1 U553 ( .A1(n622), .A2(n376), .ZN(n468) );
  NOR2_X1 U554 ( .A1(n376), .A2(KEYINPUT2), .ZN(n665) );
  NAND2_X1 U555 ( .A1(n376), .A2(n743), .ZN(n731) );
  NOR2_X2 U556 ( .A1(n757), .A2(n377), .ZN(n618) );
  XNOR2_X1 U557 ( .A(n377), .B(n756), .ZN(G21) );
  XNOR2_X1 U558 ( .A(n536), .B(n739), .ZN(n725) );
  NAND2_X1 U559 ( .A1(n392), .A2(n393), .ZN(n381) );
  OR2_X1 U560 ( .A1(n597), .A2(n359), .ZN(n479) );
  XNOR2_X2 U561 ( .A(n593), .B(KEYINPUT22), .ZN(n597) );
  NAND2_X1 U562 ( .A1(n751), .A2(n416), .ZN(n390) );
  INV_X1 U563 ( .A(n701), .ZN(n426) );
  NAND2_X2 U564 ( .A1(n382), .A2(n452), .ZN(n448) );
  NAND2_X1 U565 ( .A1(n449), .A2(n451), .ZN(n382) );
  NAND2_X1 U566 ( .A1(n723), .A2(G475), .ZN(n717) );
  NOR2_X2 U567 ( .A1(n597), .A2(n598), .ZN(n606) );
  NAND2_X1 U568 ( .A1(n585), .A2(n656), .ZN(n383) );
  XNOR2_X2 U569 ( .A(n384), .B(KEYINPUT35), .ZN(n755) );
  NAND2_X1 U570 ( .A1(n423), .A2(n422), .ZN(n384) );
  XNOR2_X1 U571 ( .A(n532), .B(n531), .ZN(n534) );
  XNOR2_X1 U572 ( .A(n534), .B(n483), .ZN(n536) );
  INV_X1 U573 ( .A(n752), .ZN(n387) );
  XNOR2_X1 U574 ( .A(n516), .B(n396), .ZN(n395) );
  XNOR2_X2 U575 ( .A(n491), .B(n490), .ZN(n400) );
  XNOR2_X1 U576 ( .A(n400), .B(n366), .ZN(n435) );
  INV_X1 U577 ( .A(n653), .ZN(n401) );
  NAND2_X1 U578 ( .A1(n658), .A2(n412), .ZN(n411) );
  INV_X1 U579 ( .A(n548), .ZN(n656) );
  NAND2_X1 U580 ( .A1(n368), .A2(n406), .ZN(n410) );
  NOR2_X1 U581 ( .A1(n658), .A2(n656), .ZN(n691) );
  XNOR2_X1 U582 ( .A(n413), .B(n458), .ZN(n708) );
  XNOR2_X1 U583 ( .A(n417), .B(KEYINPUT7), .ZN(n447) );
  XNOR2_X2 U584 ( .A(n477), .B(G143), .ZN(n417) );
  AND2_X2 U585 ( .A1(n453), .A2(n621), .ZN(n452) );
  XNOR2_X1 U586 ( .A(n618), .B(n450), .ZN(n449) );
  XNOR2_X1 U587 ( .A(n517), .B(n365), .ZN(n475) );
  XNOR2_X1 U588 ( .A(n421), .B(n420), .ZN(n423) );
  NAND2_X1 U589 ( .A1(n612), .A2(n454), .ZN(n421) );
  NOR2_X2 U590 ( .A1(n575), .A2(n590), .ZN(n654) );
  INV_X1 U591 ( .A(n672), .ZN(n438) );
  XNOR2_X1 U592 ( .A(n497), .B(n498), .ZN(n630) );
  INV_X1 U593 ( .A(n677), .ZN(n608) );
  NAND2_X1 U594 ( .A1(n723), .A2(G210), .ZN(n469) );
  XNOR2_X1 U595 ( .A(n469), .B(n639), .ZN(n640) );
  XNOR2_X1 U596 ( .A(n559), .B(n558), .ZN(n585) );
  NAND2_X1 U597 ( .A1(n688), .A2(n460), .ZN(n430) );
  NAND2_X1 U598 ( .A1(n556), .A2(n611), .ZN(n571) );
  XNOR2_X1 U599 ( .A(n604), .B(KEYINPUT66), .ZN(n451) );
  NAND2_X1 U600 ( .A1(n620), .A2(KEYINPUT44), .ZN(n453) );
  INV_X1 U601 ( .A(n700), .ZN(n454) );
  NAND2_X1 U602 ( .A1(n457), .A2(n679), .ZN(n456) );
  NAND2_X1 U603 ( .A1(n688), .A2(n687), .ZN(n462) );
  INV_X1 U604 ( .A(n687), .ZN(n461) );
  NOR2_X1 U605 ( .A1(n691), .A2(n462), .ZN(n692) );
  AND2_X2 U606 ( .A1(n474), .A2(n663), .ZN(n666) );
  NAND2_X1 U607 ( .A1(n474), .A2(n367), .ZN(n473) );
  XNOR2_X1 U608 ( .A(n473), .B(KEYINPUT83), .ZN(n625) );
  NAND2_X1 U609 ( .A1(n572), .A2(n687), .ZN(n574) );
  XNOR2_X2 U610 ( .A(KEYINPUT78), .B(G128), .ZN(n477) );
  NAND2_X1 U611 ( .A1(n597), .A2(n594), .ZN(n481) );
  NAND2_X1 U612 ( .A1(n457), .A2(n594), .ZN(n482) );
  NOR2_X2 U613 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U614 ( .A(n688), .ZN(n557) );
  AND2_X1 U615 ( .A1(G221), .A2(n533), .ZN(n483) );
  XNOR2_X1 U616 ( .A(n550), .B(n484), .ZN(n551) );
  INV_X1 U617 ( .A(KEYINPUT5), .ZN(n494) );
  XNOR2_X1 U618 ( .A(n495), .B(n494), .ZN(n496) );
  INV_X1 U619 ( .A(KEYINPUT39), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U621 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X2 U622 ( .A1(n633), .A2(n727), .ZN(n635) );
  XNOR2_X1 U623 ( .A(n485), .B(KEYINPUT73), .ZN(n546) );
  NAND2_X1 U624 ( .A1(n546), .A2(G210), .ZN(n493) );
  XOR2_X1 U625 ( .A(G113), .B(G104), .Z(n517) );
  NOR2_X1 U626 ( .A1(G902), .A2(n630), .ZN(n500) );
  XNOR2_X1 U627 ( .A(KEYINPUT70), .B(KEYINPUT94), .ZN(n499) );
  INV_X1 U628 ( .A(n600), .ZN(n598) );
  XNOR2_X1 U629 ( .A(G116), .B(n501), .ZN(n502) );
  NAND2_X1 U630 ( .A1(G217), .A2(n533), .ZN(n504) );
  NOR2_X1 U631 ( .A1(G902), .A2(n721), .ZN(n506) );
  XNOR2_X1 U632 ( .A(KEYINPUT102), .B(G478), .ZN(n505) );
  XOR2_X1 U633 ( .A(KEYINPUT98), .B(KEYINPUT13), .Z(n508) );
  XNOR2_X1 U634 ( .A(KEYINPUT97), .B(G475), .ZN(n507) );
  XNOR2_X1 U635 ( .A(n510), .B(n509), .ZN(n515) );
  NAND2_X1 U636 ( .A1(G214), .A2(n511), .ZN(n512) );
  XNOR2_X1 U637 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U638 ( .A(n515), .B(n514), .ZN(n519) );
  XNOR2_X1 U639 ( .A(n519), .B(n518), .ZN(n715) );
  XNOR2_X1 U640 ( .A(n521), .B(KEYINPUT14), .ZN(n522) );
  XNOR2_X1 U641 ( .A(KEYINPUT72), .B(n522), .ZN(n523) );
  NAND2_X1 U642 ( .A1(G952), .A2(n523), .ZN(n699) );
  NOR2_X1 U643 ( .A1(G953), .A2(n699), .ZN(n588) );
  AND2_X1 U644 ( .A1(n523), .A2(G953), .ZN(n524) );
  NAND2_X1 U645 ( .A1(G902), .A2(n524), .ZN(n586) );
  NOR2_X1 U646 ( .A1(G900), .A2(n586), .ZN(n525) );
  XNOR2_X1 U647 ( .A(n525), .B(KEYINPUT108), .ZN(n526) );
  XOR2_X1 U648 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n528) );
  XNOR2_X1 U649 ( .A(G128), .B(KEYINPUT23), .ZN(n527) );
  XNOR2_X1 U650 ( .A(n528), .B(n527), .ZN(n532) );
  XNOR2_X1 U651 ( .A(G119), .B(G110), .ZN(n530) );
  NAND2_X1 U652 ( .A1(G234), .A2(n537), .ZN(n538) );
  XNOR2_X1 U653 ( .A(n539), .B(n538), .ZN(n544) );
  NAND2_X1 U654 ( .A1(n544), .A2(G217), .ZN(n541) );
  XNOR2_X1 U655 ( .A(KEYINPUT25), .B(KEYINPUT75), .ZN(n540) );
  XNOR2_X2 U656 ( .A(n543), .B(n542), .ZN(n673) );
  NAND2_X1 U657 ( .A1(G221), .A2(n544), .ZN(n545) );
  XNOR2_X1 U658 ( .A(KEYINPUT21), .B(n545), .ZN(n672) );
  NAND2_X1 U659 ( .A1(G214), .A2(n546), .ZN(n687) );
  NAND2_X1 U660 ( .A1(n561), .A2(n687), .ZN(n547) );
  NOR2_X1 U661 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U662 ( .A1(n598), .A2(n549), .ZN(n582) );
  XNOR2_X1 U663 ( .A(n582), .B(KEYINPUT109), .ZN(n555) );
  XOR2_X1 U664 ( .A(n552), .B(G107), .Z(n553) );
  NOR2_X1 U665 ( .A1(n708), .A2(G902), .ZN(n554) );
  INV_X1 U666 ( .A(n679), .ZN(n601) );
  INV_X1 U667 ( .A(n358), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n568), .A2(n567), .ZN(n690) );
  XNOR2_X1 U669 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n560) );
  XNOR2_X1 U670 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n562) );
  XNOR2_X1 U671 ( .A(n563), .B(n562), .ZN(n565) );
  NOR2_X1 U672 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U673 ( .A(KEYINPUT107), .B(n569), .ZN(n603) );
  OR2_X1 U674 ( .A1(n603), .A2(n581), .ZN(n570) );
  NOR2_X1 U675 ( .A1(n571), .A2(n570), .ZN(n653) );
  INV_X1 U676 ( .A(n691), .ZN(n576) );
  NAND2_X1 U677 ( .A1(n576), .A2(n654), .ZN(n577) );
  NAND2_X1 U678 ( .A1(n577), .A2(KEYINPUT47), .ZN(n580) );
  NOR2_X1 U679 ( .A1(KEYINPUT47), .A2(n615), .ZN(n578) );
  NAND2_X1 U680 ( .A1(n578), .A2(n654), .ZN(n579) );
  NOR2_X1 U681 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U682 ( .A1(n658), .A2(n585), .ZN(n663) );
  XNOR2_X1 U683 ( .A(KEYINPUT74), .B(n666), .ZN(n622) );
  INV_X1 U684 ( .A(n690), .ZN(n592) );
  NOR2_X1 U685 ( .A1(G898), .A2(n586), .ZN(n587) );
  NOR2_X1 U686 ( .A1(n588), .A2(n587), .ZN(n589) );
  INV_X1 U687 ( .A(KEYINPUT105), .ZN(n594) );
  AND2_X1 U688 ( .A1(n673), .A2(n608), .ZN(n595) );
  NOR2_X1 U689 ( .A1(n457), .A2(n673), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n608), .A2(n456), .ZN(n684) );
  NAND2_X1 U692 ( .A1(n609), .A2(n684), .ZN(n610) );
  XNOR2_X1 U693 ( .A(n610), .B(KEYINPUT31), .ZN(n659) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n677), .A2(n613), .ZN(n643) );
  NOR2_X1 U696 ( .A1(n659), .A2(n643), .ZN(n614) );
  NOR2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n754), .A2(n616), .ZN(n617) );
  XNOR2_X1 U699 ( .A(n617), .B(KEYINPUT104), .ZN(n621) );
  INV_X1 U700 ( .A(n755), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U702 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n623) );
  AND2_X1 U703 ( .A1(n623), .A2(n628), .ZN(n624) );
  INV_X1 U704 ( .A(KEYINPUT2), .ZN(n626) );
  NOR2_X1 U705 ( .A1(KEYINPUT82), .A2(n626), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n723), .A2(G472), .ZN(n632) );
  XOR2_X1 U707 ( .A(KEYINPUT62), .B(KEYINPUT87), .Z(n629) );
  INV_X1 U708 ( .A(KEYINPUT63), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n635), .B(n634), .ZN(G57) );
  XNOR2_X1 U710 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT79), .ZN(n637) );
  NOR2_X2 U712 ( .A1(n640), .A2(n727), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n641), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U714 ( .A1(n656), .A2(n643), .ZN(n642) );
  XNOR2_X1 U715 ( .A(G104), .B(n642), .ZN(G6) );
  NAND2_X1 U716 ( .A1(n643), .A2(n658), .ZN(n649) );
  XOR2_X1 U717 ( .A(KEYINPUT116), .B(KEYINPUT27), .Z(n645) );
  XNOR2_X1 U718 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n645), .B(n644), .ZN(n647) );
  XOR2_X1 U720 ( .A(G107), .B(KEYINPUT26), .Z(n646) );
  XNOR2_X1 U721 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(G9) );
  XOR2_X1 U723 ( .A(KEYINPUT118), .B(KEYINPUT29), .Z(n651) );
  NAND2_X1 U724 ( .A1(n654), .A2(n658), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U726 ( .A(G128), .B(n652), .ZN(G30) );
  XOR2_X1 U727 ( .A(G143), .B(n653), .Z(G45) );
  NAND2_X1 U728 ( .A1(n654), .A2(n656), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(G146), .ZN(G48) );
  NAND2_X1 U730 ( .A1(n659), .A2(n656), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(G113), .ZN(G15) );
  NAND2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(G116), .ZN(G18) );
  XOR2_X1 U734 ( .A(G125), .B(KEYINPUT37), .Z(n661) );
  XNOR2_X1 U735 ( .A(n662), .B(n661), .ZN(G27) );
  XNOR2_X1 U736 ( .A(G134), .B(n663), .ZN(G36) );
  XOR2_X1 U737 ( .A(G140), .B(n664), .Z(G42) );
  XOR2_X1 U738 ( .A(KEYINPUT81), .B(n665), .Z(n668) );
  NOR2_X1 U739 ( .A1(n666), .A2(KEYINPUT2), .ZN(n667) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n671), .A2(n743), .ZN(n706) );
  XOR2_X1 U743 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n675) );
  NAND2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U747 ( .A(KEYINPUT120), .B(n678), .Z(n682) );
  NOR2_X1 U748 ( .A1(n679), .A2(n457), .ZN(n680) );
  XNOR2_X1 U749 ( .A(KEYINPUT50), .B(n680), .ZN(n681) );
  NOR2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U752 ( .A(KEYINPUT51), .B(n685), .Z(n686) );
  NOR2_X1 U753 ( .A1(n701), .A2(n686), .ZN(n696) );
  NOR2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n693) );
  NOR2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U757 ( .A1(n694), .A2(n700), .ZN(n695) );
  NOR2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U759 ( .A(n697), .B(KEYINPUT52), .ZN(n698) );
  NOR2_X1 U760 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U761 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U763 ( .A(n704), .B(KEYINPUT121), .ZN(n705) );
  XNOR2_X1 U764 ( .A(KEYINPUT53), .B(n707), .ZN(G75) );
  XOR2_X1 U765 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n710) );
  XNOR2_X1 U766 ( .A(n708), .B(KEYINPUT122), .ZN(n709) );
  XNOR2_X1 U767 ( .A(n710), .B(n709), .ZN(n712) );
  NAND2_X1 U768 ( .A1(n373), .A2(G469), .ZN(n711) );
  XNOR2_X1 U769 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U770 ( .A1(n727), .A2(n713), .ZN(G54) );
  XOR2_X1 U771 ( .A(KEYINPUT59), .B(KEYINPUT88), .Z(n714) );
  NOR2_X2 U772 ( .A1(n718), .A2(n727), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n719), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U774 ( .A1(G478), .A2(n373), .ZN(n720) );
  XNOR2_X1 U775 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U776 ( .A1(n727), .A2(n722), .ZN(G63) );
  NAND2_X1 U777 ( .A1(G217), .A2(n373), .ZN(n724) );
  XNOR2_X1 U778 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n727), .A2(n726), .ZN(G66) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n728) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n728), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n737) );
  XNOR2_X1 U784 ( .A(G101), .B(G110), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n733), .B(n732), .ZN(n735) );
  NOR2_X1 U786 ( .A1(G898), .A2(n743), .ZN(n734) );
  NOR2_X1 U787 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U788 ( .A(n737), .B(n736), .ZN(n738) );
  XOR2_X1 U789 ( .A(KEYINPUT123), .B(n738), .Z(G69) );
  XNOR2_X1 U790 ( .A(n740), .B(n739), .ZN(n742) );
  XNOR2_X1 U791 ( .A(n742), .B(n741), .ZN(n745) );
  XOR2_X1 U792 ( .A(n745), .B(n666), .Z(n744) );
  NAND2_X1 U793 ( .A1(n744), .A2(n743), .ZN(n749) );
  XNOR2_X1 U794 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U796 ( .A1(G953), .A2(n747), .ZN(n748) );
  NAND2_X1 U797 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U798 ( .A(G137), .B(KEYINPUT126), .Z(n750) );
  XNOR2_X1 U799 ( .A(n751), .B(n750), .ZN(G39) );
  XNOR2_X1 U800 ( .A(n357), .B(G131), .ZN(n753) );
  XNOR2_X1 U801 ( .A(n753), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U802 ( .A(n754), .B(G101), .Z(G3) );
  XOR2_X1 U803 ( .A(n755), .B(G122), .Z(G24) );
  XNOR2_X1 U804 ( .A(G119), .B(KEYINPUT125), .ZN(n756) );
  XNOR2_X1 U805 ( .A(G110), .B(KEYINPUT117), .ZN(n758) );
  XNOR2_X1 U806 ( .A(n758), .B(n757), .ZN(G12) );
endmodule

