//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n451, new_n454,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(G173));
  XNOR2_X1  g024(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n450));
  AND2_X1   g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  NAND2_X1  g027(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n451), .A2(G2106), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  NOR4_X1   g032(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  INV_X1    g035(.A(G2106), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OAI22_X1  g037(.A1(new_n457), .A2(new_n461), .B1(new_n462), .B2(new_n458), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n465), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT68), .ZN(new_n478));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n479), .A2(new_n480), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  OR3_X1    g062(.A1(new_n478), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n478), .B2(new_n486), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n466), .B2(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n484), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n512), .A2(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n510), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  OR2_X1    g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n504), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT70), .B(G51), .Z(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n515), .A2(new_n514), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n511), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n532), .A2(new_n536), .ZN(G168));
  AND2_X1   g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n507), .B2(G64), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n509), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n512), .A2(new_n541), .B1(new_n518), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(new_n525), .A2(G43), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n507), .A2(new_n511), .A3(G81), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(new_n509), .ZN(new_n548));
  INV_X1    g123(.A(G860), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  INV_X1    g131(.A(G78), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n533), .A2(new_n556), .B1(new_n557), .B2(new_n504), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n523), .A2(new_n524), .B1(new_n505), .B2(new_n506), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n558), .A2(G651), .B1(new_n559), .B2(G91), .ZN(new_n560));
  OAI211_X1 g135(.A(G53), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n559), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n525), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n507), .B2(G61), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT72), .B1(new_n572), .B2(new_n509), .ZN(new_n573));
  OAI21_X1  g148(.A(G61), .B1(new_n515), .B2(new_n514), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(new_n570), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(new_n576), .A3(G651), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n559), .A2(G86), .B1(new_n525), .B2(G48), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n509), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n512), .A2(new_n582), .B1(new_n518), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n581), .A2(new_n584), .ZN(G290));
  INV_X1    g160(.A(G868), .ZN(new_n586));
  NOR2_X1   g161(.A1(G301), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT10), .B1(new_n518), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n505), .B2(new_n506), .ZN(new_n591));
  AND2_X1   g166(.A1(G79), .A2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n525), .A2(G54), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n507), .A2(new_n511), .A3(new_n595), .A4(G92), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n589), .A2(new_n593), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT73), .Z(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n587), .B1(new_n599), .B2(new_n586), .ZN(G284));
  AOI21_X1  g175(.A(new_n587), .B1(new_n599), .B2(new_n586), .ZN(G321));
  NOR2_X1   g176(.A1(G286), .A2(new_n586), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT9), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n561), .B(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n507), .A2(new_n511), .A3(G91), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n557), .A2(new_n504), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n507), .B2(G65), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n607), .B2(new_n509), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT74), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n602), .B1(new_n610), .B2(new_n586), .ZN(G297));
  AOI21_X1  g186(.A(new_n602), .B1(new_n610), .B2(new_n586), .ZN(G280));
  AOI21_X1  g187(.A(new_n598), .B1(G559), .B2(new_n549), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT75), .ZN(G148));
  NAND2_X1  g189(.A1(new_n548), .A2(new_n586), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n598), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n586), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n484), .A2(new_n472), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT76), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n625), .A2(KEYINPUT77), .B1(new_n626), .B2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(KEYINPUT77), .B2(new_n625), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n481), .A2(G135), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n484), .A2(G123), .A3(G2105), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  OAI211_X1 g207(.A(new_n624), .B(new_n632), .C1(new_n622), .C2(new_n621), .ZN(G156));
  INV_X1    g208(.A(G14), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  INV_X1    g210(.A(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2430), .Z(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT78), .B(KEYINPUT14), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n634), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT79), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n647), .A2(new_n652), .A3(new_n649), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n647), .B2(new_n649), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT17), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT80), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT81), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n658), .A2(new_n660), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n657), .A2(new_n659), .ZN(new_n666));
  OR3_X1    g241(.A1(new_n665), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n662), .A2(new_n657), .A3(new_n659), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(KEYINPUT82), .ZN(new_n676));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(KEYINPUT82), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n673), .A2(new_n674), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n678), .B2(new_n675), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n678), .A2(KEYINPUT83), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n686), .B(new_n687), .Z(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n686), .B(new_n687), .ZN(new_n692));
  INV_X1    g267(.A(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n690), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n691), .B1(new_n690), .B2(new_n694), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT87), .Z(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  OR2_X1    g277(.A1(G6), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G305), .B2(new_n698), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  AOI22_X1  g280(.A1(new_n701), .A2(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n702), .B2(new_n701), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n698), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(G288), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n698), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT33), .B(G1976), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n704), .B2(new_n705), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n707), .A2(KEYINPUT34), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT34), .B1(new_n707), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n481), .A2(G131), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n465), .A2(G107), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n718));
  INV_X1    g293(.A(G119), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n716), .B1(new_n717), .B2(new_n718), .C1(new_n719), .C2(new_n485), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT84), .ZN(new_n721));
  MUX2_X1   g296(.A(G25), .B(new_n721), .S(G29), .Z(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(KEYINPUT85), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(KEYINPUT85), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G24), .ZN(new_n727));
  INV_X1    g302(.A(G290), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT86), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1986), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n725), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n714), .A2(new_n715), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT36), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G32), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT26), .Z(new_n738));
  INV_X1    g313(.A(G129), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n485), .B2(new_n739), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n736), .B1(new_n744), .B2(new_n735), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT27), .ZN(new_n746));
  INV_X1    g321(.A(G1996), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n698), .A2(G4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n599), .B2(new_n698), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G1348), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n750), .A2(G1348), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n748), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G168), .A2(new_n698), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n698), .B2(G21), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT90), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n735), .B1(new_n759), .B2(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n759), .B2(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G160), .B2(G29), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G2084), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT91), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n755), .A2(new_n756), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n735), .A2(G33), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n481), .A2(G139), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n768), .B(new_n769), .C1(new_n465), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n766), .B1(new_n771), .B2(G29), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(new_n442), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n698), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n698), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(G1961), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n765), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n758), .A2(new_n764), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n698), .A2(G19), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT88), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n545), .A2(new_n546), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n507), .A2(G56), .ZN(new_n782));
  NAND2_X1  g357(.A1(G68), .A2(G543), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n509), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n780), .B1(new_n785), .B2(new_n698), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1341), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n698), .A2(G20), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT23), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G299), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT93), .B(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n481), .A2(G140), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n465), .A2(G116), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n795));
  INV_X1    g370(.A(G128), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n793), .B1(new_n794), .B2(new_n795), .C1(new_n796), .C2(new_n485), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G29), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n735), .A2(G26), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT28), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT89), .B(G2067), .Z(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n735), .A2(G27), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT92), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G164), .B2(new_n735), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n803), .B1(new_n443), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n806), .A2(G2078), .B1(new_n762), .B2(G2084), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT30), .B(G28), .ZN(new_n810));
  OR2_X1    g385(.A1(KEYINPUT31), .A2(G11), .ZN(new_n811));
  NAND2_X1  g386(.A1(KEYINPUT31), .A2(G11), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n810), .A2(new_n735), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n631), .B2(new_n735), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n772), .B2(new_n442), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n802), .A2(new_n801), .B1(new_n775), .B2(G1961), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n808), .A2(new_n809), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n778), .A2(new_n787), .A3(new_n792), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(G29), .A2(G35), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G162), .B2(G29), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT29), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(G2090), .Z(new_n822));
  NAND4_X1  g397(.A1(new_n734), .A2(new_n753), .A3(new_n818), .A4(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  OAI211_X1 g399(.A(G55), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n825));
  INV_X1    g400(.A(G93), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n518), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(G67), .B1(new_n515), .B2(new_n514), .ZN(new_n828));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n509), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n549), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT37), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n599), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n785), .A2(new_n837), .A3(new_n831), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT95), .B1(new_n827), .B2(new_n830), .ZN(new_n839));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n505), .B2(new_n506), .ZN(new_n841));
  INV_X1    g416(.A(new_n829), .ZN(new_n842));
  OAI21_X1  g417(.A(G651), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n507), .A2(new_n511), .A3(G93), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n843), .A2(new_n837), .A3(new_n825), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n839), .A2(new_n548), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n838), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n836), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT96), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n549), .B1(new_n848), .B2(KEYINPUT39), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n833), .B1(new_n850), .B2(new_n851), .ZN(G145));
  INV_X1    g427(.A(G160), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n488), .B2(new_n489), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n631), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n488), .A2(new_n853), .A3(new_n489), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n856), .B1(new_n855), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT99), .ZN(new_n861));
  INV_X1    g436(.A(G130), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n465), .A2(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n485), .A2(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(G142), .B2(new_n481), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n620), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n720), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(KEYINPUT98), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n499), .A2(new_n501), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n491), .A2(new_n494), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n771), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n743), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n797), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n797), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(G164), .A3(new_n876), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n869), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n861), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n879), .A2(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n869), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n884), .A2(new_n868), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n879), .A2(new_n881), .A3(new_n868), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n887), .B(new_n888), .C1(new_n858), .C2(new_n859), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g466(.A(new_n586), .B1(new_n827), .B2(new_n830), .ZN(new_n892));
  AND4_X1   g467(.A1(new_n593), .A2(new_n589), .A3(new_n594), .A4(new_n596), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(G299), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT100), .B1(new_n609), .B2(new_n597), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(G299), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(KEYINPUT101), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n609), .A2(KEYINPUT100), .A3(new_n597), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n896), .B1(new_n893), .B2(G299), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n894), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n905), .A2(KEYINPUT41), .A3(new_n906), .A4(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n898), .A2(new_n906), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n616), .B(new_n847), .ZN(new_n912));
  MUX2_X1   g487(.A(new_n902), .B(new_n911), .S(new_n912), .Z(new_n913));
  NOR2_X1   g488(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(G290), .B(G305), .Z(new_n916));
  XNOR2_X1  g491(.A(G303), .B(new_n709), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(KEYINPUT102), .B2(KEYINPUT42), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n915), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n892), .B1(new_n920), .B2(new_n586), .ZN(G295));
  OAI21_X1  g496(.A(new_n892), .B1(new_n920), .B2(new_n586), .ZN(G331));
  INV_X1    g497(.A(new_n918), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n924));
  OAI22_X1  g499(.A1(new_n540), .A2(new_n543), .B1(new_n532), .B2(new_n536), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n539), .A2(new_n509), .ZN(new_n926));
  INV_X1    g501(.A(new_n536), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n525), .A2(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n559), .A2(G90), .B1(new_n525), .B2(G52), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  AND4_X1   g505(.A1(new_n838), .A2(new_n846), .A3(new_n925), .A4(new_n930), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n838), .A2(new_n846), .B1(new_n930), .B2(new_n925), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT104), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n925), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(new_n847), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n911), .A2(new_n924), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n847), .B(new_n935), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n901), .B2(new_n900), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n907), .A2(new_n910), .B1(new_n933), .B2(new_n936), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(new_n924), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n923), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G37), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n940), .B1(new_n943), .B2(new_n924), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n911), .A2(new_n937), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT105), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n950), .A3(new_n918), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT106), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n948), .A2(new_n950), .A3(new_n953), .A4(new_n918), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n947), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n939), .A2(KEYINPUT41), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n939), .B1(new_n959), .B2(new_n909), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n937), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n963), .B2(new_n902), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n946), .B1(new_n964), .B2(new_n918), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(new_n952), .B2(new_n954), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n957), .B(KEYINPUT44), .C1(new_n958), .C2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n952), .A2(new_n954), .ZN(new_n970));
  INV_X1    g545(.A(new_n965), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n970), .A2(new_n956), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n945), .A2(new_n946), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n956), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n968), .B(new_n969), .C1(new_n972), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n956), .A3(new_n971), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n955), .B2(new_n956), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n968), .B1(new_n978), .B2(new_n969), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n967), .B1(new_n976), .B2(new_n979), .ZN(G397));
  NOR2_X1   g555(.A1(G290), .A2(G1986), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT108), .B(G1384), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(G164), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(G160), .A2(G40), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(G1986), .A3(G290), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT110), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n743), .B(new_n747), .ZN(new_n993));
  INV_X1    g568(.A(G2067), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n797), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n723), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n720), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n987), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n992), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G303), .A2(G8), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n872), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n986), .B1(new_n1005), .B2(new_n983), .ZN(new_n1006));
  INV_X1    g581(.A(new_n984), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n872), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1971), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G40), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n470), .A2(new_n474), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n870), .B2(new_n871), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1014), .A2(new_n1015), .A3(G2090), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1003), .B(G8), .C1(new_n1009), .C2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n872), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1011), .B1(new_n1012), .B2(KEYINPUT45), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n756), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1025));
  INV_X1    g600(.A(G2084), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1011), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT114), .B(new_n756), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1023), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G286), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1017), .A2(KEYINPUT63), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n709), .A2(G1976), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1012), .A2(new_n1011), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(G8), .ZN(new_n1036));
  AOI211_X1 g611(.A(KEYINPUT111), .B(new_n1030), .C1(new_n1012), .C2(new_n1011), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1033), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT112), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n1033), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(KEYINPUT52), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  AOI211_X1 g619(.A(KEYINPUT72), .B(new_n509), .C1(new_n574), .C2(new_n570), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n1046));
  INV_X1    g621(.A(G86), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n518), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1044), .B1(new_n1049), .B2(new_n573), .ZN(new_n1050));
  AND4_X1   g625(.A1(new_n1044), .A2(new_n573), .A3(new_n577), .A4(new_n578), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1043), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G305), .A2(G1981), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1044), .A3(new_n573), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(KEYINPUT49), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1052), .B(new_n1055), .C1(new_n1037), .C2(new_n1036), .ZN(new_n1056));
  INV_X1    g631(.A(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1033), .B(new_n1058), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1003), .ZN(new_n1061));
  OAI21_X1  g636(.A(G8), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1042), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1032), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1042), .A2(new_n1060), .A3(new_n1063), .A4(KEYINPUT115), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n1038), .B2(KEYINPUT112), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1068), .B1(new_n1041), .B2(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n1017), .A4(new_n1063), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1066), .A2(new_n1067), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1056), .A2(new_n1057), .A3(new_n709), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1054), .B(KEYINPUT113), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1078), .A2(new_n1079), .B1(new_n1037), .B2(new_n1036), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT116), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1032), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1067), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1081), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1082), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1006), .A2(new_n1092), .A3(new_n443), .A4(new_n1018), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n983), .B1(G164), .B2(G1384), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1094), .A2(new_n1018), .A3(new_n443), .A4(new_n1011), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1093), .A2(new_n1096), .A3(KEYINPUT53), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1099));
  INV_X1    g674(.A(G1961), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1024), .A2(new_n1025), .A3(KEYINPUT118), .A4(new_n1011), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1103));
  NAND3_X1  g678(.A1(new_n1094), .A2(new_n1011), .A3(new_n1008), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(G2078), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(G171), .B1(new_n1097), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT123), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1109), .B(G171), .C1(new_n1097), .C2(new_n1106), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n985), .A2(new_n1008), .A3(new_n1011), .A4(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1102), .A2(new_n1105), .A3(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1108), .A2(new_n1110), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n560), .B2(KEYINPUT117), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G299), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n560), .B(new_n562), .C1(KEYINPUT117), .C2(KEYINPUT57), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1094), .A2(new_n1008), .A3(new_n1011), .A4(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1119), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1348), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1099), .A2(new_n1127), .A3(new_n1101), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1012), .A2(new_n994), .A3(new_n1011), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n598), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1123), .B1(new_n1119), .B2(new_n1125), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1126), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(KEYINPUT60), .A3(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n598), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1128), .A2(KEYINPUT60), .A3(new_n599), .A4(new_n1129), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1134), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1126), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(new_n1131), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1131), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(KEYINPUT61), .A3(new_n1126), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1012), .B2(new_n1011), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT119), .B(G1996), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1094), .A2(new_n1008), .A3(new_n1011), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1006), .A2(KEYINPUT120), .A3(new_n1008), .A4(new_n1149), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1145), .B1(new_n1154), .B2(new_n785), .ZN(new_n1155));
  AOI211_X1 g730(.A(KEYINPUT59), .B(new_n548), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1142), .B(new_n1144), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1132), .B1(new_n1139), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1029), .A2(G286), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(G8), .B1(new_n1029), .B2(G286), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT51), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1028), .A2(new_n1027), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1006), .A2(new_n1018), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT114), .B1(new_n1164), .B2(new_n756), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1030), .B1(new_n1166), .B2(G168), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT51), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1042), .A2(new_n1060), .A3(new_n1063), .A4(new_n1017), .ZN(new_n1171));
  OR3_X1    g746(.A1(new_n1097), .A2(new_n1106), .A3(G171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1116), .B1(new_n1113), .B2(G171), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1117), .A2(new_n1158), .A3(new_n1170), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1168), .B1(new_n1167), .B2(new_n1159), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1161), .A2(KEYINPUT51), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT62), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1162), .A2(new_n1179), .A3(new_n1169), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1171), .B1(new_n1110), .B2(new_n1108), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1175), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1000), .B1(new_n1091), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT48), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n989), .B(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1186), .B1(new_n1187), .B2(new_n999), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n999), .A2(new_n1187), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n721), .A2(new_n997), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n996), .A2(new_n1190), .B1(G2067), .B2(new_n797), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1188), .A2(new_n1189), .B1(new_n987), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n987), .A2(new_n747), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT46), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n995), .A2(new_n744), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n987), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT47), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1192), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT125), .ZN(new_n1200));
  OAI21_X1  g775(.A(KEYINPUT126), .B1(new_n1184), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1199), .B(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1175), .A2(new_n1182), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n1090), .B2(new_n1082), .ZN(new_n1206));
  OAI211_X1 g781(.A(new_n1202), .B(new_n1204), .C1(new_n1206), .C2(new_n1000), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1201), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g783(.A1(G227), .A2(new_n463), .ZN(new_n1210));
  OAI211_X1 g784(.A(new_n655), .B(new_n1210), .C1(new_n695), .C2(new_n696), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1211), .B1(new_n886), .B2(new_n889), .ZN(new_n1212));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1213));
  OAI211_X1 g787(.A(new_n1212), .B(new_n1213), .C1(new_n972), .C2(new_n974), .ZN(new_n1214));
  INV_X1    g788(.A(new_n1214), .ZN(new_n1215));
  AOI21_X1  g789(.A(new_n1213), .B1(new_n978), .B2(new_n1212), .ZN(new_n1216));
  NOR2_X1   g790(.A1(new_n1215), .A2(new_n1216), .ZN(G308));
  NAND2_X1  g791(.A1(new_n978), .A2(new_n1212), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1218), .A2(KEYINPUT127), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1219), .A2(new_n1214), .ZN(G225));
endmodule


