

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U557 ( .A1(n668), .A2(n548), .ZN(n657) );
  XOR2_X1 U558 ( .A(n558), .B(KEYINPUT75), .Z(n1021) );
  NOR2_X1 U559 ( .A1(n766), .A2(n765), .ZN(n768) );
  XOR2_X1 U560 ( .A(n789), .B(KEYINPUT99), .Z(n525) );
  INV_X1 U561 ( .A(KEYINPUT30), .ZN(n737) );
  XNOR2_X1 U562 ( .A(n738), .B(n737), .ZN(n739) );
  AND2_X1 U563 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U564 ( .A(KEYINPUT32), .B(KEYINPUT96), .ZN(n767) );
  XNOR2_X1 U565 ( .A(n768), .B(n767), .ZN(n782) );
  NOR2_X1 U566 ( .A1(n824), .A2(n823), .ZN(n825) );
  INV_X1 U567 ( .A(G2105), .ZN(n579) );
  AND2_X1 U568 ( .A1(n579), .A2(G2104), .ZN(n912) );
  NAND2_X1 U569 ( .A1(G102), .A2(n912), .ZN(n528) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XOR2_X2 U571 ( .A(n526), .B(KEYINPUT17), .Z(n913) );
  NAND2_X1 U572 ( .A1(G138), .A2(n913), .ZN(n527) );
  NAND2_X1 U573 ( .A1(n528), .A2(n527), .ZN(n533) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n908) );
  NAND2_X1 U575 ( .A1(n908), .A2(G114), .ZN(n531) );
  NOR2_X1 U576 ( .A1(n579), .A2(G2104), .ZN(n529) );
  XNOR2_X2 U577 ( .A(n529), .B(KEYINPUT66), .ZN(n909) );
  NAND2_X1 U578 ( .A1(G126), .A2(n909), .ZN(n530) );
  NAND2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U580 ( .A1(n533), .A2(n532), .ZN(G164) );
  XOR2_X1 U581 ( .A(G2438), .B(G2454), .Z(n535) );
  XNOR2_X1 U582 ( .A(G2435), .B(G2430), .ZN(n534) );
  XNOR2_X1 U583 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U584 ( .A(n536), .B(KEYINPUT106), .Z(n538) );
  XNOR2_X1 U585 ( .A(G1348), .B(G1341), .ZN(n537) );
  XNOR2_X1 U586 ( .A(n538), .B(n537), .ZN(n542) );
  XOR2_X1 U587 ( .A(G2446), .B(G2451), .Z(n540) );
  XNOR2_X1 U588 ( .A(G2443), .B(G2427), .ZN(n539) );
  XNOR2_X1 U589 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U590 ( .A(n542), .B(n541), .Z(n543) );
  AND2_X1 U591 ( .A1(G14), .A2(n543), .ZN(G401) );
  INV_X1 U592 ( .A(G651), .ZN(n548) );
  NOR2_X1 U593 ( .A1(G543), .A2(n548), .ZN(n544) );
  XOR2_X2 U594 ( .A(KEYINPUT1), .B(n544), .Z(n667) );
  NAND2_X1 U595 ( .A1(G56), .A2(n667), .ZN(n545) );
  XNOR2_X1 U596 ( .A(n545), .B(KEYINPUT73), .ZN(n546) );
  XNOR2_X1 U597 ( .A(n546), .B(KEYINPUT14), .ZN(n553) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U599 ( .A1(n654), .A2(G81), .ZN(n547) );
  XNOR2_X1 U600 ( .A(n547), .B(KEYINPUT12), .ZN(n550) );
  XOR2_X1 U601 ( .A(KEYINPUT0), .B(G543), .Z(n668) );
  NAND2_X1 U602 ( .A1(G68), .A2(n657), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U604 ( .A(KEYINPUT13), .B(n551), .Z(n552) );
  NOR2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U606 ( .A(n554), .B(KEYINPUT74), .ZN(n557) );
  NOR2_X1 U607 ( .A1(G651), .A2(n668), .ZN(n555) );
  XOR2_X1 U608 ( .A(KEYINPUT65), .B(n555), .Z(n663) );
  NAND2_X1 U609 ( .A1(G43), .A2(n663), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n558) );
  INV_X1 U611 ( .A(G860), .ZN(n610) );
  OR2_X1 U612 ( .A1(n1021), .A2(n610), .ZN(G153) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  INV_X1 U614 ( .A(G82), .ZN(G220) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G120), .ZN(G236) );
  NAND2_X1 U617 ( .A1(G64), .A2(n667), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G52), .A2(n663), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n566) );
  NAND2_X1 U620 ( .A1(G90), .A2(n654), .ZN(n562) );
  NAND2_X1 U621 ( .A1(G77), .A2(n657), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  XNOR2_X1 U624 ( .A(KEYINPUT70), .B(n564), .ZN(n565) );
  NOR2_X1 U625 ( .A1(n566), .A2(n565), .ZN(G171) );
  INV_X1 U626 ( .A(G171), .ZN(G301) );
  NAND2_X1 U627 ( .A1(n654), .A2(G89), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G76), .A2(n657), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT5), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n667), .A2(G63), .ZN(n571) );
  XNOR2_X1 U633 ( .A(n571), .B(KEYINPUT78), .ZN(n573) );
  NAND2_X1 U634 ( .A1(G51), .A2(n663), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT6), .B(n574), .Z(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U638 ( .A(n577), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(G125), .A2(n909), .ZN(n583) );
  AND2_X1 U641 ( .A1(G2104), .A2(G101), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U643 ( .A(n580), .B(KEYINPUT67), .ZN(n581) );
  XNOR2_X1 U644 ( .A(n581), .B(KEYINPUT23), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U646 ( .A(n584), .B(KEYINPUT68), .ZN(n700) );
  NAND2_X1 U647 ( .A1(G137), .A2(n913), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G113), .A2(n908), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n698) );
  NOR2_X1 U650 ( .A1(n700), .A2(n698), .ZN(G160) );
  NAND2_X1 U651 ( .A1(G94), .A2(G452), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n588), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U655 ( .A(G223), .B(KEYINPUT72), .Z(n849) );
  NAND2_X1 U656 ( .A1(n849), .A2(G567), .ZN(n589) );
  XOR2_X1 U657 ( .A(KEYINPUT11), .B(n589), .Z(G234) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U659 ( .A1(G92), .A2(n654), .ZN(n591) );
  NAND2_X1 U660 ( .A1(G66), .A2(n667), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U662 ( .A(KEYINPUT76), .B(n592), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G79), .A2(n657), .ZN(n594) );
  NAND2_X1 U664 ( .A1(G54), .A2(n663), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n598) );
  XNOR2_X1 U667 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n598), .B(n597), .ZN(n857) );
  INV_X1 U669 ( .A(n857), .ZN(n1024) );
  INV_X1 U670 ( .A(G868), .ZN(n607) );
  NAND2_X1 U671 ( .A1(n1024), .A2(n607), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U673 ( .A1(G65), .A2(n667), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G53), .A2(n663), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G91), .A2(n654), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G78), .A2(n657), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n1008) );
  INV_X1 U680 ( .A(n1008), .ZN(G299) );
  NOR2_X1 U681 ( .A1(G868), .A2(G299), .ZN(n609) );
  NOR2_X1 U682 ( .A1(G286), .A2(n607), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n610), .A2(G559), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n611), .A2(n857), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n612), .B(KEYINPUT16), .ZN(n613) );
  XOR2_X1 U687 ( .A(KEYINPUT79), .B(n613), .Z(G148) );
  NAND2_X1 U688 ( .A1(n857), .A2(G868), .ZN(n614) );
  NOR2_X1 U689 ( .A1(G559), .A2(n614), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n615), .B(KEYINPUT80), .ZN(n617) );
  NOR2_X1 U691 ( .A1(n1021), .A2(G868), .ZN(n616) );
  NOR2_X1 U692 ( .A1(n617), .A2(n616), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G99), .A2(n912), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT82), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G111), .A2(n908), .ZN(n619) );
  XOR2_X1 U696 ( .A(KEYINPUT81), .B(n619), .Z(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n909), .A2(G123), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(KEYINPUT18), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n913), .A2(G135), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n944) );
  XNOR2_X1 U703 ( .A(n944), .B(G2096), .ZN(n628) );
  INV_X1 U704 ( .A(G2100), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(G156) );
  NAND2_X1 U706 ( .A1(G559), .A2(n857), .ZN(n629) );
  XNOR2_X1 U707 ( .A(n629), .B(KEYINPUT83), .ZN(n678) );
  XOR2_X1 U708 ( .A(n1021), .B(n678), .Z(n630) );
  NOR2_X1 U709 ( .A1(G860), .A2(n630), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n663), .A2(G55), .ZN(n631) );
  XNOR2_X1 U711 ( .A(n631), .B(KEYINPUT86), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G67), .A2(n667), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G93), .A2(n654), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G80), .A2(n657), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT85), .B(n636), .Z(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n680) );
  XOR2_X1 U719 ( .A(n639), .B(n680), .Z(n640) );
  XOR2_X1 U720 ( .A(KEYINPUT84), .B(n640), .Z(G145) );
  NAND2_X1 U721 ( .A1(G88), .A2(n654), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G75), .A2(n657), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G62), .A2(n667), .ZN(n644) );
  NAND2_X1 U725 ( .A1(G50), .A2(n663), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U727 ( .A1(n646), .A2(n645), .ZN(G166) );
  NAND2_X1 U728 ( .A1(G85), .A2(n654), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G72), .A2(n657), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n663), .A2(G47), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n667), .A2(G60), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U735 ( .A(KEYINPUT69), .B(n653), .ZN(G290) );
  NAND2_X1 U736 ( .A1(G86), .A2(n654), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G61), .A2(n667), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n657), .A2(G73), .ZN(n658) );
  XOR2_X1 U740 ( .A(KEYINPUT2), .B(n658), .Z(n659) );
  NOR2_X1 U741 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n663), .A2(G48), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n662), .A2(n661), .ZN(G305) );
  NAND2_X1 U744 ( .A1(G49), .A2(n663), .ZN(n665) );
  NAND2_X1 U745 ( .A1(G74), .A2(G651), .ZN(n664) );
  NAND2_X1 U746 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U747 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U748 ( .A1(n668), .A2(G87), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n670), .A2(n669), .ZN(G288) );
  XNOR2_X1 U750 ( .A(G166), .B(n1008), .ZN(n676) );
  XNOR2_X1 U751 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n672) );
  XOR2_X1 U752 ( .A(G305), .B(G288), .Z(n671) );
  XNOR2_X1 U753 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U754 ( .A(n680), .B(n673), .Z(n674) );
  XNOR2_X1 U755 ( .A(G290), .B(n674), .ZN(n675) );
  XNOR2_X1 U756 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U757 ( .A(n677), .B(n1021), .ZN(n856) );
  XNOR2_X1 U758 ( .A(n678), .B(n856), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n679), .A2(G868), .ZN(n682) );
  OR2_X1 U760 ( .A1(G868), .A2(n680), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n682), .A2(n681), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2078), .A2(G2084), .ZN(n683) );
  XOR2_X1 U763 ( .A(KEYINPUT20), .B(n683), .Z(n684) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n684), .ZN(n685) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n685), .ZN(n686) );
  NAND2_X1 U766 ( .A1(n686), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U767 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U768 ( .A1(G236), .A2(G237), .ZN(n687) );
  NAND2_X1 U769 ( .A1(G69), .A2(n687), .ZN(n688) );
  XNOR2_X1 U770 ( .A(KEYINPUT89), .B(n688), .ZN(n689) );
  NAND2_X1 U771 ( .A1(n689), .A2(G108), .ZN(n855) );
  NAND2_X1 U772 ( .A1(n855), .A2(G567), .ZN(n695) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n690) );
  XOR2_X1 U774 ( .A(KEYINPUT22), .B(n690), .Z(n691) );
  NOR2_X1 U775 ( .A1(G218), .A2(n691), .ZN(n692) );
  NAND2_X1 U776 ( .A1(G96), .A2(n692), .ZN(n854) );
  NAND2_X1 U777 ( .A1(G2106), .A2(n854), .ZN(n693) );
  XNOR2_X1 U778 ( .A(KEYINPUT88), .B(n693), .ZN(n694) );
  NAND2_X1 U779 ( .A1(n695), .A2(n694), .ZN(n929) );
  NAND2_X1 U780 ( .A1(G483), .A2(G661), .ZN(n696) );
  NOR2_X1 U781 ( .A1(n929), .A2(n696), .ZN(n853) );
  NAND2_X1 U782 ( .A1(n853), .A2(G36), .ZN(G176) );
  INV_X1 U783 ( .A(G166), .ZN(G303) );
  INV_X1 U784 ( .A(KEYINPUT33), .ZN(n772) );
  NOR2_X1 U785 ( .A1(G1976), .A2(G288), .ZN(n705) );
  INV_X1 U786 ( .A(G40), .ZN(n697) );
  OR2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n699) );
  OR2_X1 U788 ( .A1(n700), .A2(n699), .ZN(n810) );
  NOR2_X1 U789 ( .A1(G164), .A2(G1384), .ZN(n701) );
  INV_X1 U790 ( .A(n701), .ZN(n809) );
  NOR2_X2 U791 ( .A1(n810), .A2(n809), .ZN(n731) );
  INV_X1 U792 ( .A(n731), .ZN(n749) );
  NAND2_X1 U793 ( .A1(n749), .A2(G8), .ZN(n779) );
  INV_X1 U794 ( .A(n779), .ZN(n786) );
  NAND2_X1 U795 ( .A1(n705), .A2(n786), .ZN(n702) );
  NOR2_X1 U796 ( .A1(n772), .A2(n702), .ZN(n703) );
  XNOR2_X1 U797 ( .A(n703), .B(KEYINPUT97), .ZN(n775) );
  NOR2_X1 U798 ( .A1(G1971), .A2(G303), .ZN(n704) );
  NOR2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n1013) );
  NOR2_X1 U800 ( .A1(n749), .A2(G2084), .ZN(n706) );
  XNOR2_X1 U801 ( .A(n706), .B(KEYINPUT94), .ZN(n734) );
  NAND2_X1 U802 ( .A1(n734), .A2(G8), .ZN(n748) );
  NOR2_X1 U803 ( .A1(G1966), .A2(n779), .ZN(n746) );
  AND2_X1 U804 ( .A1(n731), .A2(G1996), .ZN(n707) );
  XOR2_X1 U805 ( .A(n707), .B(KEYINPUT26), .Z(n709) );
  NAND2_X1 U806 ( .A1(n749), .A2(G1341), .ZN(n708) );
  NAND2_X1 U807 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U808 ( .A1(n1021), .A2(n710), .ZN(n711) );
  XOR2_X1 U809 ( .A(n711), .B(KEYINPUT64), .Z(n715) );
  XOR2_X1 U810 ( .A(KEYINPUT95), .B(n749), .Z(n730) );
  INV_X1 U811 ( .A(n730), .ZN(n719) );
  NAND2_X1 U812 ( .A1(G2067), .A2(n719), .ZN(n713) );
  NAND2_X1 U813 ( .A1(G1348), .A2(n749), .ZN(n712) );
  NAND2_X1 U814 ( .A1(n713), .A2(n712), .ZN(n716) );
  OR2_X1 U815 ( .A1(n1024), .A2(n716), .ZN(n714) );
  NAND2_X1 U816 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U817 ( .A1(n1024), .A2(n716), .ZN(n717) );
  NAND2_X1 U818 ( .A1(n718), .A2(n717), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n719), .A2(G2072), .ZN(n720) );
  XNOR2_X1 U820 ( .A(n720), .B(KEYINPUT27), .ZN(n722) );
  AND2_X1 U821 ( .A1(G1956), .A2(n730), .ZN(n721) );
  NOR2_X1 U822 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U823 ( .A1(n725), .A2(n1008), .ZN(n723) );
  NAND2_X1 U824 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U825 ( .A1(n725), .A2(n1008), .ZN(n726) );
  XOR2_X1 U826 ( .A(n726), .B(KEYINPUT28), .Z(n727) );
  NAND2_X1 U827 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U828 ( .A(n729), .B(KEYINPUT29), .ZN(n758) );
  XOR2_X1 U829 ( .A(G2078), .B(KEYINPUT25), .Z(n961) );
  NOR2_X1 U830 ( .A1(n961), .A2(n730), .ZN(n733) );
  NOR2_X1 U831 ( .A1(n731), .A2(G1961), .ZN(n732) );
  NOR2_X1 U832 ( .A1(n733), .A2(n732), .ZN(n740) );
  NOR2_X1 U833 ( .A1(G301), .A2(n740), .ZN(n756) );
  NOR2_X1 U834 ( .A1(n758), .A2(n756), .ZN(n744) );
  INV_X1 U835 ( .A(n734), .ZN(n735) );
  NAND2_X1 U836 ( .A1(G8), .A2(n735), .ZN(n736) );
  NOR2_X1 U837 ( .A1(n746), .A2(n736), .ZN(n738) );
  NOR2_X1 U838 ( .A1(G168), .A2(n739), .ZN(n742) );
  AND2_X1 U839 ( .A1(G301), .A2(n740), .ZN(n741) );
  NOR2_X1 U840 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U841 ( .A(n743), .B(KEYINPUT31), .ZN(n759) );
  NOR2_X1 U842 ( .A1(n744), .A2(n759), .ZN(n745) );
  NOR2_X1 U843 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U844 ( .A1(n748), .A2(n747), .ZN(n780) );
  INV_X1 U845 ( .A(G8), .ZN(n754) );
  NOR2_X1 U846 ( .A1(G1971), .A2(n779), .ZN(n751) );
  NOR2_X1 U847 ( .A1(G2090), .A2(n749), .ZN(n750) );
  NOR2_X1 U848 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U849 ( .A1(n752), .A2(G303), .ZN(n753) );
  NOR2_X1 U850 ( .A1(n754), .A2(n753), .ZN(n760) );
  OR2_X1 U851 ( .A1(n760), .A2(G286), .ZN(n764) );
  INV_X1 U852 ( .A(n764), .ZN(n755) );
  OR2_X1 U853 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U854 ( .A1(n758), .A2(n757), .ZN(n766) );
  INV_X1 U855 ( .A(n759), .ZN(n762) );
  INV_X1 U856 ( .A(n760), .ZN(n761) );
  NAND2_X1 U857 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U858 ( .A1(n780), .A2(n782), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n1013), .A2(n769), .ZN(n771) );
  AND2_X1 U860 ( .A1(G288), .A2(G1976), .ZN(n1012) );
  NOR2_X1 U861 ( .A1(n1012), .A2(n779), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U865 ( .A(G1981), .B(G305), .ZN(n1017) );
  NOR2_X1 U866 ( .A1(n776), .A2(n1017), .ZN(n792) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XNOR2_X1 U868 ( .A(n777), .B(KEYINPUT24), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n778), .A2(n786), .ZN(n790) );
  AND2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n788) );
  NOR2_X1 U872 ( .A1(G2090), .A2(G303), .ZN(n783) );
  NAND2_X1 U873 ( .A1(G8), .A2(n783), .ZN(n784) );
  XNOR2_X1 U874 ( .A(n784), .B(KEYINPUT98), .ZN(n785) );
  OR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n787) );
  AND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n525), .ZN(n791) );
  NOR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n824) );
  NAND2_X1 U879 ( .A1(n908), .A2(G107), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G119), .A2(n909), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G95), .A2(n912), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G131), .A2(n913), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n797) );
  OR2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n898) );
  NAND2_X1 U886 ( .A1(n898), .A2(G1991), .ZN(n807) );
  NAND2_X1 U887 ( .A1(n908), .A2(G117), .ZN(n800) );
  NAND2_X1 U888 ( .A1(G129), .A2(n909), .ZN(n799) );
  NAND2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n912), .A2(G105), .ZN(n801) );
  XOR2_X1 U891 ( .A(KEYINPUT38), .B(n801), .Z(n802) );
  NOR2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n913), .A2(G141), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n899) );
  NAND2_X1 U895 ( .A1(G1996), .A2(n899), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n808), .B(KEYINPUT93), .ZN(n939) );
  INV_X1 U898 ( .A(n939), .ZN(n811) );
  NOR2_X1 U899 ( .A1(n701), .A2(n810), .ZN(n843) );
  NAND2_X1 U900 ( .A1(n811), .A2(n843), .ZN(n829) );
  NAND2_X1 U901 ( .A1(G104), .A2(n912), .ZN(n813) );
  NAND2_X1 U902 ( .A1(G140), .A2(n913), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U904 ( .A(KEYINPUT34), .B(n814), .ZN(n820) );
  NAND2_X1 U905 ( .A1(n908), .A2(G116), .ZN(n815) );
  XOR2_X1 U906 ( .A(KEYINPUT91), .B(n815), .Z(n817) );
  NAND2_X1 U907 ( .A1(G128), .A2(n909), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U909 ( .A(n818), .B(KEYINPUT35), .Z(n819) );
  NOR2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U911 ( .A(KEYINPUT36), .B(n821), .Z(n822) );
  XNOR2_X1 U912 ( .A(KEYINPUT92), .B(n822), .ZN(n895) );
  XOR2_X1 U913 ( .A(KEYINPUT37), .B(G2067), .Z(n839) );
  AND2_X1 U914 ( .A1(n895), .A2(n839), .ZN(n942) );
  NAND2_X1 U915 ( .A1(n843), .A2(n942), .ZN(n837) );
  NAND2_X1 U916 ( .A1(n829), .A2(n837), .ZN(n823) );
  XNOR2_X1 U917 ( .A(n825), .B(KEYINPUT100), .ZN(n828) );
  XNOR2_X1 U918 ( .A(KEYINPUT90), .B(G1986), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n826), .B(G290), .ZN(n1030) );
  NAND2_X1 U920 ( .A1(n1030), .A2(n843), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n847) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n899), .ZN(n935) );
  INV_X1 U923 ( .A(n829), .ZN(n834) );
  NOR2_X1 U924 ( .A1(G1991), .A2(n898), .ZN(n830) );
  XNOR2_X1 U925 ( .A(KEYINPUT102), .B(n830), .ZN(n943) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n831) );
  XOR2_X1 U927 ( .A(n831), .B(KEYINPUT101), .Z(n832) );
  NOR2_X1 U928 ( .A1(n943), .A2(n832), .ZN(n833) );
  NOR2_X1 U929 ( .A1(n834), .A2(n833), .ZN(n835) );
  NOR2_X1 U930 ( .A1(n935), .A2(n835), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n836), .B(KEYINPUT39), .ZN(n838) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(n841) );
  NOR2_X1 U933 ( .A1(n895), .A2(n839), .ZN(n840) );
  XNOR2_X1 U934 ( .A(n840), .B(KEYINPUT103), .ZN(n950) );
  NAND2_X1 U935 ( .A1(n841), .A2(n950), .ZN(n842) );
  XNOR2_X1 U936 ( .A(KEYINPUT104), .B(n842), .ZN(n844) );
  NAND2_X1 U937 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U938 ( .A(KEYINPUT105), .B(n845), .Z(n846) );
  NAND2_X1 U939 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U940 ( .A(n848), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U941 ( .A1(n849), .A2(G2106), .ZN(n850) );
  XOR2_X1 U942 ( .A(KEYINPUT107), .B(n850), .Z(G217) );
  AND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U944 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U946 ( .A1(n853), .A2(n852), .ZN(G188) );
  INV_X1 U948 ( .A(G108), .ZN(G238) );
  INV_X1 U949 ( .A(G96), .ZN(G221) );
  NOR2_X1 U950 ( .A1(n855), .A2(n854), .ZN(G325) );
  INV_X1 U951 ( .A(G325), .ZN(G261) );
  XOR2_X1 U952 ( .A(KEYINPUT113), .B(n856), .Z(n859) );
  XNOR2_X1 U953 ( .A(G171), .B(n857), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U955 ( .A(n860), .B(G286), .ZN(n861) );
  NOR2_X1 U956 ( .A1(G37), .A2(n861), .ZN(G397) );
  XOR2_X1 U957 ( .A(G2100), .B(G2096), .Z(n863) );
  XNOR2_X1 U958 ( .A(KEYINPUT42), .B(G2678), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U960 ( .A(KEYINPUT43), .B(G2072), .Z(n865) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2090), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U963 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U964 ( .A(G2078), .B(G2084), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n869), .B(n868), .ZN(G227) );
  XOR2_X1 U966 ( .A(G1956), .B(G1961), .Z(n871) );
  XNOR2_X1 U967 ( .A(G1986), .B(G1981), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U969 ( .A(n872), .B(G2474), .Z(n874) );
  XNOR2_X1 U970 ( .A(G1976), .B(G1971), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U972 ( .A(KEYINPUT41), .B(G1966), .Z(n876) );
  XNOR2_X1 U973 ( .A(G1991), .B(G1996), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(G229) );
  NAND2_X1 U976 ( .A1(G100), .A2(n912), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G112), .A2(n908), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U979 ( .A1(n909), .A2(G124), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n881), .B(KEYINPUT44), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n913), .A2(G136), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(G162) );
  NAND2_X1 U984 ( .A1(n912), .A2(G103), .ZN(n886) );
  XOR2_X1 U985 ( .A(KEYINPUT109), .B(n886), .Z(n888) );
  NAND2_X1 U986 ( .A1(n913), .A2(G139), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U988 ( .A(KEYINPUT110), .B(n889), .ZN(n894) );
  NAND2_X1 U989 ( .A1(n908), .A2(G115), .ZN(n891) );
  NAND2_X1 U990 ( .A1(G127), .A2(n909), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n930) );
  XOR2_X1 U994 ( .A(n930), .B(G162), .Z(n897) );
  XOR2_X1 U995 ( .A(n895), .B(n944), .Z(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n902) );
  XNOR2_X1 U997 ( .A(G164), .B(n898), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U999 ( .A(n902), .B(n901), .Z(n907) );
  XOR2_X1 U1000 ( .A(KEYINPUT108), .B(KEYINPUT111), .Z(n904) );
  XNOR2_X1 U1001 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(KEYINPUT46), .B(n905), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n921) );
  NAND2_X1 U1005 ( .A1(n908), .A2(G118), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(G130), .A2(n909), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(G106), .A2(n912), .ZN(n915) );
  NAND2_X1 U1009 ( .A1(G142), .A2(n913), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1011 ( .A(KEYINPUT45), .B(n916), .Z(n917) );
  NOR2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1013 ( .A(G160), .B(n919), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n922), .ZN(G395) );
  NOR2_X1 U1016 ( .A1(G401), .A2(n929), .ZN(n926) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G397), .A2(n924), .ZN(n925) );
  NAND2_X1 U1020 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1021 ( .A1(n927), .A2(G395), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(n928), .B(KEYINPUT114), .ZN(G308) );
  INV_X1 U1023 ( .A(G308), .ZN(G225) );
  INV_X1 U1024 ( .A(n929), .ZN(G319) );
  INV_X1 U1025 ( .A(G69), .ZN(G235) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n955) );
  XOR2_X1 U1027 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n953) );
  XOR2_X1 U1028 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n933), .ZN(n938) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n936), .Z(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n949) );
  XNOR2_X1 U1036 ( .A(G160), .B(G2084), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1041 ( .A(KEYINPUT115), .B(n947), .Z(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(n953), .B(n952), .ZN(n954) );
  NAND2_X1 U1045 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1046 ( .A1(n956), .A2(G29), .ZN(n982) );
  XNOR2_X1 U1047 ( .A(G2084), .B(G34), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(n957), .B(KEYINPUT54), .ZN(n975) );
  XOR2_X1 U1049 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n958) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n958), .ZN(n970) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G32), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n965) );
  XNOR2_X1 U1054 ( .A(G2067), .B(G26), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G27), .B(n961), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1058 ( .A(G1991), .B(G25), .Z(n966) );
  NAND2_X1 U1059 ( .A1(G28), .A2(n966), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n970), .B(n969), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G35), .B(G2090), .ZN(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(n973), .B(KEYINPUT119), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(KEYINPUT55), .B(n976), .ZN(n978) );
  INV_X1 U1067 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n979), .A2(G11), .ZN(n980) );
  XOR2_X1 U1070 ( .A(KEYINPUT120), .B(n980), .Z(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n1038) );
  XNOR2_X1 U1072 ( .A(G1976), .B(G23), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G22), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1075 ( .A(KEYINPUT126), .B(n985), .Z(n987) );
  XNOR2_X1 U1076 ( .A(G1986), .B(G24), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1078 ( .A(KEYINPUT58), .B(n988), .Z(n1005) );
  XOR2_X1 U1079 ( .A(G1961), .B(G5), .Z(n1000) );
  XNOR2_X1 U1080 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n998) );
  XNOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(G4), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(G1956), .B(G20), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(G19), .B(G1341), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n996) );
  XOR2_X1 U1087 ( .A(KEYINPUT123), .B(G1981), .Z(n994) );
  XNOR2_X1 U1088 ( .A(G6), .B(n994), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(n998), .B(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G21), .B(G1966), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(KEYINPUT125), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1006), .Z(n1007) );
  NOR2_X1 U1097 ( .A1(G16), .A2(n1007), .ZN(n1035) );
  XOR2_X1 U1098 ( .A(G16), .B(KEYINPUT56), .Z(n1032) );
  XNOR2_X1 U1099 ( .A(G1956), .B(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(G1971), .A2(G303), .ZN(n1009) );
  NAND2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(n1015), .B(KEYINPUT121), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(G168), .B(G1966), .Z(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT57), .B(n1018), .Z(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(G1341), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(G301), .B(G1961), .ZN(n1026) );
  XNOR2_X1 U1112 ( .A(n1024), .B(G1348), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1117 ( .A(n1033), .B(KEYINPUT122), .ZN(n1034) );
  NOR2_X1 U1118 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1119 ( .A(n1036), .B(KEYINPUT127), .ZN(n1037) );
  NOR2_X1 U1120 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1039), .ZN(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

