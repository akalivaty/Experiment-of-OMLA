//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n445, new_n449, new_n451, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  INV_X1    g025(.A(G567), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI21_X1  g035(.A(KEYINPUT69), .B1(new_n456), .B2(G2106), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n456), .A2(KEYINPUT69), .A3(G2106), .ZN(new_n462));
  AOI211_X1 g037(.A(new_n461), .B(new_n462), .C1(G567), .C2(new_n458), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT70), .ZN(G319));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(KEYINPUT71), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n476), .A3(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n477), .A2(G137), .A3(new_n478), .A4(new_n467), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT71), .B(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n473), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  INV_X1    g059(.A(KEYINPUT72), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n477), .A2(new_n467), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(new_n478), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n477), .A2(KEYINPUT72), .A3(G2105), .A4(new_n467), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n486), .A2(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n478), .A2(G112), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n491), .A2(G136), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  AND2_X1   g072(.A1(new_n478), .A2(G138), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n477), .A2(new_n467), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(new_n478), .A3(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n470), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n477), .A2(G126), .A3(G2105), .A4(new_n467), .ZN(new_n506));
  OR2_X1    g081(.A1(G102), .A2(G2105), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n507), .B(G2104), .C1(G114), .C2(new_n478), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n517), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n524), .A2(KEYINPUT73), .A3(G50), .ZN(new_n525));
  AOI21_X1  g100(.A(KEYINPUT73), .B1(new_n524), .B2(G50), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n515), .B1(new_n516), .B2(new_n521), .C1(new_n525), .C2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT6), .B(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n519), .A2(new_n520), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n534), .A2(new_n538), .ZN(G168));
  XOR2_X1   g114(.A(KEYINPUT74), .B(G52), .Z(new_n540));
  NAND2_X1  g115(.A1(new_n524), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n542), .B2(new_n521), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n514), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n514), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT75), .B(G81), .Z(new_n550));
  OAI22_X1  g125(.A1(new_n532), .A2(new_n549), .B1(new_n521), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT76), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n532), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n532), .B2(new_n559), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n521), .A2(KEYINPUT77), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n512), .A2(new_n531), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(G91), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n514), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n562), .A2(new_n566), .A3(new_n568), .ZN(G299));
  INV_X1    g144(.A(new_n545), .ZN(new_n570));
  INV_X1    g145(.A(new_n521), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G90), .B1(new_n524), .B2(new_n540), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n570), .A2(KEYINPUT78), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT78), .B1(new_n570), .B2(new_n572), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n514), .B1(new_n535), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(G49), .B2(new_n524), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n563), .A2(G87), .A3(new_n565), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n583), .A2(new_n514), .B1(new_n584), .B2(new_n532), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n563), .A2(G86), .A3(new_n565), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT79), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n563), .A2(new_n588), .A3(G86), .A4(new_n565), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n585), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT80), .ZN(G305));
  AOI22_X1  g166(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n514), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT81), .B(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n532), .A2(new_n594), .B1(new_n521), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND3_X1  g173(.A1(new_n563), .A2(G92), .A3(new_n565), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n535), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n524), .B2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n575), .ZN(G284));
  AOI21_X1  g183(.A(new_n607), .B1(G868), .B2(new_n575), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n562), .A2(new_n566), .A3(new_n568), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  INV_X1    g191(.A(new_n552), .ZN(new_n617));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n606), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g197(.A1(new_n481), .A2(new_n467), .A3(new_n469), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n489), .A2(G123), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n478), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n491), .A2(G135), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g206(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2096), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n626), .A2(new_n634), .A3(new_n635), .ZN(G156));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  OAI21_X1  g223(.A(G14), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NOR2_X1   g228(.A1(G2072), .A2(G2078), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n442), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(KEYINPUT83), .ZN(new_n658));
  INV_X1    g233(.A(new_n655), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n655), .B(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n652), .A3(new_n658), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g243(.A1(new_n657), .A2(new_n663), .A3(new_n664), .A4(new_n666), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G1986), .ZN(new_n673));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n679), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n675), .A2(new_n678), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G1981), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(G1981), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n673), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n690), .A2(new_n686), .A3(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT85), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n689), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n689), .B2(new_n691), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n672), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n689), .A2(new_n691), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(new_n693), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n689), .A2(new_n691), .A3(new_n694), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n699), .A2(new_n700), .A3(new_n671), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(new_n701), .ZN(G229));
  NAND2_X1  g277(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n703));
  OR2_X1    g278(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G23), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT86), .Z(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(G288), .B2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT33), .B(G1976), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n707), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G1971), .ZN(new_n713));
  INV_X1    g288(.A(G1971), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n714), .B(new_n711), .C1(G166), .C2(new_n707), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n710), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n717), .B2(new_n716), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT80), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n590), .B(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(new_n707), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G6), .B2(new_n707), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT32), .B(G1981), .Z(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n719), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G25), .A2(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n489), .A2(G119), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n478), .A2(G107), .ZN(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n491), .A2(G131), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n730), .B1(new_n737), .B2(G29), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n738), .A2(new_n740), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n707), .A2(G24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n597), .B2(new_n707), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1986), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n741), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n727), .B2(KEYINPUT34), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n703), .B(new_n704), .C1(new_n729), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n632), .A2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT95), .Z(new_n750));
  NOR2_X1   g325(.A1(G168), .A2(new_n707), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n707), .B2(G21), .ZN(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT97), .Z(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT96), .B(G28), .Z(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n757), .B2(KEYINPUT30), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(KEYINPUT30), .B2(new_n757), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n759), .C1(new_n752), .C2(new_n753), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n707), .A2(G5), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G171), .B2(new_n707), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT98), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n760), .B1(new_n763), .B2(G1961), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n750), .A2(new_n755), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT99), .ZN(new_n766));
  NOR2_X1   g341(.A1(G4), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n614), .B2(G16), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(G1348), .ZN(new_n769));
  NAND2_X1  g344(.A1(G162), .A2(G29), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G29), .B2(G35), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT29), .B(G2090), .Z(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G34), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n774), .B2(KEYINPUT24), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(KEYINPUT24), .B2(new_n774), .ZN(new_n776));
  INV_X1    g351(.A(G29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n483), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT100), .Z(new_n781));
  XOR2_X1   g356(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n707), .A2(G20), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n611), .B2(new_n707), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1956), .Z(new_n786));
  AND4_X1   g361(.A1(new_n769), .A2(new_n773), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n707), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n552), .B2(new_n707), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1341), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  NOR2_X1   g366(.A1(G27), .A2(G29), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G164), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n790), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n763), .A2(G1961), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G2078), .B2(new_n793), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n778), .A2(new_n779), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT91), .Z(new_n799));
  INV_X1    g374(.A(G2067), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n777), .A2(G26), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT28), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n489), .A2(G128), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n478), .A2(G116), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n491), .A2(G140), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n802), .B1(new_n808), .B2(G29), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n799), .B1(new_n800), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n787), .A2(new_n795), .A3(new_n797), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n491), .A2(G139), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT89), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(G115), .A2(G2104), .ZN(new_n815));
  INV_X1    g390(.A(G127), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n470), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n818));
  NAND2_X1  g393(.A1(G103), .A2(G2104), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(G2105), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n478), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n817), .A2(G2105), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n814), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G29), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n777), .A2(G33), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n826), .A2(KEYINPUT90), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(KEYINPUT90), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n827), .A2(new_n828), .A3(G2072), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n777), .A2(G32), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n487), .A2(G129), .A3(new_n488), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT92), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n491), .A2(G141), .B1(G105), .B2(new_n481), .ZN(new_n833));
  NAND3_X1  g408(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT93), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT26), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n830), .B1(new_n839), .B2(new_n777), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT27), .B(G1996), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT94), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(G2072), .B1(new_n827), .B2(new_n828), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n829), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n768), .A2(G1348), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n809), .A2(new_n800), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n771), .A2(new_n772), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n848), .B(new_n849), .C1(new_n842), .C2(new_n840), .ZN(new_n850));
  NOR4_X1   g425(.A1(new_n766), .A2(new_n811), .A3(new_n845), .A4(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n852));
  INV_X1    g427(.A(new_n703), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n852), .A2(new_n728), .A3(new_n746), .A4(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n748), .A2(new_n851), .A3(new_n854), .ZN(G311));
  NAND3_X1  g430(.A1(new_n748), .A2(new_n851), .A3(new_n854), .ZN(G150));
  AOI22_X1  g431(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(new_n514), .ZN(new_n858));
  INV_X1    g433(.A(G55), .ZN(new_n859));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n532), .A2(new_n859), .B1(new_n521), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g442(.A(KEYINPUT103), .B(new_n858), .C1(new_n863), .C2(new_n864), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n552), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n617), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n614), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  AOI21_X1  g450(.A(G860), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n875), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n865), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(G145));
  NAND2_X1  g455(.A1(new_n489), .A2(G130), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n491), .A2(G142), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n478), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n624), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n838), .A2(new_n823), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n838), .A2(new_n823), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n886), .B1(new_n892), .B2(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n808), .A2(new_n510), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n803), .A2(G164), .A3(new_n807), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n895), .A2(new_n736), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n736), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n891), .A2(new_n893), .A3(new_n899), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n483), .B(KEYINPUT104), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n496), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n633), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n906), .A3(new_n902), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g487(.A1(G305), .A2(G290), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n721), .A2(new_n597), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G288), .B(KEYINPUT106), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(G303), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n916), .B(G166), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n913), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n871), .B1(G559), .B2(new_n606), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n869), .A2(new_n620), .A3(new_n870), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n614), .A2(new_n611), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n606), .A2(G299), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n606), .A2(G299), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n611), .B1(new_n601), .B2(new_n605), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT41), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n934), .A3(KEYINPUT105), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n929), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n927), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n936), .B1(new_n925), .B2(new_n926), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n922), .B(new_n924), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n922), .A2(new_n924), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n939), .B2(new_n927), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(G868), .ZN(new_n947));
  INV_X1    g522(.A(new_n865), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(G868), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(G295));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n952), .A3(new_n950), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n618), .B1(new_n942), .B2(new_n945), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT107), .B1(new_n954), .B2(new_n949), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(G331));
  OAI21_X1  g531(.A(G168), .B1(new_n573), .B2(new_n574), .ZN(new_n957));
  INV_X1    g532(.A(G171), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(G286), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n869), .A2(new_n960), .A3(new_n870), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n960), .B1(new_n870), .B2(new_n869), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n936), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n931), .A2(new_n934), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n963), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n936), .A2(KEYINPUT108), .A3(new_n929), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n968), .A2(new_n961), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n964), .A2(new_n965), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n921), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n920), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n919), .B1(new_n914), .B2(new_n913), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n935), .A2(new_n938), .A3(new_n961), .A4(new_n969), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n964), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n974), .A2(KEYINPUT43), .A3(new_n910), .A4(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n910), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n978), .B2(new_n964), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n974), .A2(new_n981), .A3(new_n910), .A4(new_n979), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT43), .B1(new_n982), .B2(new_n983), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n986), .A2(new_n991), .ZN(G397));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n503), .B1(new_n499), .B2(KEYINPUT4), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n506), .A2(new_n508), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT110), .B(G40), .Z(new_n999));
  NAND4_X1  g574(.A1(new_n473), .A2(new_n479), .A3(new_n482), .A4(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n808), .B(new_n800), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n736), .B(new_n739), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n839), .A2(G1996), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n838), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1002), .B(new_n1003), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n597), .B(new_n673), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1001), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1981), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G73), .A2(G543), .ZN(new_n1011));
  INV_X1    g586(.A(G61), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n535), .B2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1013), .A2(G651), .B1(new_n524), .B2(G48), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n571), .A2(G86), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1010), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT114), .B(G1981), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n590), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT49), .B1(new_n1019), .B2(KEYINPUT115), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n585), .B(new_n1017), .C1(new_n587), .C2(new_n589), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1021), .B(new_n1022), .C1(new_n1023), .C2(new_n1016), .ZN(new_n1024));
  OAI21_X1  g599(.A(G8), .B1(new_n996), .B2(new_n1000), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1020), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1976), .B1(new_n580), .B2(new_n581), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(G8), .C1(new_n996), .C2(new_n1000), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n1032));
  INV_X1    g607(.A(G1976), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(G288), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1025), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1029), .B(new_n1030), .C1(new_n1025), .C2(new_n1034), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1027), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT118), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1027), .A2(new_n1041), .A3(new_n1038), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n997), .A2(G1384), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n994), .B2(new_n995), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1000), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT111), .B(new_n1044), .C1(new_n994), .C2(new_n995), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n998), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n714), .ZN(new_n1051));
  INV_X1    g626(.A(G2090), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1000), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(new_n993), .C1(new_n994), .C2(new_n995), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1052), .B(new_n1053), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1051), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1051), .A2(new_n1059), .A3(KEYINPUT117), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G303), .A2(G8), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT55), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1053), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1051), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT112), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1066), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1051), .A2(new_n1072), .A3(new_n1068), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1070), .A2(new_n1071), .A3(G8), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1053), .A2(new_n779), .A3(new_n1055), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1000), .B1(new_n510), .B2(new_n1044), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1966), .B1(new_n1077), .B2(new_n998), .ZN(new_n1078));
  OAI21_X1  g653(.A(G8), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(G286), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1043), .A2(new_n1067), .A3(new_n1074), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT63), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR4_X1   g658(.A1(new_n1039), .A2(new_n1082), .A3(G286), .A4(new_n1079), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1070), .A2(G8), .A3(new_n1073), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1066), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1074), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(G288), .A2(G1976), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1023), .B1(new_n1027), .B2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1074), .A2(new_n1039), .B1(new_n1090), .B2(new_n1025), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G168), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(KEYINPUT51), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1079), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT45), .B1(new_n510), .B2(new_n993), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1048), .A2(new_n1045), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n753), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1092), .B1(new_n1098), .B2(new_n1075), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1093), .B(KEYINPUT123), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT51), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1092), .B(G168), .C1(new_n1098), .C2(new_n1075), .ZN(new_n1102));
  OAI211_X1 g677(.A(KEYINPUT62), .B(new_n1095), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1046), .A2(new_n1045), .B1(new_n996), .B2(new_n997), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1104), .A2(new_n791), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  INV_X1    g681(.A(G1961), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1105), .A2(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1077), .A2(KEYINPUT53), .A3(new_n791), .A4(new_n998), .ZN(new_n1110));
  AOI21_X1  g685(.A(G301), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1103), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(G8), .B(G286), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(KEYINPUT51), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT62), .B1(new_n1114), .B2(new_n1095), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1027), .A2(new_n1041), .A3(new_n1038), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1041), .B1(new_n1027), .B2(new_n1038), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1074), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1092), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1071), .B1(new_n1120), .B2(new_n1063), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1091), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1088), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n998), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1126));
  NAND2_X1  g701(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n791), .A2(KEYINPUT124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n791), .A2(KEYINPUT124), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(G160), .A3(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1109), .A2(G301), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1125), .B1(new_n1132), .B2(new_n1111), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1106), .B1(new_n1050), .B2(G2078), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1108), .A2(new_n1107), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(new_n1110), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT54), .B1(new_n1136), .B2(new_n575), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n958), .B1(new_n1109), .B2(new_n1131), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1114), .A2(new_n1095), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1122), .A2(new_n1133), .A3(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(G299), .B(KEYINPUT57), .ZN(new_n1143));
  AOI21_X1  g718(.A(G1384), .B1(new_n505), .B2(new_n509), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(KEYINPUT116), .A3(new_n1054), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(G1956), .B1(new_n1147), .B2(new_n1053), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT56), .B(G2072), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1050), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1143), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1126), .A2(new_n1048), .A3(new_n1149), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1143), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1053), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1153), .B(new_n1154), .C1(new_n1156), .C2(G1956), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(G1348), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n996), .A2(new_n1000), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1108), .A2(new_n1159), .B1(new_n800), .B2(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1161), .A2(new_n606), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1152), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1126), .A2(new_n1164), .A3(new_n1005), .A4(new_n1048), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT119), .B1(new_n1050), .B2(G1996), .ZN(new_n1166));
  XOR2_X1   g741(.A(KEYINPUT58), .B(G1341), .Z(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n996), .B2(new_n1000), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1165), .A2(new_n1166), .A3(new_n1170), .ZN(new_n1171));
  AND2_X1   g746(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1171), .A2(new_n552), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1161), .A2(KEYINPUT60), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1108), .A2(new_n1159), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1160), .A2(new_n800), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1175), .A2(KEYINPUT60), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n614), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1161), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1174), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n1171), .B2(new_n552), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1173), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1157), .A2(new_n1152), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1152), .A2(KEYINPUT122), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(new_n1185), .A3(KEYINPUT61), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1157), .B(new_n1152), .C1(KEYINPUT122), .C2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1163), .B1(new_n1183), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1142), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1009), .B1(new_n1124), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1001), .A2(new_n673), .A3(new_n597), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT48), .Z(new_n1194));
  AOI21_X1  g769(.A(new_n1194), .B1(new_n1007), .B2(new_n1001), .ZN(new_n1195));
  AOI21_X1  g770(.A(KEYINPUT46), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT125), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1005), .A2(KEYINPUT46), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n839), .A2(new_n1002), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1197), .B1(new_n1199), .B2(new_n1001), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT47), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1002), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n737), .A2(new_n739), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1202), .A2(new_n1203), .B1(G2067), .B2(new_n808), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n1195), .B(new_n1201), .C1(new_n1001), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1192), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g781(.A1(new_n463), .A2(new_n669), .A3(new_n668), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1208), .A2(KEYINPUT126), .ZN(new_n1209));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n1210));
  NAND4_X1  g784(.A1(new_n463), .A2(new_n668), .A3(new_n1210), .A4(new_n669), .ZN(new_n1211));
  AOI21_X1  g785(.A(G401), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n697), .A2(new_n701), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n1213), .A2(KEYINPUT127), .ZN(new_n1214));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n1215));
  NAND4_X1  g789(.A1(new_n697), .A2(new_n701), .A3(new_n1215), .A4(new_n1212), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  AND3_X1   g791(.A1(new_n1217), .A2(new_n989), .A3(new_n911), .ZN(G308));
  NAND3_X1  g792(.A1(new_n1217), .A2(new_n989), .A3(new_n911), .ZN(G225));
endmodule


