

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U561 ( .A1(n653), .A2(n550), .ZN(n547) );
  AND2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n911) );
  INV_X1 U563 ( .A(n994), .ZN(n726) );
  XNOR2_X1 U564 ( .A(n539), .B(KEYINPUT65), .ZN(G160) );
  AND2_X2 U565 ( .A1(n533), .A2(G2105), .ZN(n910) );
  OR2_X1 U566 ( .A1(n744), .A2(n743), .ZN(n797) );
  INV_X1 U567 ( .A(KEYINPUT17), .ZN(n529) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  AND2_X1 U569 ( .A1(n541), .A2(n540), .ZN(n528) );
  INV_X1 U570 ( .A(KEYINPUT104), .ZN(n715) );
  XNOR2_X1 U571 ( .A(KEYINPUT30), .B(KEYINPUT106), .ZN(n746) );
  XNOR2_X1 U572 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U573 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U574 ( .A1(G1966), .A2(n797), .ZN(n769) );
  INV_X1 U575 ( .A(n993), .ZN(n776) );
  AND2_X1 U576 ( .A1(n778), .A2(n777), .ZN(n779) );
  OR2_X1 U577 ( .A1(KEYINPUT33), .A2(n780), .ZN(n787) );
  INV_X1 U578 ( .A(G1384), .ZN(n706) );
  INV_X1 U579 ( .A(G164), .ZN(n707) );
  NAND2_X1 U580 ( .A1(n665), .A2(G66), .ZN(n605) );
  NAND2_X1 U581 ( .A1(n907), .A2(G137), .ZN(n532) );
  INV_X1 U582 ( .A(KEYINPUT1), .ZN(n551) );
  NOR2_X1 U583 ( .A1(G651), .A2(n653), .ZN(n664) );
  NOR2_X1 U584 ( .A1(G543), .A2(G651), .ZN(n663) );
  AND2_X1 U585 ( .A1(n546), .A2(n545), .ZN(G164) );
  INV_X1 U586 ( .A(G2104), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G113), .A2(n911), .ZN(n538) );
  XNOR2_X2 U588 ( .A(n530), .B(n529), .ZN(n907) );
  NAND2_X1 U589 ( .A1(G125), .A2(n910), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n536) );
  NOR2_X1 U591 ( .A1(n533), .A2(G2105), .ZN(n636) );
  NAND2_X1 U592 ( .A1(G101), .A2(n636), .ZN(n534) );
  XNOR2_X1 U593 ( .A(KEYINPUT23), .B(n534), .ZN(n535) );
  NOR2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n907), .A2(G138), .ZN(n546) );
  NAND2_X1 U597 ( .A1(G126), .A2(n910), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G114), .A2(n911), .ZN(n540) );
  AND2_X1 U599 ( .A1(n636), .A2(G102), .ZN(n543) );
  INV_X1 U600 ( .A(KEYINPUT96), .ZN(n542) );
  XNOR2_X1 U601 ( .A(n543), .B(n542), .ZN(n544) );
  AND2_X1 U602 ( .A1(n528), .A2(n544), .ZN(n545) );
  XOR2_X1 U603 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  NAND2_X1 U604 ( .A1(n664), .A2(G47), .ZN(n549) );
  XOR2_X1 U605 ( .A(KEYINPUT66), .B(G651), .Z(n550) );
  NAND2_X1 U606 ( .A1(G72), .A2(n547), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n556) );
  NAND2_X1 U608 ( .A1(n663), .A2(G85), .ZN(n554) );
  NOR2_X1 U609 ( .A1(G543), .A2(n550), .ZN(n552) );
  XNOR2_X2 U610 ( .A(n552), .B(n551), .ZN(n665) );
  NAND2_X1 U611 ( .A1(G60), .A2(n665), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U613 ( .A1(n556), .A2(n555), .ZN(G290) );
  XOR2_X1 U614 ( .A(G2446), .B(KEYINPUT114), .Z(n558) );
  XNOR2_X1 U615 ( .A(G2451), .B(G2430), .ZN(n557) );
  XNOR2_X1 U616 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U617 ( .A(n559), .B(G2427), .Z(n561) );
  XNOR2_X1 U618 ( .A(G1341), .B(G1348), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n561), .B(n560), .ZN(n565) );
  XOR2_X1 U620 ( .A(G2443), .B(G2435), .Z(n563) );
  XNOR2_X1 U621 ( .A(G2438), .B(G2454), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U623 ( .A(n565), .B(n564), .Z(n566) );
  AND2_X1 U624 ( .A1(G14), .A2(n566), .ZN(G401) );
  INV_X1 U625 ( .A(G108), .ZN(G238) );
  INV_X1 U626 ( .A(G120), .ZN(G236) );
  INV_X1 U627 ( .A(G57), .ZN(G237) );
  INV_X1 U628 ( .A(G82), .ZN(G220) );
  NAND2_X1 U629 ( .A1(G52), .A2(n664), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G64), .A2(n665), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n663), .A2(G90), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT67), .B(n569), .Z(n571) );
  NAND2_X1 U634 ( .A1(G77), .A2(n547), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n572), .Z(n573) );
  NOR2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT68), .B(n575), .Z(G301) );
  INV_X1 U639 ( .A(G301), .ZN(G171) );
  NAND2_X1 U640 ( .A1(G89), .A2(n663), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT4), .B(n576), .Z(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT79), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G76), .A2(n547), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT5), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n664), .A2(G51), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT80), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G63), .A2(n665), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U650 ( .A(KEYINPUT6), .B(n584), .Z(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U653 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U654 ( .A1(G94), .A2(G452), .ZN(n588) );
  XNOR2_X1 U655 ( .A(n588), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n589) );
  XOR2_X1 U657 ( .A(n589), .B(KEYINPUT10), .Z(n855) );
  INV_X1 U658 ( .A(n855), .ZN(G223) );
  INV_X1 U659 ( .A(G567), .ZN(n699) );
  NOR2_X1 U660 ( .A1(n699), .A2(G223), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U662 ( .A1(n664), .A2(G43), .ZN(n601) );
  NAND2_X1 U663 ( .A1(n663), .A2(G81), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT12), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G68), .A2(n547), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U667 ( .A(KEYINPUT13), .B(n594), .ZN(n598) );
  XOR2_X1 U668 ( .A(KEYINPUT14), .B(KEYINPUT73), .Z(n596) );
  NAND2_X1 U669 ( .A1(G56), .A2(n665), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n596), .B(n595), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U672 ( .A(KEYINPUT74), .B(n599), .Z(n600) );
  AND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n1001) );
  NAND2_X1 U674 ( .A1(G860), .A2(n1001), .ZN(n602) );
  XOR2_X1 U675 ( .A(KEYINPUT75), .B(n602), .Z(G153) );
  NAND2_X1 U676 ( .A1(n664), .A2(G54), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G79), .A2(n547), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n663), .A2(G92), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X2 U682 ( .A(KEYINPUT15), .B(n609), .Z(n610) );
  XOR2_X2 U683 ( .A(KEYINPUT77), .B(n610), .Z(n994) );
  INV_X1 U684 ( .A(G868), .ZN(n684) );
  NAND2_X1 U685 ( .A1(n726), .A2(n684), .ZN(n611) );
  XNOR2_X1 U686 ( .A(KEYINPUT78), .B(n611), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G301), .A2(G868), .ZN(n612) );
  XNOR2_X1 U688 ( .A(KEYINPUT76), .B(n612), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(G284) );
  NAND2_X1 U690 ( .A1(G53), .A2(n664), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G65), .A2(n665), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U693 ( .A(KEYINPUT71), .B(n617), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n663), .A2(G91), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G78), .A2(n547), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U697 ( .A(KEYINPUT70), .B(n620), .Z(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(G299) );
  NOR2_X1 U699 ( .A1(G286), .A2(n684), .ZN(n624) );
  NOR2_X1 U700 ( .A1(G868), .A2(G299), .ZN(n623) );
  NOR2_X1 U701 ( .A1(n624), .A2(n623), .ZN(G297) );
  INV_X1 U702 ( .A(G860), .ZN(n861) );
  NAND2_X1 U703 ( .A1(n861), .A2(G559), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n625), .A2(n994), .ZN(n626) );
  XNOR2_X1 U705 ( .A(n626), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U706 ( .A1(n1001), .A2(n684), .ZN(n627) );
  XNOR2_X1 U707 ( .A(KEYINPUT81), .B(n627), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G868), .A2(n994), .ZN(n628) );
  NOR2_X1 U709 ( .A1(G559), .A2(n628), .ZN(n629) );
  NOR2_X1 U710 ( .A1(n630), .A2(n629), .ZN(G282) );
  XOR2_X1 U711 ( .A(G2100), .B(KEYINPUT82), .Z(n640) );
  NAND2_X1 U712 ( .A1(G135), .A2(n907), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G111), .A2(n911), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n910), .A2(G123), .ZN(n633) );
  XOR2_X1 U716 ( .A(KEYINPUT18), .B(n633), .Z(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n638) );
  BUF_X1 U718 ( .A(n636), .Z(n906) );
  NAND2_X1 U719 ( .A1(n906), .A2(G99), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n950) );
  XOR2_X1 U721 ( .A(G2096), .B(n950), .Z(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(G156) );
  XOR2_X1 U723 ( .A(KEYINPUT87), .B(KEYINPUT2), .Z(n642) );
  NAND2_X1 U724 ( .A1(G73), .A2(n547), .ZN(n641) );
  XNOR2_X1 U725 ( .A(n642), .B(n641), .ZN(n649) );
  NAND2_X1 U726 ( .A1(G48), .A2(n664), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G86), .A2(n663), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n665), .A2(G61), .ZN(n645) );
  XOR2_X1 U730 ( .A(KEYINPUT86), .B(n645), .Z(n646) );
  NOR2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U732 ( .A1(n649), .A2(n648), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G49), .A2(n664), .ZN(n651) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U736 ( .A1(n665), .A2(n652), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G87), .A2(n653), .ZN(n654) );
  XOR2_X1 U738 ( .A(KEYINPUT85), .B(n654), .Z(n655) );
  NAND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(G288) );
  NAND2_X1 U740 ( .A1(n663), .A2(G88), .ZN(n658) );
  NAND2_X1 U741 ( .A1(G75), .A2(n547), .ZN(n657) );
  NAND2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U743 ( .A1(G50), .A2(n664), .ZN(n660) );
  NAND2_X1 U744 ( .A1(G62), .A2(n665), .ZN(n659) );
  NAND2_X1 U745 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U746 ( .A1(n662), .A2(n661), .ZN(G166) );
  INV_X1 U747 ( .A(G166), .ZN(G303) );
  NAND2_X1 U748 ( .A1(G93), .A2(n663), .ZN(n672) );
  NAND2_X1 U749 ( .A1(G55), .A2(n664), .ZN(n667) );
  NAND2_X1 U750 ( .A1(G67), .A2(n665), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U752 ( .A1(G80), .A2(n547), .ZN(n668) );
  XNOR2_X1 U753 ( .A(KEYINPUT83), .B(n668), .ZN(n669) );
  NOR2_X1 U754 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U755 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U756 ( .A(n673), .B(KEYINPUT84), .ZN(n862) );
  XNOR2_X1 U757 ( .A(KEYINPUT88), .B(G305), .ZN(n674) );
  XNOR2_X1 U758 ( .A(n674), .B(G288), .ZN(n675) );
  XNOR2_X1 U759 ( .A(KEYINPUT19), .B(n675), .ZN(n677) );
  XOR2_X1 U760 ( .A(G290), .B(G303), .Z(n676) );
  XNOR2_X1 U761 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U762 ( .A(n862), .B(n678), .ZN(n679) );
  INV_X1 U763 ( .A(G299), .ZN(n731) );
  XOR2_X1 U764 ( .A(n679), .B(n731), .Z(n931) );
  NAND2_X1 U765 ( .A1(G559), .A2(n994), .ZN(n680) );
  XNOR2_X1 U766 ( .A(n680), .B(n1001), .ZN(n860) );
  XNOR2_X1 U767 ( .A(n931), .B(n860), .ZN(n681) );
  XNOR2_X1 U768 ( .A(n681), .B(KEYINPUT89), .ZN(n682) );
  NAND2_X1 U769 ( .A1(n682), .A2(G868), .ZN(n683) );
  XNOR2_X1 U770 ( .A(n683), .B(KEYINPUT90), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n862), .A2(n684), .ZN(n685) );
  NAND2_X1 U772 ( .A1(n686), .A2(n685), .ZN(G295) );
  NAND2_X1 U773 ( .A1(G2078), .A2(G2084), .ZN(n687) );
  XOR2_X1 U774 ( .A(KEYINPUT20), .B(n687), .Z(n688) );
  NAND2_X1 U775 ( .A1(G2090), .A2(n688), .ZN(n690) );
  XOR2_X1 U776 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n689) );
  XNOR2_X1 U777 ( .A(n690), .B(n689), .ZN(n691) );
  NAND2_X1 U778 ( .A1(G2072), .A2(n691), .ZN(G158) );
  XNOR2_X1 U779 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U780 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  NOR2_X1 U781 ( .A1(G219), .A2(G220), .ZN(n692) );
  XNOR2_X1 U782 ( .A(KEYINPUT22), .B(n692), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n693), .A2(G96), .ZN(n694) );
  NOR2_X1 U784 ( .A1(G218), .A2(n694), .ZN(n695) );
  XOR2_X1 U785 ( .A(KEYINPUT92), .B(n695), .Z(n865) );
  NAND2_X1 U786 ( .A1(n865), .A2(G2106), .ZN(n696) );
  XNOR2_X1 U787 ( .A(n696), .B(KEYINPUT93), .ZN(n701) );
  NOR2_X1 U788 ( .A1(G236), .A2(G238), .ZN(n697) );
  NAND2_X1 U789 ( .A1(G69), .A2(n697), .ZN(n698) );
  NOR2_X1 U790 ( .A1(G237), .A2(n698), .ZN(n864) );
  NOR2_X1 U791 ( .A1(n699), .A2(n864), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n701), .A2(n700), .ZN(G319) );
  NAND2_X1 U793 ( .A1(G483), .A2(G661), .ZN(n703) );
  INV_X1 U794 ( .A(G319), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U796 ( .A(n704), .B(KEYINPUT94), .ZN(n859) );
  NAND2_X1 U797 ( .A1(n859), .A2(G36), .ZN(n705) );
  XOR2_X1 U798 ( .A(KEYINPUT95), .B(n705), .Z(G176) );
  INV_X1 U799 ( .A(G40), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n800) );
  NOR2_X1 U801 ( .A1(n708), .A2(n800), .ZN(n709) );
  AND2_X2 U802 ( .A1(n709), .A2(G160), .ZN(n743) );
  NAND2_X1 U803 ( .A1(n743), .A2(G1996), .ZN(n710) );
  XNOR2_X1 U804 ( .A(n710), .B(KEYINPUT26), .ZN(n712) );
  INV_X1 U805 ( .A(n743), .ZN(n753) );
  NAND2_X1 U806 ( .A1(G1341), .A2(n753), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U808 ( .A(n713), .B(KEYINPUT103), .ZN(n714) );
  NAND2_X1 U809 ( .A1(n714), .A2(n1001), .ZN(n727) );
  NOR2_X1 U810 ( .A1(n727), .A2(n726), .ZN(n716) );
  XNOR2_X1 U811 ( .A(n716), .B(n715), .ZN(n724) );
  NOR2_X1 U812 ( .A1(n743), .A2(G1348), .ZN(n718) );
  NOR2_X1 U813 ( .A1(G2067), .A2(n753), .ZN(n717) );
  NOR2_X1 U814 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n743), .A2(G2072), .ZN(n719) );
  XNOR2_X1 U816 ( .A(n719), .B(KEYINPUT27), .ZN(n721) );
  XOR2_X1 U817 ( .A(G1956), .B(KEYINPUT102), .Z(n1010) );
  NOR2_X1 U818 ( .A1(n743), .A2(n1010), .ZN(n720) );
  NOR2_X1 U819 ( .A1(n721), .A2(n720), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n725) );
  AND2_X1 U821 ( .A1(n722), .A2(n725), .ZN(n723) );
  NAND2_X1 U822 ( .A1(n724), .A2(n723), .ZN(n736) );
  INV_X1 U823 ( .A(n725), .ZN(n729) );
  NAND2_X1 U824 ( .A1(n727), .A2(n726), .ZN(n728) );
  OR2_X1 U825 ( .A1(n729), .A2(n728), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U827 ( .A(n732), .B(KEYINPUT28), .Z(n733) );
  AND2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U830 ( .A(n737), .B(KEYINPUT29), .ZN(n741) );
  XNOR2_X1 U831 ( .A(G2078), .B(KEYINPUT25), .ZN(n974) );
  NOR2_X1 U832 ( .A1(n753), .A2(n974), .ZN(n739) );
  AND2_X1 U833 ( .A1(n753), .A2(G1961), .ZN(n738) );
  NOR2_X1 U834 ( .A1(n739), .A2(n738), .ZN(n749) );
  AND2_X1 U835 ( .A1(n749), .A2(G171), .ZN(n740) );
  NOR2_X1 U836 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U837 ( .A(n742), .B(KEYINPUT105), .ZN(n767) );
  INV_X1 U838 ( .A(G8), .ZN(n744) );
  NOR2_X1 U839 ( .A1(G2084), .A2(n753), .ZN(n765) );
  NOR2_X1 U840 ( .A1(n769), .A2(n765), .ZN(n745) );
  NAND2_X1 U841 ( .A1(G8), .A2(n745), .ZN(n747) );
  NOR2_X1 U842 ( .A1(G168), .A2(n748), .ZN(n751) );
  NOR2_X1 U843 ( .A1(n749), .A2(G171), .ZN(n750) );
  XOR2_X1 U844 ( .A(KEYINPUT31), .B(n752), .Z(n766) );
  NOR2_X1 U845 ( .A1(G1971), .A2(n797), .ZN(n755) );
  NOR2_X1 U846 ( .A1(G2090), .A2(n753), .ZN(n754) );
  NOR2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n756), .A2(G303), .ZN(n758) );
  AND2_X1 U849 ( .A1(n766), .A2(n758), .ZN(n757) );
  NAND2_X1 U850 ( .A1(n767), .A2(n757), .ZN(n762) );
  INV_X1 U851 ( .A(n758), .ZN(n759) );
  OR2_X1 U852 ( .A1(n759), .A2(G286), .ZN(n760) );
  AND2_X1 U853 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n764) );
  XOR2_X1 U855 ( .A(KEYINPUT32), .B(KEYINPUT107), .Z(n763) );
  XNOR2_X1 U856 ( .A(n764), .B(n763), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G8), .A2(n765), .ZN(n771) );
  AND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n788) );
  NOR2_X1 U862 ( .A1(G1976), .A2(G288), .ZN(n781) );
  NOR2_X1 U863 ( .A1(G1971), .A2(G303), .ZN(n774) );
  OR2_X1 U864 ( .A1(n781), .A2(n774), .ZN(n991) );
  XOR2_X1 U865 ( .A(KEYINPUT108), .B(n991), .Z(n775) );
  NAND2_X1 U866 ( .A1(n788), .A2(n775), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NOR2_X1 U868 ( .A1(n797), .A2(n776), .ZN(n777) );
  XNOR2_X1 U869 ( .A(n779), .B(KEYINPUT64), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(KEYINPUT33), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n782), .A2(n797), .ZN(n785) );
  XNOR2_X1 U872 ( .A(G1981), .B(KEYINPUT109), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n783), .B(G305), .ZN(n987) );
  INV_X1 U874 ( .A(n987), .ZN(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n793) );
  NOR2_X1 U877 ( .A1(G2090), .A2(G303), .ZN(n789) );
  NAND2_X1 U878 ( .A1(G8), .A2(n789), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n788), .A2(n790), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n791), .A2(n797), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U882 ( .A(n794), .B(KEYINPUT110), .ZN(n799) );
  NOR2_X1 U883 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XOR2_X1 U884 ( .A(n795), .B(KEYINPUT24), .Z(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n834) );
  INV_X1 U887 ( .A(n800), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G160), .A2(G40), .ZN(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n850) );
  NAND2_X1 U890 ( .A1(G128), .A2(n910), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G116), .A2(n911), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U893 ( .A(KEYINPUT35), .B(n805), .ZN(n811) );
  NAND2_X1 U894 ( .A1(n907), .A2(G140), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n806), .B(KEYINPUT98), .ZN(n808) );
  NAND2_X1 U896 ( .A1(G104), .A2(n906), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U898 ( .A(KEYINPUT34), .B(n809), .Z(n810) );
  NAND2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U900 ( .A(KEYINPUT36), .B(n812), .Z(n922) );
  XNOR2_X1 U901 ( .A(G2067), .B(KEYINPUT37), .ZN(n813) );
  XOR2_X1 U902 ( .A(n813), .B(KEYINPUT97), .Z(n837) );
  NOR2_X1 U903 ( .A1(n922), .A2(n837), .ZN(n961) );
  NAND2_X1 U904 ( .A1(n850), .A2(n961), .ZN(n847) );
  NAND2_X1 U905 ( .A1(n911), .A2(G107), .ZN(n816) );
  NAND2_X1 U906 ( .A1(G131), .A2(n907), .ZN(n814) );
  XOR2_X1 U907 ( .A(KEYINPUT99), .B(n814), .Z(n815) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n820) );
  NAND2_X1 U909 ( .A1(G95), .A2(n906), .ZN(n818) );
  NAND2_X1 U910 ( .A1(G119), .A2(n910), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  OR2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n925) );
  AND2_X1 U913 ( .A1(n925), .A2(G1991), .ZN(n831) );
  XOR2_X1 U914 ( .A(KEYINPUT101), .B(KEYINPUT38), .Z(n822) );
  NAND2_X1 U915 ( .A1(G105), .A2(n906), .ZN(n821) );
  XNOR2_X1 U916 ( .A(n822), .B(n821), .ZN(n829) );
  NAND2_X1 U917 ( .A1(G141), .A2(n907), .ZN(n824) );
  NAND2_X1 U918 ( .A1(G129), .A2(n910), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n911), .A2(G117), .ZN(n825) );
  XOR2_X1 U921 ( .A(KEYINPUT100), .B(n825), .Z(n826) );
  NOR2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n901) );
  AND2_X1 U924 ( .A1(n901), .A2(G1996), .ZN(n830) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n955) );
  INV_X1 U926 ( .A(n955), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n832), .A2(n850), .ZN(n839) );
  NAND2_X1 U928 ( .A1(n847), .A2(n839), .ZN(n833) );
  NOR2_X1 U929 ( .A1(n834), .A2(n833), .ZN(n836) );
  XNOR2_X1 U930 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U931 ( .A1(n990), .A2(n850), .ZN(n835) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(n853) );
  AND2_X1 U933 ( .A1(n837), .A2(n922), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n838), .B(KEYINPUT113), .ZN(n958) );
  NOR2_X1 U935 ( .A1(G1996), .A2(n901), .ZN(n940) );
  INV_X1 U936 ( .A(n839), .ZN(n842) );
  NOR2_X1 U937 ( .A1(G1991), .A2(n925), .ZN(n953) );
  NOR2_X1 U938 ( .A1(G1986), .A2(G290), .ZN(n840) );
  NOR2_X1 U939 ( .A1(n953), .A2(n840), .ZN(n841) );
  NOR2_X1 U940 ( .A1(n842), .A2(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(KEYINPUT111), .B(n843), .Z(n844) );
  NOR2_X1 U942 ( .A1(n940), .A2(n844), .ZN(n845) );
  XNOR2_X1 U943 ( .A(KEYINPUT112), .B(n845), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n846), .B(KEYINPUT39), .ZN(n848) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n958), .A2(n849), .ZN(n851) );
  NAND2_X1 U947 ( .A1(n851), .A2(n850), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n854), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U950 ( .A1(G2106), .A2(n855), .ZN(G217) );
  NAND2_X1 U951 ( .A1(G15), .A2(G2), .ZN(n856) );
  XNOR2_X1 U952 ( .A(KEYINPUT115), .B(n856), .ZN(n857) );
  NAND2_X1 U953 ( .A1(n857), .A2(G661), .ZN(G259) );
  NAND2_X1 U954 ( .A1(G3), .A2(G1), .ZN(n858) );
  NAND2_X1 U955 ( .A1(n859), .A2(n858), .ZN(G188) );
  NAND2_X1 U957 ( .A1(n861), .A2(n860), .ZN(n863) );
  XNOR2_X1 U958 ( .A(n863), .B(n862), .ZN(G145) );
  INV_X1 U959 ( .A(G96), .ZN(G221) );
  INV_X1 U960 ( .A(n864), .ZN(n866) );
  NOR2_X1 U961 ( .A1(n866), .A2(n865), .ZN(G325) );
  INV_X1 U962 ( .A(G325), .ZN(G261) );
  XOR2_X1 U963 ( .A(G2096), .B(G2100), .Z(n868) );
  XNOR2_X1 U964 ( .A(KEYINPUT42), .B(G2678), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U966 ( .A(KEYINPUT43), .B(G2090), .Z(n870) );
  XNOR2_X1 U967 ( .A(G2067), .B(G2072), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U969 ( .A(n872), .B(n871), .Z(n874) );
  XNOR2_X1 U970 ( .A(G2078), .B(G2084), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(G227) );
  XOR2_X1 U972 ( .A(G2474), .B(G1956), .Z(n876) );
  XNOR2_X1 U973 ( .A(G1986), .B(G1961), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U975 ( .A(n877), .B(KEYINPUT41), .Z(n879) );
  XNOR2_X1 U976 ( .A(G1996), .B(G1991), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n883) );
  XOR2_X1 U978 ( .A(G1971), .B(G1966), .Z(n881) );
  XNOR2_X1 U979 ( .A(G1981), .B(G1976), .ZN(n880) );
  XNOR2_X1 U980 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U981 ( .A(n883), .B(n882), .Z(n885) );
  XNOR2_X1 U982 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(G229) );
  NAND2_X1 U984 ( .A1(G124), .A2(n910), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n886), .B(KEYINPUT44), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n887), .B(KEYINPUT118), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G112), .A2(n911), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n893) );
  NAND2_X1 U989 ( .A1(G100), .A2(n906), .ZN(n891) );
  NAND2_X1 U990 ( .A1(G136), .A2(n907), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n892) );
  NOR2_X1 U992 ( .A1(n893), .A2(n892), .ZN(G162) );
  NAND2_X1 U993 ( .A1(G130), .A2(n910), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G118), .A2(n911), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n900) );
  NAND2_X1 U996 ( .A1(G106), .A2(n906), .ZN(n897) );
  NAND2_X1 U997 ( .A1(G142), .A2(n907), .ZN(n896) );
  NAND2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U999 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n921) );
  XOR2_X1 U1002 ( .A(KEYINPUT46), .B(KEYINPUT120), .Z(n904) );
  XNOR2_X1 U1003 ( .A(KEYINPUT121), .B(KEYINPUT48), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n950), .B(n905), .ZN(n919) );
  NAND2_X1 U1006 ( .A1(G103), .A2(n906), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(G139), .A2(n907), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n917) );
  NAND2_X1 U1009 ( .A1(G127), .A2(n910), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(G115), .A2(n911), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT119), .B(n914), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT47), .B(n915), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n942) );
  XNOR2_X1 U1015 ( .A(G164), .B(n942), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1017 ( .A(n921), .B(n920), .Z(n924) );
  XOR2_X1 U1018 ( .A(n922), .B(G162), .Z(n923) );
  XNOR2_X1 U1019 ( .A(n924), .B(n923), .ZN(n927) );
  XOR2_X1 U1020 ( .A(n925), .B(G160), .Z(n926) );
  XNOR2_X1 U1021 ( .A(n927), .B(n926), .ZN(n928) );
  NOR2_X1 U1022 ( .A1(G37), .A2(n928), .ZN(G395) );
  XOR2_X1 U1023 ( .A(G286), .B(n1001), .Z(n930) );
  XOR2_X1 U1024 ( .A(G171), .B(n994), .Z(n929) );
  XNOR2_X1 U1025 ( .A(n930), .B(n929), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(n932), .B(n931), .ZN(n933) );
  NOR2_X1 U1027 ( .A1(G37), .A2(n933), .ZN(G397) );
  NOR2_X1 U1028 ( .A1(G227), .A2(G229), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(KEYINPUT49), .B(n934), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(G401), .A2(n935), .ZN(n936) );
  AND2_X1 U1031 ( .A1(G319), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(G395), .A2(G397), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(G225) );
  INV_X1 U1034 ( .A(G225), .ZN(G308) );
  INV_X1 U1035 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1038 ( .A(KEYINPUT51), .B(n941), .Z(n948) );
  XNOR2_X1 U1039 ( .A(KEYINPUT123), .B(KEYINPUT50), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G2072), .B(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G164), .B(G2078), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n946), .B(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n957) );
  XNOR2_X1 U1045 ( .A(G160), .B(G2084), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(n949), .B(KEYINPUT122), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(KEYINPUT52), .B(n962), .ZN(n964) );
  INV_X1 U1054 ( .A(KEYINPUT55), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n965), .A2(G29), .ZN(n1040) );
  XNOR2_X1 U1057 ( .A(G2090), .B(G35), .ZN(n979) );
  XNOR2_X1 U1058 ( .A(G1991), .B(G25), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(G33), .B(G2072), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n973) );
  XOR2_X1 U1061 ( .A(G2067), .B(G26), .Z(n968) );
  NAND2_X1 U1062 ( .A1(n968), .A2(G28), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G32), .B(G1996), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(KEYINPUT124), .B(n969), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1067 ( .A(G27), .B(n974), .Z(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(KEYINPUT53), .B(n977), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1071 ( .A(G2084), .B(KEYINPUT54), .Z(n980) );
  XNOR2_X1 U1072 ( .A(G34), .B(n980), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1074 ( .A(KEYINPUT55), .B(n983), .Z(n985) );
  INV_X1 U1075 ( .A(G29), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(G11), .A2(n986), .ZN(n1038) );
  INV_X1 U1078 ( .A(G16), .ZN(n1034) );
  XOR2_X1 U1079 ( .A(n1034), .B(KEYINPUT56), .Z(n1009) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(KEYINPUT57), .ZN(n1007) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n1000) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(n994), .B(G1348), .ZN(n996) );
  XOR2_X1 U1087 ( .A(G299), .B(G1956), .Z(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1001), .B(G1341), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(G301), .B(G1961), .Z(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1036) );
  XOR2_X1 U1097 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n1020) );
  XOR2_X1 U1098 ( .A(G1341), .B(G19), .Z(n1012) );
  XNOR2_X1 U1099 ( .A(n1010), .B(G20), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G6), .B(G1981), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(G4), .B(KEYINPUT125), .Z(n1016) );
  XNOR2_X1 U1104 ( .A(G1348), .B(KEYINPUT59), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1016), .B(n1015), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(n1020), .B(n1019), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(G1966), .B(G21), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(G5), .B(G1961), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1031) );
  XNOR2_X1 U1112 ( .A(G1976), .B(G23), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(G1971), .B(G22), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XOR2_X1 U1115 ( .A(G1986), .B(G24), .Z(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1117 ( .A(KEYINPUT58), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1119 ( .A(KEYINPUT61), .B(n1032), .ZN(n1033) );
  NAND2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1122 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1123 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1124 ( .A(n1041), .B(KEYINPUT127), .ZN(n1042) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1042), .Z(G150) );
  INV_X1 U1126 ( .A(G150), .ZN(G311) );
endmodule

