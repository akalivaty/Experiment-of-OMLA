//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  XNOR2_X1  g000(.A(KEYINPUT88), .B(G29gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT89), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n202), .A2(KEYINPUT89), .A3(G36gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT90), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT15), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT91), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n213), .B(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n206), .A2(new_n209), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT91), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n205), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n211), .A2(new_n212), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n210), .A2(KEYINPUT15), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT92), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n221), .A2(new_n226), .A3(new_n223), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G1gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G1gat), .B2(new_n228), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(G8gat), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n225), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n221), .A2(new_n226), .A3(new_n223), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n226), .B1(new_n221), .B2(new_n223), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT17), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n221), .A2(KEYINPUT17), .A3(new_n223), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n232), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n234), .B(new_n235), .C1(new_n238), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n227), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n232), .B(new_n239), .C1(new_n244), .C2(KEYINPUT17), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n245), .A2(KEYINPUT18), .A3(new_n235), .A4(new_n234), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n235), .B(KEYINPUT13), .Z(new_n247));
  NOR2_X1   g046(.A1(new_n236), .A2(new_n237), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(new_n233), .ZN(new_n249));
  INV_X1    g048(.A(new_n234), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G197gat), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT11), .B(G169gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n258), .B(KEYINPUT12), .Z(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n259), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n252), .A2(new_n253), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT83), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT31), .B(G50gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(G228gat), .A2(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(G155gat), .ZN(new_n267));
  INV_X1    g066(.A(G162gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT78), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(KEYINPUT78), .A3(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(KEYINPUT2), .ZN(new_n275));
  INV_X1    g074(.A(G141gat), .ZN(new_n276));
  INV_X1    g075(.A(G148gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G141gat), .A2(G148gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n273), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n271), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n278), .A2(new_n279), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT78), .A4(new_n275), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n287));
  XNOR2_X1  g086(.A(G197gat), .B(G204gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT22), .ZN(new_n289));
  INV_X1    g088(.A(G211gat), .ZN(new_n290));
  INV_X1    g089(.A(G218gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT29), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n287), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n294), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n293), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT82), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n286), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n300), .B1(new_n306), .B2(new_n301), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n266), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n305), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n286), .B1(new_n296), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n308), .A2(new_n311), .A3(new_n266), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n265), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(G22gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n265), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT3), .B1(new_n302), .B2(KEYINPUT82), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n296), .A2(new_n297), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n307), .B1(new_n320), .B2(new_n286), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n312), .B(new_n317), .C1(new_n321), .C2(new_n266), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n314), .A2(new_n316), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n316), .B1(new_n314), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(G1gat), .B(G29gat), .Z(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G57gat), .B(G85gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  XOR2_X1   g130(.A(G127gat), .B(G134gat), .Z(new_n332));
  INV_X1    g131(.A(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G113gat), .ZN(new_n334));
  INV_X1    g133(.A(G113gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G120gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT71), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n337), .A2(KEYINPUT71), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n332), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n332), .A2(KEYINPUT1), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n335), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n334), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n286), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT1), .B1(new_n337), .B2(KEYINPUT71), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(KEYINPUT71), .B2(new_n337), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n352), .A2(new_n332), .B1(new_n347), .B2(new_n343), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n285), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n331), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n349), .B(new_n306), .C1(new_n287), .C2(new_n285), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n360), .B1(new_n353), .B2(new_n285), .ZN(new_n361));
  AND4_X1   g160(.A1(new_n360), .A2(new_n342), .A3(new_n285), .A4(new_n348), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n359), .B(new_n356), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT80), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n363), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n354), .A2(KEYINPUT4), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n353), .A2(new_n360), .A3(new_n285), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n369), .A2(new_n331), .A3(new_n356), .A4(new_n359), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n330), .B(new_n365), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n374));
  INV_X1    g173(.A(new_n330), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n372), .B1(new_n366), .B2(new_n370), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n364), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n373), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(KEYINPUT6), .B(new_n375), .C1(new_n376), .C2(new_n364), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT68), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT27), .B(G183gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G190gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT28), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n381), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n382), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n384), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT67), .B1(new_n388), .B2(G183gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n384), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n383), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n386), .B(new_n387), .C1(new_n392), .C2(KEYINPUT28), .ZN(new_n393));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT26), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G169gat), .ZN(new_n398));
  INV_X1    g197(.A(G176gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT69), .B1(new_n400), .B2(KEYINPUT26), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT69), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n395), .A2(new_n402), .A3(new_n396), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n397), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT70), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT70), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n404), .A2(new_n409), .A3(new_n406), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n393), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT23), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n412), .A2(G169gat), .A3(G176gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n394), .A2(KEYINPUT23), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n400), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n405), .ZN(new_n417));
  NAND3_X1  g216(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT25), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT64), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n417), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n395), .A2(KEYINPUT23), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n412), .B1(G169gat), .B2(G176gat), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT25), .B(new_n425), .C1(new_n426), .C2(new_n395), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT65), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n417), .A2(new_n421), .A3(new_n423), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n415), .A2(new_n429), .A3(new_n430), .A4(KEYINPUT25), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT66), .B(new_n420), .C1(new_n428), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT66), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n431), .ZN(new_n434));
  INV_X1    g233(.A(new_n420), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n411), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT75), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(KEYINPUT75), .B(new_n411), .C1(new_n432), .C2(new_n436), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(G226gat), .A3(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n434), .A2(new_n435), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n411), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(G226gat), .A2(G233gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n301), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n295), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n439), .A2(new_n301), .A3(new_n440), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT76), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT76), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n451), .A3(new_n445), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n445), .B1(new_n411), .B2(new_n443), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n447), .B1(new_n455), .B2(new_n295), .ZN(new_n456));
  XOR2_X1   g255(.A(G8gat), .B(G36gat), .Z(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(KEYINPUT77), .ZN(new_n458));
  XNOR2_X1  g257(.A(G64gat), .B(G92gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n380), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n455), .A2(new_n295), .ZN(new_n465));
  INV_X1    g264(.A(new_n447), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n465), .A2(KEYINPUT30), .A3(new_n466), .A4(new_n461), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n453), .B1(new_n449), .B2(KEYINPUT76), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n300), .B1(new_n468), .B2(new_n452), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n460), .B1(new_n469), .B2(new_n447), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n325), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT74), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n437), .A2(new_n353), .ZN(new_n474));
  INV_X1    g273(.A(G227gat), .ZN(new_n475));
  INV_X1    g274(.A(G233gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n349), .B(new_n411), .C1(new_n432), .C2(new_n436), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT32), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT33), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G71gat), .B(G99gat), .Z(new_n483));
  XNOR2_X1  g282(.A(G15gat), .B(G43gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n480), .B1(new_n485), .B2(KEYINPUT33), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n479), .A2(KEYINPUT73), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT73), .B1(new_n479), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n478), .ZN(new_n492));
  INV_X1    g291(.A(new_n477), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI211_X1 g293(.A(KEYINPUT34), .B(new_n477), .C1(new_n474), .C2(new_n478), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n494), .A2(new_n495), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n487), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT73), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n479), .A2(KEYINPUT73), .A3(new_n487), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n498), .B1(new_n503), .B2(new_n486), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n473), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n496), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n498), .B(new_n486), .C1(new_n489), .C2(new_n488), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n473), .A3(KEYINPUT36), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n264), .B1(new_n472), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n325), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n378), .A2(new_n379), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n469), .A2(new_n447), .A3(new_n460), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(KEYINPUT30), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n467), .A2(new_n470), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT83), .A3(new_n511), .A4(new_n507), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT40), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n356), .B1(new_n369), .B2(new_n359), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n522), .A2(KEYINPUT84), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n369), .A2(new_n359), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(KEYINPUT84), .A3(new_n357), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n350), .A2(new_n354), .A3(new_n356), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n523), .A2(KEYINPUT39), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n330), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT39), .B1(new_n523), .B2(new_n525), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n529), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n531), .A2(KEYINPUT40), .A3(new_n330), .A4(new_n527), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n530), .A2(new_n377), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT30), .B1(new_n456), .B2(new_n461), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n518), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT38), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n461), .B1(new_n456), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT37), .B1(new_n469), .B2(new_n447), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n515), .B1(new_n456), .B2(new_n461), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n448), .A2(new_n451), .A3(new_n445), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n451), .B1(new_n448), .B2(new_n445), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n542), .A2(new_n543), .A3(new_n453), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n537), .B(new_n466), .C1(new_n544), .C2(new_n300), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n442), .A2(new_n446), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n537), .B1(new_n546), .B2(new_n295), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n544), .B2(new_n295), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n545), .A2(new_n548), .A3(new_n536), .A4(new_n460), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n541), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n535), .B(new_n325), .C1(new_n540), .C2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n513), .A2(new_n520), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n508), .A2(new_n509), .A3(new_n325), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT86), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n508), .A2(new_n509), .A3(new_n325), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n534), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n557), .A2(new_n471), .A3(new_n515), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT35), .ZN(new_n560));
  INV_X1    g359(.A(new_n553), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT85), .B(KEYINPUT35), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n464), .A2(new_n471), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n263), .B1(new_n552), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n239), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n567));
  NAND3_X1  g366(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(KEYINPUT7), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(KEYINPUT8), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n572), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G99gat), .B(G106gat), .Z(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(KEYINPUT99), .A3(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT99), .B1(new_n579), .B2(new_n580), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n567), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(new_n581), .A3(KEYINPUT100), .A4(new_n582), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OR3_X1    g387(.A1(new_n238), .A2(new_n566), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G232gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(new_n476), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n248), .A2(new_n588), .B1(KEYINPUT41), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n595), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n599), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n593), .A2(new_n597), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n603), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n604), .B1(new_n593), .B2(new_n597), .ZN(new_n608));
  AOI211_X1 g407(.A(new_n596), .B(new_n599), .C1(new_n589), .C2(new_n592), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G57gat), .B(G64gat), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n613), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G71gat), .B(G78gat), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n618), .A2(KEYINPUT93), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(KEYINPUT93), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT95), .ZN(new_n622));
  INV_X1    g421(.A(new_n617), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n618), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n617), .A2(new_n619), .A3(new_n625), .A4(new_n620), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n622), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G127gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n232), .B1(new_n627), .B2(new_n628), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT96), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n634), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(new_n267), .ZN(new_n638));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  AND3_X1   g439(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n635), .B2(new_n636), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n611), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(KEYINPUT103), .Z(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n580), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n579), .B(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n650), .A2(new_n626), .A3(new_n624), .A4(new_n622), .ZN(new_n651));
  INV_X1    g450(.A(new_n627), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n583), .A2(new_n584), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n647), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n585), .A2(new_n652), .A3(KEYINPUT10), .A4(new_n587), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n646), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n646), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n659), .B(new_n660), .Z(new_n661));
  OR2_X1    g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n654), .A2(new_n655), .ZN(new_n663));
  INV_X1    g462(.A(new_n646), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n657), .A2(new_n646), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n661), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n644), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n565), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n515), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(G1gat), .Z(G1324gat));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n518), .A2(new_n534), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n565), .A2(new_n675), .A3(new_n669), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n673), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT104), .Z(new_n679));
  OR3_X1    g478(.A1(new_n676), .A2(new_n673), .A3(new_n677), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT105), .B1(new_n676), .B2(G8gat), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n676), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n679), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT36), .B1(new_n510), .B2(new_n473), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT74), .B(new_n506), .C1(new_n508), .C2(new_n509), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n507), .A2(KEYINPUT106), .A3(new_n511), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n670), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n510), .A2(G15gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n670), .B2(new_n691), .ZN(G1326gat));
  NOR2_X1   g491(.A1(new_n670), .A2(new_n325), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  NOR3_X1   g494(.A1(new_n611), .A2(new_n643), .A3(new_n668), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT107), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n565), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(new_n515), .A3(new_n202), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT45), .Z(new_n700));
  NAND3_X1  g499(.A1(new_n689), .A2(new_n519), .A3(new_n551), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n564), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n606), .A2(new_n610), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n552), .A2(new_n564), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n611), .A2(new_n705), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n704), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n643), .A2(new_n263), .A3(new_n668), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n202), .B1(new_n710), .B2(new_n515), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n700), .A2(new_n711), .ZN(G1328gat));
  NOR3_X1   g511(.A1(new_n698), .A2(G36gat), .A3(new_n674), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT46), .ZN(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n710), .B2(new_n674), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1329gat));
  INV_X1    g515(.A(G43gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n706), .A2(new_n707), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n519), .A2(new_n687), .A3(new_n688), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n719), .A2(new_n551), .B1(new_n560), .B2(new_n563), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n705), .B1(new_n720), .B2(new_n611), .ZN(new_n721));
  INV_X1    g520(.A(new_n689), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n718), .A2(new_n721), .A3(new_n722), .A4(new_n709), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n708), .A2(KEYINPUT108), .A3(new_n722), .A4(new_n709), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n510), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n565), .A2(new_n717), .A3(new_n728), .A4(new_n697), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT47), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n723), .A2(G43gat), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT47), .B1(new_n734), .B2(new_n729), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n730), .B1(new_n725), .B2(new_n726), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT109), .B1(new_n738), .B2(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1330gat));
  INV_X1    g539(.A(new_n698), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n325), .A2(G50gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n741), .A2(new_n742), .B1(KEYINPUT110), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n718), .A2(new_n721), .A3(new_n514), .A4(new_n709), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n744), .B2(new_n746), .ZN(new_n749));
  OAI22_X1  g548(.A1(new_n748), .A2(new_n749), .B1(KEYINPUT110), .B2(new_n743), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n746), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT111), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n743), .A2(KEYINPUT110), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n750), .A2(new_n755), .ZN(G1331gat));
  INV_X1    g555(.A(new_n644), .ZN(new_n757));
  INV_X1    g556(.A(new_n263), .ZN(new_n758));
  INV_X1    g557(.A(new_n668), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n702), .A2(KEYINPUT112), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n757), .A2(new_n760), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n720), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n380), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g567(.A1(new_n765), .A2(new_n674), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(G1333gat));
  OAI21_X1  g572(.A(G71gat), .B1(new_n765), .B2(new_n689), .ZN(new_n774));
  INV_X1    g573(.A(G71gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n728), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n765), .B2(new_n776), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g577(.A1(new_n765), .A2(new_n325), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT113), .B(G78gat), .Z(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1335gat));
  INV_X1    g580(.A(new_n643), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n760), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n708), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(G85gat), .B1(new_n785), .B2(new_n515), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n263), .ZN(new_n787));
  AOI211_X1 g586(.A(new_n611), .B(new_n787), .C1(new_n701), .C2(new_n564), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n380), .A2(new_n576), .A3(new_n668), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n786), .B1(new_n790), .B2(new_n791), .ZN(G1336gat));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n718), .A2(new_n721), .A3(new_n675), .A4(new_n784), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n674), .A2(G92gat), .A3(new_n759), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n793), .B(new_n795), .C1(new_n790), .C2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT114), .B1(new_n800), .B2(KEYINPUT51), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n611), .B1(new_n701), .B2(new_n564), .ZN(new_n802));
  INV_X1    g601(.A(new_n787), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT115), .B1(new_n788), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n805), .B(new_n796), .C1(new_n807), .C2(KEYINPUT51), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n795), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n799), .B1(new_n809), .B2(KEYINPUT52), .ZN(new_n810));
  AOI211_X1 g609(.A(KEYINPUT116), .B(new_n793), .C1(new_n808), .C2(new_n795), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n798), .B1(new_n810), .B2(new_n811), .ZN(G1337gat));
  OAI21_X1  g611(.A(G99gat), .B1(new_n785), .B2(new_n689), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n510), .A2(new_n759), .A3(G99gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n790), .B2(new_n814), .ZN(G1338gat));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n759), .A2(new_n325), .A3(G106gat), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n790), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n718), .A2(new_n721), .A3(new_n514), .A4(new_n784), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n702), .A2(new_n806), .A3(new_n703), .A4(new_n803), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n800), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n804), .B1(new_n824), .B2(new_n789), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT117), .B1(new_n825), .B2(new_n817), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT51), .B1(new_n823), .B2(new_n800), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n827), .A2(new_n828), .A3(new_n804), .A4(new_n818), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n826), .A2(new_n829), .A3(new_n821), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n822), .B1(new_n830), .B2(new_n816), .ZN(G1339gat));
  NAND4_X1  g630(.A1(new_n243), .A2(new_n246), .A3(new_n251), .A4(new_n261), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n235), .B1(new_n245), .B2(new_n234), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n249), .A2(new_n250), .A3(new_n247), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n258), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n654), .A2(new_n655), .A3(new_n646), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n661), .B1(new_n656), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n843), .A2(new_n667), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n703), .A2(new_n836), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n252), .A2(new_n253), .A3(new_n261), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n261), .B1(new_n252), .B2(new_n253), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n667), .A3(new_n844), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n668), .A2(new_n835), .A3(new_n832), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n611), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n643), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n644), .A2(new_n758), .A3(new_n668), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n515), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n856), .A2(new_n674), .A3(new_n557), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT118), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n335), .A3(new_n758), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n674), .A2(new_n380), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n855), .A2(new_n553), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n263), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(G1340gat));
  NAND3_X1  g662(.A1(new_n858), .A2(new_n333), .A3(new_n668), .ZN(new_n864));
  OAI21_X1  g663(.A(G120gat), .B1(new_n861), .B2(new_n759), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1341gat));
  INV_X1    g665(.A(G127gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n857), .A2(new_n867), .A3(new_n643), .ZN(new_n868));
  OAI21_X1  g667(.A(G127gat), .B1(new_n861), .B2(new_n782), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1342gat));
  INV_X1    g669(.A(G134gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n857), .A2(new_n871), .A3(new_n703), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n861), .B2(new_n611), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  NOR3_X1   g675(.A1(new_n722), .A2(new_n675), .A3(new_n325), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n856), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n263), .A2(G141gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n850), .B2(new_n851), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n836), .A2(new_n668), .ZN(new_n886));
  OAI211_X1 g685(.A(KEYINPUT120), .B(new_n886), .C1(new_n263), .C2(new_n849), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n611), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n643), .B1(new_n888), .B2(new_n846), .ZN(new_n889));
  OAI211_X1 g688(.A(KEYINPUT57), .B(new_n514), .C1(new_n889), .C2(new_n854), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n514), .B1(new_n853), .B2(new_n854), .ZN(new_n891));
  XOR2_X1   g690(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n689), .A2(new_n380), .A3(new_n674), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n758), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n276), .B1(new_n897), .B2(KEYINPUT121), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n263), .B(new_n895), .C1(new_n890), .C2(new_n893), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n883), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n897), .A2(G141gat), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n882), .B1(new_n903), .B2(new_n881), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT122), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n883), .ZN(new_n906));
  OAI21_X1  g705(.A(G141gat), .B1(new_n899), .B2(new_n900), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n903), .A2(new_n881), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT58), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n905), .A2(new_n913), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n879), .A2(new_n277), .A3(new_n668), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n889), .A2(new_n854), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT57), .B1(new_n917), .B2(new_n514), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n891), .A2(new_n892), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n668), .A3(new_n896), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n916), .B1(new_n921), .B2(G148gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n895), .B1(new_n890), .B2(new_n893), .ZN(new_n923));
  AOI211_X1 g722(.A(KEYINPUT59), .B(new_n277), .C1(new_n923), .C2(new_n668), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n915), .B1(new_n922), .B2(new_n924), .ZN(G1345gat));
  AND2_X1   g724(.A1(new_n923), .A2(new_n643), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n643), .A2(new_n267), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n926), .A2(new_n267), .B1(new_n878), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT123), .ZN(G1346gat));
  AOI21_X1  g728(.A(G162gat), .B1(new_n879), .B2(new_n703), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n611), .A2(new_n268), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n923), .B2(new_n931), .ZN(G1347gat));
  NOR3_X1   g731(.A1(new_n855), .A2(new_n380), .A3(new_n674), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n561), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n398), .A3(new_n263), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n557), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n758), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n935), .B1(new_n398), .B2(new_n938), .ZN(G1348gat));
  OAI21_X1  g738(.A(new_n399), .B1(new_n936), .B2(new_n759), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT124), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n934), .A2(new_n399), .A3(new_n759), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n934), .B2(new_n782), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n643), .A2(new_n382), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n936), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n946), .B(new_n947), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n937), .A2(new_n384), .A3(new_n703), .ZN(new_n949));
  OAI21_X1  g748(.A(G190gat), .B1(new_n934), .B2(new_n611), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(KEYINPUT61), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(KEYINPUT61), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1351gat));
  INV_X1    g752(.A(G197gat), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n674), .A2(new_n380), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n689), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n758), .B(new_n957), .C1(new_n918), .C2(new_n919), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n959), .B2(new_n958), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n891), .A2(new_n956), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n954), .A3(new_n758), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT126), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n961), .A2(new_n964), .ZN(G1352gat));
  INV_X1    g764(.A(G204gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n962), .A2(new_n966), .A3(new_n668), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT62), .Z(new_n968));
  INV_X1    g767(.A(new_n920), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n969), .A2(new_n759), .A3(new_n956), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n970), .B2(new_n966), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n962), .A2(new_n290), .A3(new_n643), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n920), .A2(new_n643), .A3(new_n957), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  NAND3_X1  g775(.A1(new_n962), .A2(new_n291), .A3(new_n703), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n969), .A2(new_n611), .A3(new_n956), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n291), .ZN(G1355gat));
endmodule


