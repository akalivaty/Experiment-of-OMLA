//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G116), .B2(G270), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G77), .A2(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n203), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n212), .B(new_n227), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT65), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n220), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT66), .B1(new_n251), .B2(new_n253), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G226), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G222), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n263), .B(new_n265), .C1(new_n266), .C2(new_n264), .ZN(new_n267));
  INV_X1    g0067(.A(new_n251), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n267), .B(new_n268), .C1(G77), .C2(new_n263), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n259), .A2(new_n262), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G190), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(G200), .ZN(new_n273));
  OAI21_X1  g0073(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT67), .ZN(new_n275));
  XOR2_X1   g0075(.A(KEYINPUT8), .B(G58), .Z(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n276), .A2(new_n278), .B1(G150), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n228), .B1(new_n209), .B2(new_n277), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n252), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n281), .A2(new_n282), .B1(new_n220), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT9), .ZN(new_n290));
  INV_X1    g0090(.A(new_n282), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n229), .A2(G1), .ZN(new_n293));
  OR3_X1    g0093(.A1(new_n292), .A2(new_n220), .A3(new_n293), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n289), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n290), .B1(new_n289), .B2(new_n294), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n272), .B(new_n273), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n270), .A2(KEYINPUT70), .A3(G200), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT70), .B1(new_n270), .B2(G200), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT10), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n272), .C1(new_n296), .C2(new_n295), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n261), .B1(new_n258), .B2(G244), .ZN(new_n304));
  AND2_X1   g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(G238), .B2(G1698), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n224), .B2(G1698), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G107), .B2(new_n263), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n304), .B1(new_n310), .B2(new_n251), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n287), .A2(KEYINPUT69), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT69), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n285), .A2(new_n314), .A3(new_n286), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n316), .A2(new_n293), .A3(new_n282), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT15), .B(G87), .Z(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n278), .ZN(new_n319));
  INV_X1    g0119(.A(G77), .ZN(new_n320));
  INV_X1    g0120(.A(new_n276), .ZN(new_n321));
  INV_X1    g0121(.A(new_n279), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n319), .B1(new_n229), .B2(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n317), .A2(G77), .B1(new_n282), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n316), .A2(new_n320), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n311), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n312), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n289), .A2(new_n294), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n270), .A2(new_n327), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(G179), .B2(new_n270), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n324), .B(new_n325), .C1(new_n311), .C2(new_n271), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n311), .A2(G200), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n303), .A2(new_n329), .A3(new_n334), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT71), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n298), .B2(new_n302), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT71), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n329), .A4(new_n337), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n317), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n215), .B1(new_n344), .B2(KEYINPUT12), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n278), .A2(G77), .B1(G20), .B2(new_n215), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n220), .B2(new_n322), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n282), .ZN(new_n348));
  XOR2_X1   g0148(.A(new_n348), .B(KEYINPUT11), .Z(new_n349));
  NAND3_X1  g0149(.A1(new_n316), .A2(KEYINPUT12), .A3(new_n215), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n288), .A2(KEYINPUT12), .ZN(new_n352));
  NOR4_X1   g0152(.A1(new_n345), .A2(new_n349), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT72), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  OAI21_X1  g0156(.A(G238), .B1(new_n256), .B2(new_n257), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n224), .A2(G1698), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n358), .B1(G226), .B2(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n268), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n357), .A2(new_n362), .A3(new_n262), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n357), .A2(new_n362), .A3(new_n365), .A4(new_n262), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n356), .B1(new_n367), .B2(G169), .ZN(new_n368));
  AOI211_X1 g0168(.A(KEYINPUT14), .B(new_n327), .C1(new_n364), .C2(new_n366), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(G179), .A3(new_n366), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n355), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n371), .ZN(new_n373));
  NOR4_X1   g0173(.A1(new_n368), .A2(new_n369), .A3(new_n373), .A4(KEYINPUT72), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n354), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n367), .A2(G200), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n353), .B(new_n376), .C1(new_n271), .C2(new_n367), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT78), .ZN(new_n379));
  AND2_X1   g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n380), .B2(new_n202), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n279), .A2(G159), .ZN(new_n384));
  OAI211_X1 g0184(.A(KEYINPUT73), .B(G20), .C1(new_n380), .C2(new_n202), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT74), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT74), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n383), .A2(new_n388), .A3(new_n384), .A4(new_n385), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n307), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n307), .B2(new_n229), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT75), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  INV_X1    g0197(.A(new_n394), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n386), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n390), .A2(new_n400), .A3(KEYINPUT16), .A4(new_n394), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n396), .A2(new_n282), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n292), .A2(new_n293), .A3(new_n321), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n288), .B2(new_n321), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n266), .A2(new_n264), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n221), .A2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(new_n407), .C1(new_n305), .C2(new_n306), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n261), .B1(new_n410), .B2(new_n268), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n251), .A2(G232), .A3(new_n253), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n327), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n251), .B1(new_n408), .B2(new_n409), .ZN(new_n414));
  INV_X1    g0214(.A(new_n412), .ZN(new_n415));
  INV_X1    g0215(.A(G179), .ZN(new_n416));
  NOR4_X1   g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(new_n261), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT76), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n411), .A2(G179), .A3(new_n412), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT76), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n414), .A2(new_n261), .A3(new_n415), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n420), .C1(new_n327), .C2(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT18), .B1(new_n405), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  AOI211_X1 g0226(.A(new_n426), .B(new_n423), .C1(new_n402), .C2(new_n404), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n421), .A2(new_n271), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G200), .B2(new_n421), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n402), .A2(new_n404), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(KEYINPUT77), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n402), .A2(new_n435), .A3(new_n404), .A4(new_n430), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n379), .B1(new_n428), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n405), .A2(new_n424), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n426), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n405), .A2(KEYINPUT18), .A3(new_n424), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n433), .A2(new_n436), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT78), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n378), .B1(new_n438), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n343), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(KEYINPUT79), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n343), .B2(new_n445), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n277), .A2(G1), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n292), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G107), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n287), .A2(G107), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT25), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT24), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(KEYINPUT89), .ZN(new_n457));
  AND2_X1   g0257(.A1(KEYINPUT88), .A2(G87), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n229), .B(new_n458), .C1(new_n305), .C2(new_n306), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n263), .A2(new_n461), .A3(new_n229), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n206), .A2(G20), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n465), .B(KEYINPUT23), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n456), .A2(KEYINPUT89), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n466), .B1(new_n460), .B2(new_n462), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(new_n469), .A3(new_n464), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n457), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n453), .B(new_n455), .C1(new_n474), .C2(new_n291), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n263), .B1(G257), .B2(new_n264), .ZN(new_n476));
  NOR2_X1   g0276(.A1(G250), .A2(G1698), .ZN(new_n477));
  INV_X1    g0277(.A(G294), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n476), .A2(new_n477), .B1(new_n277), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n268), .ZN(new_n480));
  INV_X1    g0280(.A(G41), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n252), .B(G45), .C1(new_n481), .C2(KEYINPUT5), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G41), .ZN(new_n484));
  OAI211_X1 g0284(.A(G264), .B(new_n251), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(KEYINPUT80), .ZN(new_n486));
  AND2_X1   g0286(.A1(G1), .A2(G13), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n250), .B1(KEYINPUT5), .B2(new_n481), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n483), .A2(G41), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n252), .A4(G45), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n486), .A2(new_n488), .A3(new_n491), .A4(G274), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n480), .A2(new_n485), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT90), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n485), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n480), .A3(new_n492), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n493), .A2(new_n327), .B1(new_n496), .B2(new_n416), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n475), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n457), .ZN(new_n499));
  AND4_X1   g0299(.A1(new_n469), .A2(new_n463), .A3(new_n464), .A4(new_n467), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n469), .B1(new_n472), .B2(new_n464), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n282), .ZN(new_n503));
  INV_X1    g0303(.A(G200), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n480), .A2(new_n271), .A3(new_n485), .A4(new_n492), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n503), .A2(new_n507), .A3(new_n453), .A4(new_n455), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n498), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(G107), .B1(new_n392), .B2(new_n393), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n279), .A2(G77), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT6), .B1(new_n207), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n205), .A2(G107), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(KEYINPUT6), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n510), .B(new_n511), .C1(new_n229), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n282), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n287), .A2(G97), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n292), .A2(new_n205), .A3(new_n451), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n492), .ZN(new_n523));
  OAI21_X1  g0323(.A(G244), .B1(new_n305), .B2(new_n306), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n524), .A2(new_n525), .B1(G33), .B2(G283), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n264), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n525), .B1(new_n263), .B2(G250), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n264), .C2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n523), .B1(new_n529), .B2(new_n268), .ZN(new_n530));
  OAI211_X1 g0330(.A(G257), .B(new_n251), .C1(new_n482), .C2(new_n484), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n327), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n416), .A3(new_n531), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n522), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(G200), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n520), .B1(new_n516), .B2(new_n282), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n530), .A2(G190), .A3(new_n531), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n536), .A2(new_n519), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n285), .A2(new_n314), .A3(new_n286), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n314), .B1(new_n285), .B2(new_n286), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G116), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n451), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(KEYINPUT85), .A3(new_n291), .A4(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n313), .A2(new_n315), .A3(new_n291), .A4(new_n547), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT85), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n316), .A2(new_n546), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G283), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n553), .B(new_n229), .C1(G33), .C2(new_n205), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n546), .A2(G20), .ZN(new_n555));
  OR2_X1    g0355(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n554), .A2(new_n282), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n557), .B(new_n558), .ZN(new_n559));
  AND4_X1   g0359(.A1(new_n548), .A2(new_n551), .A3(new_n552), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n264), .A2(G257), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G264), .A2(G1698), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n305), .C2(new_n306), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n563), .B(new_n268), .C1(G303), .C2(new_n263), .ZN(new_n564));
  OAI211_X1 g0364(.A(G270), .B(new_n251), .C1(new_n482), .C2(new_n484), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n492), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT84), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT84), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n564), .A2(new_n492), .A3(new_n568), .A4(new_n565), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(G169), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n542), .B1(new_n560), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n567), .A2(KEYINPUT21), .A3(G169), .A4(new_n569), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n566), .A2(new_n416), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n548), .A2(new_n551), .A3(new_n552), .A4(new_n559), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n567), .A2(new_n569), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n567), .A2(G200), .A3(new_n569), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n560), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n571), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  OAI211_X1 g0383(.A(G244), .B(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT81), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n263), .A2(KEYINPUT81), .A3(G244), .A4(G1698), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G116), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n263), .A2(G238), .A3(new_n264), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n268), .ZN(new_n591));
  INV_X1    g0391(.A(G250), .ZN(new_n592));
  INV_X1    g0392(.A(G45), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(G1), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n252), .A2(new_n260), .A3(G45), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n251), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n327), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n596), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n416), .B(new_n598), .C1(new_n590), .C2(new_n268), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n583), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n591), .A2(G179), .A3(new_n596), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n590), .B2(new_n268), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(KEYINPUT82), .C1(new_n327), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n452), .A2(new_n318), .ZN(new_n604));
  INV_X1    g0404(.A(new_n318), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n543), .B2(new_n544), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT83), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n360), .A2(new_n229), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n608), .B(KEYINPUT19), .C1(new_n207), .C2(G87), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n229), .B(G68), .C1(new_n305), .C2(new_n306), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT19), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n360), .B2(G20), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n282), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n606), .A2(new_n607), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n607), .B1(new_n606), .B2(new_n614), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n604), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n600), .A2(new_n603), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n606), .A2(new_n614), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT83), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n606), .A2(new_n607), .A3(new_n614), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n602), .A2(new_n504), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n602), .A2(G190), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n452), .A2(G87), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n582), .A2(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n450), .A2(new_n509), .A3(new_n541), .A4(new_n628), .ZN(G372));
  NOR2_X1   g0429(.A1(new_n627), .A2(new_n535), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n601), .B1(new_n327), .B2(new_n602), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n617), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n635), .B2(new_n535), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT91), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n533), .A2(new_n534), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(new_n522), .A3(new_n626), .A4(new_n634), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(KEYINPUT91), .A3(new_n632), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n631), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n634), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n505), .A2(new_n506), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n475), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n540), .A2(new_n645), .A3(new_n635), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n567), .A2(new_n569), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n576), .A2(new_n647), .A3(G169), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n542), .B1(new_n575), .B2(new_n576), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n498), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n643), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n642), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n450), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n413), .A2(new_n417), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n402), .B2(new_n404), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  INV_X1    g0456(.A(new_n375), .ZN(new_n657));
  INV_X1    g0457(.A(new_n329), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n377), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n656), .B1(new_n659), .B2(new_n437), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n333), .B1(new_n660), .B2(new_n303), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(G369));
  INV_X1    g0462(.A(G13), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n252), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT95), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n475), .A2(new_n497), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n670), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n498), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n475), .A2(new_n670), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n509), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT93), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n509), .A2(KEYINPUT93), .A3(new_n676), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n649), .A2(new_n670), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT94), .Z(new_n683));
  OAI21_X1  g0483(.A(new_n673), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n576), .A2(new_n670), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n649), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n649), .A2(new_n581), .A3(new_n685), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(KEYINPUT92), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n689));
  OAI21_X1  g0489(.A(G330), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n681), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n684), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n210), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G1), .ZN(new_n696));
  INV_X1    g0496(.A(G87), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n697), .A2(new_n205), .A3(new_n206), .A4(new_n546), .ZN(new_n698));
  OAI22_X1  g0498(.A1(new_n696), .A2(new_n698), .B1(new_n231), .B2(new_n695), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n650), .B(KEYINPUT96), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n646), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n630), .A2(new_n632), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n643), .B1(new_n640), .B2(KEYINPUT26), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(KEYINPUT29), .A3(new_n674), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n671), .B1(new_n642), .B2(new_n651), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n628), .A2(new_n509), .A3(new_n541), .A4(new_n672), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n530), .A2(new_n495), .A3(new_n531), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n602), .A2(new_n480), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n573), .A4(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n530), .A2(new_n495), .A3(new_n573), .A4(new_n531), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n711), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n647), .A2(new_n532), .A3(new_n416), .A4(new_n496), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n713), .B(new_n716), .C1(new_n602), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n670), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n709), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n706), .A2(new_n708), .B1(G330), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n700), .B1(new_n724), .B2(G1), .ZN(G364));
  AOI21_X1  g0525(.A(new_n696), .B1(G45), .B2(new_n664), .ZN(new_n726));
  XOR2_X1   g0526(.A(G355), .B(KEYINPUT97), .Z(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n210), .A3(new_n263), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n245), .A2(new_n593), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n693), .A2(new_n263), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(G45), .B2(new_n231), .ZN(new_n731));
  OAI221_X1 g0531(.A(new_n728), .B1(G116), .B2(new_n210), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n228), .B1(G20), .B2(new_n327), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n229), .A2(new_n271), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n416), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G322), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n307), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n416), .A2(new_n504), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n229), .A2(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G317), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT33), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n748), .A2(KEYINPUT33), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n744), .A2(new_n739), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G326), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n745), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G329), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n504), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n745), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G283), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n751), .A2(new_n754), .A3(new_n758), .A4(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n229), .B1(new_n755), .B2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n743), .B(new_n763), .C1(G294), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G303), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n739), .A2(new_n759), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n745), .A2(new_n740), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n766), .B1(new_n767), .B2(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n757), .A2(G159), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n760), .A2(new_n206), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n752), .A2(new_n220), .B1(new_n768), .B2(new_n697), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n263), .B1(new_n764), .B2(new_n205), .C1(new_n320), .C2(new_n770), .ZN(new_n776));
  NOR4_X1   g0576(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n777), .B1(new_n223), .B2(new_n741), .C1(new_n215), .C2(new_n746), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n736), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n726), .B(new_n738), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n688), .A2(new_n689), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n735), .B(KEYINPUT99), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n726), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n690), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G330), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(new_n789), .B2(new_n784), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  NOR2_X1   g0592(.A1(new_n329), .A2(new_n670), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n326), .A2(new_n670), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n335), .B2(new_n336), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n329), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n707), .A2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n671), .B(new_n798), .C1(new_n642), .C2(new_n651), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n723), .A2(G330), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n787), .ZN(new_n805));
  INV_X1    g0605(.A(new_n741), .ZN(new_n806));
  INV_X1    g0606(.A(new_n770), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G143), .A2(new_n806), .B1(new_n807), .B2(G159), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  INV_X1    g0609(.A(G150), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n752), .C1(new_n810), .C2(new_n746), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT34), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n764), .A2(new_n223), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n760), .A2(new_n215), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n811), .C2(new_n812), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n263), .C1(new_n817), .C2(new_n756), .ZN(new_n818));
  INV_X1    g0618(.A(new_n768), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n813), .B(new_n818), .C1(G50), .C2(new_n819), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n752), .A2(new_n767), .B1(new_n770), .B2(new_n546), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G283), .B2(new_n747), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT100), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n741), .A2(new_n478), .B1(new_n764), .B2(new_n205), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT101), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n263), .B1(new_n824), .B2(KEYINPUT101), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n827), .B1(new_n697), .B2(new_n760), .C1(new_n769), .C2(new_n756), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n823), .B(new_n828), .C1(G107), .C2(new_n819), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n736), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n798), .A2(new_n733), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n736), .A2(new_n733), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n320), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n830), .A2(new_n831), .A3(new_n726), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n805), .A2(new_n834), .ZN(G384));
  NAND3_X1  g0635(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n709), .A2(new_n721), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT107), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT107), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n709), .A2(new_n839), .A3(new_n721), .A4(new_n836), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n450), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n390), .A2(new_n394), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n397), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n396), .A2(new_n844), .A3(new_n282), .A4(new_n401), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n668), .B1(new_n845), .B2(new_n404), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n428), .B2(new_n437), .ZN(new_n847));
  INV_X1    g0647(.A(new_n668), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n405), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n439), .A2(new_n849), .A3(new_n850), .A4(new_n431), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n402), .A2(new_n404), .A3(new_n430), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n654), .B1(new_n845), .B2(new_n404), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n852), .A2(new_n846), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n851), .B1(new_n854), .B2(new_n850), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n847), .A2(new_n855), .A3(KEYINPUT38), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT106), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n437), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n433), .A2(KEYINPUT106), .A3(new_n436), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n656), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n668), .B1(new_n402), .B2(new_n404), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT105), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n852), .A2(new_n655), .A3(new_n861), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n864), .B2(new_n850), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n849), .A2(new_n431), .ZN(new_n866));
  OAI211_X1 g0666(.A(KEYINPUT105), .B(KEYINPUT37), .C1(new_n866), .C2(new_n655), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n851), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n856), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n798), .B1(new_n838), .B2(new_n840), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n354), .A2(new_n670), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n375), .A2(new_n377), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n354), .B(new_n670), .C1(new_n372), .C2(new_n374), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT40), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  AOI221_X4 g0678(.A(new_n798), .B1(new_n874), .B2(new_n875), .C1(new_n838), .C2(new_n840), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT104), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n847), .A2(new_n855), .A3(new_n881), .A4(KEYINPUT38), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n852), .A2(new_n846), .ZN(new_n883));
  INV_X1    g0683(.A(new_n853), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n850), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND4_X1   g0685(.A1(new_n850), .A2(new_n439), .A3(new_n849), .A4(new_n431), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n846), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n442), .B2(new_n443), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n870), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n847), .A2(new_n855), .A3(KEYINPUT38), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(KEYINPUT104), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n879), .A2(new_n880), .A3(new_n882), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n878), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(G330), .B1(new_n842), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT108), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n895), .A2(new_n896), .B1(new_n894), .B2(new_n842), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n896), .B2(new_n895), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n656), .A2(new_n848), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT103), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n801), .A2(new_n900), .A3(new_n793), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n707), .A2(new_n799), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT103), .B1(new_n902), .B2(new_n794), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n876), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n892), .A2(new_n882), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n375), .A2(new_n670), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n871), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n892), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n706), .A2(new_n708), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n447), .B2(new_n449), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n661), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n913), .B(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n898), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n252), .B2(new_n664), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT35), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n515), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(G116), .A3(new_n230), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT102), .Z(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n920), .B2(new_n515), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT36), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n231), .A2(new_n320), .A3(new_n380), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n201), .A2(new_n215), .ZN(new_n927));
  OAI211_X1 g0727(.A(G1), .B(new_n663), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n919), .A2(new_n925), .A3(new_n928), .ZN(G367));
  OAI22_X1  g0729(.A1(new_n760), .A2(new_n205), .B1(new_n756), .B2(new_n748), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n307), .B1(new_n764), .B2(new_n206), .C1(new_n767), .C2(new_n741), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n930), .B(new_n931), .C1(G283), .C2(new_n807), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n753), .A2(G311), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n819), .A2(G116), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT46), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n747), .A2(G294), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n932), .A2(new_n933), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n753), .A2(G143), .B1(new_n765), .B2(G68), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n809), .B2(new_n756), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G159), .B2(new_n747), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n761), .A2(G77), .ZN(new_n941));
  INV_X1    g0741(.A(new_n201), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n940), .B(new_n941), .C1(new_n942), .C2(new_n770), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n263), .B1(new_n741), .B2(new_n810), .C1(new_n223), .C2(new_n768), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT47), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n736), .ZN(new_n947));
  INV_X1    g0747(.A(new_n730), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n737), .B1(new_n210), .B2(new_n605), .C1(new_n241), .C2(new_n948), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n947), .A2(new_n726), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n622), .A2(new_n625), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n643), .A2(new_n951), .A3(new_n670), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n670), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n626), .A3(new_n634), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n954), .A3(new_n785), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT111), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n522), .A2(new_n671), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n541), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n639), .A2(new_n522), .A3(new_n671), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n684), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT44), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n673), .B(new_n961), .C1(new_n681), .C2(new_n683), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT45), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n691), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n966), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT44), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n963), .B(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n691), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n683), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n681), .A2(new_n690), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n973), .B1(new_n975), .B2(new_n691), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n683), .A3(new_n974), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n724), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n967), .A2(new_n972), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n724), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n694), .B(KEYINPUT41), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n252), .B1(new_n664), .B2(G45), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n952), .A2(new_n954), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT109), .Z(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n535), .B1(new_n959), .B2(new_n498), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n672), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n681), .A2(new_n683), .A3(new_n962), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT42), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(new_n994), .ZN(new_n998));
  OAI211_X1 g0798(.A(KEYINPUT110), .B(new_n992), .C1(new_n993), .C2(new_n994), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n691), .A2(new_n961), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1001), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n990), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1005), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(new_n989), .A3(new_n1003), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n957), .B1(new_n986), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n985), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n982), .B2(new_n983), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1013), .A2(new_n1009), .A3(KEYINPUT111), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n956), .B1(new_n1011), .B2(new_n1014), .ZN(G387));
  NAND2_X1  g0815(.A1(new_n978), .A2(new_n1012), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n276), .A2(new_n220), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT50), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n215), .A2(new_n320), .ZN(new_n1019));
  NOR4_X1   g0819(.A1(new_n1018), .A2(G45), .A3(new_n1019), .A4(new_n698), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n730), .B1(new_n237), .B2(new_n593), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n263), .A2(new_n698), .A3(new_n210), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n210), .A2(G107), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n737), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n787), .B1(new_n681), .B2(new_n785), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G322), .A2(new_n753), .B1(new_n747), .B2(G311), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n767), .B2(new_n770), .C1(new_n748), .C2(new_n741), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  INV_X1    g0829(.A(G283), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n764), .C1(new_n478), .C2(new_n768), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n263), .B1(new_n757), .B2(G326), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n546), .C2(new_n760), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n263), .B1(new_n760), .B2(new_n205), .C1(new_n220), .C2(new_n741), .ZN(new_n1035));
  INV_X1    g0835(.A(G159), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n752), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT114), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n215), .B2(new_n770), .C1(new_n321), .C2(new_n746), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1035), .B(new_n1039), .C1(new_n318), .C2(new_n765), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(KEYINPUT112), .B(G150), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n768), .A2(new_n320), .B1(new_n756), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT113), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1040), .B(new_n1043), .C1(KEYINPUT114), .C2(new_n1037), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1034), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1025), .B(new_n1026), .C1(new_n1045), .C2(new_n780), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n694), .B1(new_n978), .B2(new_n724), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1016), .B(new_n1046), .C1(new_n980), .C2(new_n1047), .ZN(G393));
  INV_X1    g0848(.A(KEYINPUT115), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n972), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n971), .B1(new_n968), .B2(new_n970), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n967), .A2(new_n972), .A3(KEYINPUT115), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n1012), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n979), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n694), .A3(new_n981), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n787), .B1(new_n962), .B2(new_n735), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n737), .B1(new_n205), .B2(new_n210), .C1(new_n248), .C2(new_n948), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n760), .A2(new_n206), .B1(new_n756), .B2(new_n742), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1059), .A2(new_n263), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n478), .B2(new_n770), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n752), .A2(new_n748), .B1(new_n741), .B2(new_n769), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT52), .Z(new_n1063));
  AOI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(G116), .C2(new_n765), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n1030), .B2(new_n768), .C1(new_n767), .C2(new_n746), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n752), .A2(new_n810), .B1(new_n741), .B2(new_n1036), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  NOR2_X1   g0867(.A1(new_n321), .A2(new_n770), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n764), .A2(new_n320), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n942), .B2(new_n746), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n307), .B1(new_n757), .B2(G143), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n215), .B2(new_n768), .C1(new_n697), .C2(new_n760), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT116), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1065), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n736), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1057), .A2(new_n1058), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1054), .A2(new_n1056), .A3(new_n1077), .ZN(G390));
  NAND3_X1  g0878(.A1(new_n872), .A2(G330), .A3(new_n876), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n876), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n900), .B1(new_n801), .B2(new_n793), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n902), .A2(KEYINPUT103), .A3(new_n794), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n911), .B(new_n910), .C1(new_n1083), .C2(new_n907), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n871), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n705), .A2(new_n674), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n793), .B1(new_n1086), .B2(new_n797), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1085), .B(new_n908), .C1(new_n1087), .C2(new_n1080), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1079), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1080), .A2(new_n803), .A3(new_n798), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1084), .A2(new_n1092), .A3(new_n1088), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1090), .A2(new_n1012), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n910), .A2(new_n733), .A3(new_n911), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n832), .A2(new_n321), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT54), .B(G143), .Z(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1098), .A2(new_n770), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n768), .A2(new_n1041), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT53), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n765), .A2(G159), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n263), .B1(new_n741), .B2(new_n817), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G125), .B2(new_n757), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G128), .A2(new_n753), .B1(new_n761), .B2(new_n201), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1099), .B(new_n1106), .C1(G137), .C2(new_n747), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1069), .B(new_n815), .C1(G87), .C2(new_n819), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n753), .A2(G283), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n263), .B1(new_n747), .B2(G107), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G97), .A2(new_n807), .B1(new_n757), .B2(G294), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G116), .B2(new_n806), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n736), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1095), .A2(new_n726), .A3(new_n1096), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1094), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1084), .A2(new_n1092), .A3(new_n1088), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n1089), .ZN(new_n1118));
  OAI211_X1 g0918(.A(G330), .B(new_n841), .C1(new_n447), .C2(new_n449), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n661), .A3(new_n915), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n872), .A2(G330), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1091), .B1(new_n1121), .B2(new_n1080), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1080), .B1(new_n803), .B2(new_n798), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1079), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1122), .A2(new_n1087), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1118), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n695), .B1(new_n1118), .B2(new_n1127), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1116), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(G378));
  NAND3_X1  g0931(.A1(new_n1090), .A2(new_n1127), .A3(new_n1093), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1120), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n340), .B(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n330), .A2(new_n668), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n892), .A2(new_n880), .A3(new_n882), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT38), .B1(new_n862), .B2(new_n868), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n872), .B(new_n876), .C1(new_n1141), .C2(new_n856), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1140), .A2(new_n879), .B1(new_n1142), .B2(KEYINPUT40), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1139), .B1(new_n1143), .B2(new_n789), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1139), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n894), .A2(G330), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n913), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n910), .A2(new_n911), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n907), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1083), .A2(new_n882), .A3(new_n892), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n899), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1145), .B1(new_n894), .B2(G330), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n789), .B(new_n1139), .C1(new_n878), .C2(new_n893), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1134), .A2(KEYINPUT57), .A3(new_n1147), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1120), .B1(new_n1118), .B2(new_n1127), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT119), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n913), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1147), .A2(new_n1154), .A3(KEYINPUT119), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1156), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n694), .B(new_n1155), .C1(new_n1162), .C2(KEYINPUT57), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1147), .A2(new_n1154), .A3(KEYINPUT119), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT119), .B1(new_n1147), .B2(new_n1154), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1012), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n320), .A2(new_n768), .B1(new_n741), .B2(new_n206), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G41), .B(new_n1167), .C1(G68), .C2(new_n765), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n760), .A2(new_n223), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1169), .A2(new_n263), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n807), .A2(new_n318), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n747), .A2(G97), .B1(new_n757), .B2(G283), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G116), .B2(new_n753), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT117), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n220), .B1(new_n305), .B2(G41), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1174), .A2(KEYINPUT58), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G33), .B1(new_n757), .B2(G124), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n481), .C1(new_n1036), .C2(new_n760), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT118), .ZN(new_n1180));
  INV_X1    g0980(.A(G128), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n741), .A2(new_n1181), .B1(new_n770), .B2(new_n809), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1098), .A2(new_n768), .B1(new_n810), .B2(new_n764), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(G125), .C2(new_n753), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n817), .B2(new_n746), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT59), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1177), .B1(new_n1175), .B2(new_n1176), .C1(new_n1180), .C2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1174), .A2(KEYINPUT58), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n736), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n787), .B1(new_n942), .B2(new_n832), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n1139), .C2(new_n734), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1166), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1163), .A2(new_n1192), .ZN(G375));
  INV_X1    g0993(.A(KEYINPUT120), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1120), .A2(new_n1194), .A3(new_n1126), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n983), .B1(new_n1120), .B2(new_n1126), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n752), .A2(new_n817), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n768), .A2(new_n1036), .B1(new_n756), .B2(new_n1181), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT122), .Z(new_n1200));
  AOI22_X1  g1000(.A1(G137), .A2(new_n806), .B1(new_n747), .B2(new_n1097), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n810), .B2(new_n770), .ZN(new_n1202));
  OR4_X1    g1002(.A1(new_n307), .A2(new_n1200), .A3(new_n1169), .A4(new_n1202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1198), .B(new_n1203), .C1(G50), .C2(new_n765), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n819), .A2(G97), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G107), .A2(new_n807), .B1(new_n757), .B2(G303), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n1030), .B2(new_n741), .C1(new_n478), .C2(new_n752), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n941), .A2(new_n307), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT121), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n605), .B2(new_n764), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1207), .B(new_n1210), .C1(G116), .C2(new_n747), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1204), .B1(new_n1205), .B2(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT123), .Z(new_n1213));
  OAI221_X1 g1013(.A(new_n726), .B1(new_n734), .B2(new_n876), .C1(new_n1213), .C2(new_n780), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n215), .B2(new_n832), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1126), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n1012), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1197), .A2(new_n1217), .ZN(G381));
  NAND3_X1  g1018(.A1(new_n986), .A2(new_n1010), .A3(new_n957), .ZN(new_n1219));
  OAI21_X1  g1019(.A(KEYINPUT111), .B1(new_n1013), .B2(new_n1009), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(G390), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n956), .A3(new_n1222), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1223), .A2(G396), .A3(G393), .ZN(new_n1224));
  INV_X1    g1024(.A(G384), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(new_n1217), .A4(new_n1197), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT124), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1166), .A2(new_n1191), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1134), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT57), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n695), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1230), .B1(new_n1233), .B2(new_n1155), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1130), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1228), .A2(new_n1229), .A3(new_n1235), .ZN(G407));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G343), .C2(new_n1235), .ZN(G409));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1130), .B1(new_n1163), .B2(new_n1192), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1195), .A2(new_n1196), .B1(new_n1127), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n1126), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n694), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G384), .B1(new_n1243), .B2(new_n1217), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(G384), .A3(new_n1217), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n983), .B(new_n1134), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1147), .A2(new_n1154), .A3(new_n1012), .ZN(new_n1249));
  AND4_X1   g1049(.A1(new_n1130), .A2(new_n1248), .A3(new_n1191), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G213), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(G343), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1239), .A2(new_n1247), .A3(new_n1250), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1239), .A2(new_n1252), .A3(new_n1250), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1246), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G2897), .B(new_n1252), .C1(new_n1256), .C2(new_n1244), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1252), .A2(G2897), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1245), .A2(new_n1246), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1253), .A2(new_n1254), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G375), .A2(G378), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1247), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1252), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1250), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1262), .B1(new_n1267), .B2(KEYINPUT62), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1238), .B1(new_n1261), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1266), .B(new_n1265), .C1(new_n1234), .C2(new_n1130), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1260), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1267), .A2(KEYINPUT62), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1273), .A3(KEYINPUT126), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1222), .B1(new_n1221), .B2(new_n956), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n956), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1277), .B(G390), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1275), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(G390), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(KEYINPUT125), .A3(new_n1223), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(G393), .B(new_n791), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1283), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1280), .A2(new_n1223), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1284), .B1(new_n1290), .B2(new_n1275), .ZN(new_n1291));
  OAI21_X1  g1091(.A(KEYINPUT127), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1269), .A2(new_n1274), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1253), .A2(KEYINPUT63), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1295), .B(new_n1296), .C1(new_n1253), .C2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(G405));
  NAND2_X1  g1100(.A1(new_n1235), .A2(new_n1263), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1264), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1235), .A2(new_n1263), .A3(new_n1247), .ZN(new_n1303));
  AND4_X1   g1103(.A1(new_n1292), .A2(new_n1288), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1288), .A2(new_n1292), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(G402));
endmodule


