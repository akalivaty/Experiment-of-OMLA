//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G57), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(G567), .A2(new_n454), .B1(new_n456), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n465), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  AND2_X1   g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(new_n474), .B2(G112), .ZN(new_n478));
  OAI22_X1  g053(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n479), .B1(G124), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT69), .ZN(G162));
  NAND3_X1  g058(.A1(new_n468), .A2(G138), .A3(new_n474), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT3), .B1(new_n463), .B2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(G126), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n474), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(G2105), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .A3(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G62), .ZN(new_n504));
  INV_X1    g079(.A(G75), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(new_n498), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G651), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT70), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(new_n509), .A3(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n503), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n514), .ZN(new_n518));
  INV_X1    g093(.A(new_n510), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(G543), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n516), .A2(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n508), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  INV_X1    g099(.A(new_n516), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  AOI211_X1 g101(.A(new_n498), .B(new_n510), .C1(new_n512), .C2(new_n514), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n526), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n516), .A2(new_n534), .B1(new_n520), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n511), .B2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n511), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n525), .A2(G81), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n527), .A2(G43), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  AND2_X1   g129(.A1(new_n525), .A2(G91), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n500), .A2(KEYINPUT76), .A3(new_n502), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT76), .B1(new_n500), .B2(new_n502), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  NOR3_X1   g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT77), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n564), .B(G651), .C1(new_n559), .C2(new_n561), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n555), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n518), .A2(G53), .A3(G543), .A4(new_n519), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT73), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(new_n570), .A3(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n527), .A2(new_n574), .A3(new_n575), .A4(G53), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n515), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n572), .A2(new_n573), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n573), .B1(new_n572), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n566), .B1(new_n580), .B2(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n525), .A2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n527), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  AOI22_X1  g161(.A1(new_n503), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n511), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n525), .A2(G86), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n527), .A2(G48), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G305));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n516), .A2(new_n592), .B1(new_n520), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n511), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n520), .A2(KEYINPUT79), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n520), .A2(KEYINPUT79), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n601), .A2(G54), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n518), .A2(new_n503), .A3(G92), .A4(new_n519), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  NOR3_X1   g182(.A1(new_n556), .A2(new_n557), .A3(new_n607), .ZN(new_n608));
  AND2_X1   g183(.A1(G79), .A2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n603), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n603), .A2(new_n606), .A3(KEYINPUT80), .A4(new_n610), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n600), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n600), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND3_X1  g199(.A1(new_n613), .A2(new_n623), .A3(new_n614), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g202(.A1(new_n613), .A2(KEYINPUT81), .A3(new_n623), .A4(new_n614), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n481), .A2(G123), .ZN(new_n633));
  INV_X1    g208(.A(new_n475), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G135), .ZN(new_n635));
  NOR2_X1   g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n633), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(G2096), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2430), .Z(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(new_n652));
  INV_X1    g227(.A(G2438), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(KEYINPUT84), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(KEYINPUT84), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G2438), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n650), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n649), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n650), .ZN(new_n661));
  INV_X1    g236(.A(new_n657), .ZN(new_n662));
  AOI21_X1  g237(.A(G2438), .B1(new_n655), .B2(new_n656), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n664), .A2(KEYINPUT85), .A3(KEYINPUT14), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n654), .A2(new_n650), .A3(new_n657), .ZN(new_n667));
  XOR2_X1   g242(.A(G2451), .B(G2454), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT83), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT16), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1341), .B(G1348), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n671), .B1(new_n666), .B2(new_n667), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(KEYINPUT85), .B1(new_n664), .B2(KEYINPUT14), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n658), .A2(new_n649), .A3(new_n659), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n667), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(new_n670), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n674), .B1(new_n681), .B2(new_n672), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n648), .B1(new_n677), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n675), .B1(new_n673), .B2(new_n676), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n674), .A3(new_n672), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(new_n685), .A3(new_n647), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(G14), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G401));
  INV_X1    g263(.A(G2100), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  XNOR2_X1  g265(.A(G2072), .B(G2078), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(KEYINPUT86), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(KEYINPUT86), .B2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(G2084), .B(G2090), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n690), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT17), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n691), .B(new_n697), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n693), .B(new_n695), .C1(new_n696), .C2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(KEYINPUT87), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(KEYINPUT87), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n698), .A2(new_n694), .A3(new_n696), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT88), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n694), .A2(new_n690), .A3(new_n691), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT18), .Z(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G2096), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n704), .B1(new_n701), .B2(new_n700), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n639), .B1(new_n710), .B2(new_n707), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n689), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(G2096), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n639), .A3(new_n707), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n713), .A2(G2100), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n715), .ZN(G227));
  XNOR2_X1  g291(.A(KEYINPUT22), .B(G1981), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(G1971), .B(G1976), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT19), .ZN(new_n720));
  XOR2_X1   g295(.A(G1956), .B(G2474), .Z(new_n721));
  XOR2_X1   g296(.A(G1961), .B(G1966), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT20), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n721), .A2(new_n722), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n720), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n724), .B2(new_n725), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n720), .A2(new_n727), .A3(new_n723), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n726), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT21), .B(G1986), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(G1991), .B(G1996), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n726), .A2(new_n729), .A3(new_n730), .A4(new_n732), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n736), .B1(new_n734), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n718), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n734), .A2(new_n737), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(new_n735), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n743), .A2(new_n717), .A3(new_n738), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(G229));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(G34), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n472), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G2084), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n548), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G16), .B2(G19), .ZN(new_n755));
  INV_X1    g330(.A(G1341), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT30), .B(G28), .Z(new_n757));
  OAI22_X1  g332(.A1(new_n755), .A2(new_n756), .B1(G29), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n756), .B2(new_n755), .ZN(new_n759));
  INV_X1    g334(.A(G16), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G4), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n615), .B2(G16), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AND4_X1   g341(.A1(new_n753), .A2(new_n759), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n634), .A2(G141), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT97), .Z(new_n769));
  AND3_X1   g344(.A1(new_n474), .A2(G105), .A3(G2104), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT26), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n770), .B(new_n772), .C1(new_n481), .C2(G129), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G29), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G29), .B2(G32), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT98), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G29), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G27), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n781), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2078), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G2084), .B2(new_n752), .ZN(new_n785));
  NOR2_X1   g360(.A1(G5), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G171), .B2(G16), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G1961), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n767), .A2(new_n780), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n787), .A2(G1961), .ZN(new_n790));
  INV_X1    g365(.A(G11), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n790), .B1(KEYINPUT31), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT25), .Z(new_n794));
  INV_X1    g369(.A(G139), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n794), .B1(new_n795), .B2(new_n475), .C1(new_n474), .C2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G33), .B(new_n797), .S(G29), .Z(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G2072), .Z(new_n799));
  OAI211_X1 g374(.A(new_n792), .B(new_n799), .C1(KEYINPUT31), .C2(new_n791), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT99), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G16), .B2(G21), .ZN(new_n802));
  NOR2_X1   g377(.A1(G286), .A2(new_n760), .ZN(new_n803));
  MUX2_X1   g378(.A(new_n802), .B(new_n801), .S(new_n803), .Z(new_n804));
  INV_X1    g379(.A(G1966), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n781), .A2(G26), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(new_n474), .B2(G116), .ZN(new_n808));
  INV_X1    g383(.A(G104), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n474), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n481), .B2(G128), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n812));
  INV_X1    g387(.A(G140), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n475), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n634), .A2(KEYINPUT96), .A3(G140), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n811), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n807), .B1(new_n817), .B2(new_n781), .ZN(new_n818));
  MUX2_X1   g393(.A(new_n807), .B(new_n818), .S(KEYINPUT28), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G2067), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n789), .A2(new_n800), .A3(new_n806), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(G29), .A2(G35), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G162), .B2(G29), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT29), .B(G2090), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n638), .A2(new_n781), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n776), .A2(new_n779), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n821), .A2(new_n825), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT92), .B1(G16), .B2(G23), .ZN(new_n831));
  OR3_X1    g406(.A1(KEYINPUT92), .A2(G16), .A3(G23), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n831), .B(new_n832), .C1(G288), .C2(new_n760), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT93), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT33), .B(G1976), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n760), .A2(G22), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G166), .B2(new_n760), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G1971), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  MUX2_X1   g415(.A(G6), .B(G305), .S(G16), .Z(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT32), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G1981), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT34), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n838), .A2(G1971), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n840), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G1981), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n842), .B(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n836), .A2(new_n845), .A3(new_n839), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT34), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(new_n474), .B2(G107), .ZN(new_n851));
  INV_X1    g426(.A(G95), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(new_n474), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n634), .B2(G131), .ZN(new_n854));
  INV_X1    g429(.A(G119), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n480), .A2(KEYINPUT90), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT90), .B1(new_n480), .B2(new_n855), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G29), .ZN(new_n859));
  INV_X1    g434(.A(G25), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT89), .B1(new_n860), .B2(G29), .ZN(new_n861));
  OR3_X1    g436(.A1(new_n860), .A2(KEYINPUT89), .A3(G29), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(KEYINPUT35), .B(G1991), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n863), .B(new_n864), .Z(new_n865));
  INV_X1    g440(.A(KEYINPUT91), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n760), .A2(G24), .ZN(new_n867));
  AOI211_X1 g442(.A(new_n866), .B(new_n867), .C1(G290), .C2(G16), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  INV_X1    g444(.A(G1986), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n846), .A2(new_n850), .A3(new_n865), .A4(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n873));
  NAND2_X1  g448(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT95), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n872), .B2(new_n873), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n760), .A2(KEYINPUT23), .A3(G20), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT23), .ZN(new_n879));
  INV_X1    g454(.A(G20), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(G16), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n878), .B(new_n881), .C1(new_n620), .C2(new_n760), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G1956), .ZN(new_n883));
  NOR4_X1   g458(.A1(new_n830), .A2(new_n876), .A3(new_n877), .A4(new_n883), .ZN(G311));
  NOR2_X1   g459(.A1(new_n830), .A2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n876), .A2(new_n877), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(G150));
  AOI22_X1  g462(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n888), .A2(KEYINPUT101), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(KEYINPUT101), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(G651), .A3(new_n890), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n525), .A2(G93), .B1(new_n527), .B2(G55), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G860), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT37), .Z(new_n895));
  NOR2_X1   g470(.A1(new_n615), .A2(new_n623), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n548), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n547), .A2(new_n891), .A3(new_n892), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n898), .B(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT102), .ZN(new_n906));
  INV_X1    g481(.A(G860), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n895), .B1(new_n906), .B2(new_n908), .ZN(G145));
  XOR2_X1   g484(.A(new_n858), .B(new_n642), .Z(new_n910));
  NAND2_X1  g485(.A1(new_n481), .A2(G130), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n634), .A2(G142), .ZN(new_n912));
  OR2_X1    g487(.A1(G106), .A2(G2105), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n913), .B(G2104), .C1(G118), .C2(new_n474), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n910), .B(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n491), .A2(KEYINPUT103), .A3(new_n495), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n919));
  INV_X1    g494(.A(new_n484), .ZN(new_n920));
  INV_X1    g495(.A(G126), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n462), .B2(new_n464), .ZN(new_n922));
  INV_X1    g497(.A(new_n488), .ZN(new_n923));
  OAI21_X1  g498(.A(G2105), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n920), .B1(new_n924), .B2(KEYINPUT4), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n919), .B1(new_n925), .B2(new_n494), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n918), .A2(new_n926), .A3(new_n816), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n816), .B1(new_n918), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n774), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n929), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n769), .A2(new_n773), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n927), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n797), .A2(KEYINPUT104), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n930), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n797), .A2(KEYINPUT104), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n930), .A2(new_n933), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n917), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n934), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n910), .B(new_n915), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n930), .A2(new_n933), .A3(new_n934), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n638), .B(new_n472), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(G162), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G37), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n938), .A2(new_n944), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g528(.A(G290), .B(G288), .ZN(new_n954));
  XNOR2_X1  g529(.A(G303), .B(G305), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n954), .B(new_n955), .Z(new_n956));
  NAND2_X1  g531(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n629), .A2(new_n901), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n627), .A2(new_n628), .A3(new_n902), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n566), .B(new_n611), .C1(new_n580), .C2(new_n581), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n577), .A2(KEYINPUT74), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n577), .A2(KEYINPUT74), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n567), .A2(new_n570), .A3(KEYINPUT9), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n570), .B1(new_n567), .B2(KEYINPUT9), .ZN(new_n966));
  OAI22_X1  g541(.A1(new_n963), .A2(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT75), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n572), .A2(new_n579), .A3(new_n573), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n611), .B1(new_n970), .B2(new_n566), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n962), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(KEYINPUT105), .ZN(new_n973));
  INV_X1    g548(.A(new_n611), .ZN(new_n974));
  NAND2_X1  g549(.A1(G299), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n961), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n959), .B(new_n960), .C1(new_n973), .C2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n959), .A2(new_n960), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT41), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n975), .B2(new_n961), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n961), .A2(new_n982), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n981), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n972), .A2(KEYINPUT41), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n958), .A2(new_n979), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n958), .B1(new_n979), .B2(new_n988), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n990), .A2(new_n991), .B1(KEYINPUT107), .B2(KEYINPUT42), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n979), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n957), .A3(new_n956), .ZN(new_n994));
  NOR2_X1   g569(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n995), .A3(new_n989), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(G868), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G868), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT108), .B1(new_n893), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n992), .A2(KEYINPUT108), .A3(new_n996), .A4(G868), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(G295));
  AND2_X1   g577(.A1(new_n1000), .A2(new_n1001), .ZN(G331));
  AND3_X1   g578(.A1(new_n899), .A2(G286), .A3(new_n900), .ZN(new_n1004));
  AOI21_X1  g579(.A(G286), .B1(new_n899), .B2(new_n900), .ZN(new_n1005));
  OAI21_X1  g580(.A(G301), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n901), .A2(G168), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n899), .A2(G286), .A3(new_n900), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(G171), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(new_n972), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n986), .A2(new_n987), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(new_n1010), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n954), .B(new_n955), .ZN(new_n1014));
  AOI21_X1  g589(.A(G37), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n976), .A2(new_n981), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT106), .B1(new_n962), .B2(new_n971), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n984), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1010), .B(new_n1016), .C1(new_n1018), .C2(new_n981), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n973), .B2(new_n978), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n956), .A3(new_n1021), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1015), .A2(KEYINPUT43), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n986), .B2(new_n987), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n956), .B1(new_n1024), .B2(new_n1011), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT43), .B1(new_n1015), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT44), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1011), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n976), .A2(new_n981), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n1018), .B2(new_n981), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1014), .B(new_n1028), .C1(new_n1030), .C2(new_n1020), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1025), .A2(new_n1031), .A3(new_n950), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT43), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT43), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1031), .A2(new_n1022), .A3(new_n1034), .A4(new_n950), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1027), .B1(new_n1037), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g613(.A(G1996), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n932), .B(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n816), .B(G2067), .Z(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n858), .A2(new_n864), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n1042), .A2(new_n1043), .B1(G2067), .B2(new_n816), .ZN(new_n1044));
  INV_X1    g619(.A(G1384), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT103), .B1(new_n491), .B2(new_n495), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n925), .A2(new_n919), .A3(new_n494), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g623(.A(new_n1048), .B(KEYINPUT109), .Z(new_n1049));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1044), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G290), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n870), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n1058), .B(new_n1059), .Z(new_n1060));
  AOI21_X1  g635(.A(new_n1042), .B1(new_n864), .B2(new_n858), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1053), .B1(new_n1061), .B2(new_n1043), .ZN(new_n1062));
  NAND2_X1  g637(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1041), .A2(new_n774), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1063), .B1(new_n1053), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1054), .A2(new_n1039), .A3(new_n1067), .ZN(new_n1068));
  OAI22_X1  g643(.A1(new_n1053), .A2(G1996), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT47), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI221_X1 g648(.A(new_n1055), .B1(new_n1060), .B2(new_n1062), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1045), .B1(new_n925), .B2(new_n494), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT110), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT110), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n1045), .C1(new_n925), .C2(new_n494), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1050), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G2078), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1384), .B1(new_n491), .B2(new_n495), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1051), .B1(new_n1082), .B2(KEYINPUT45), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT122), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1080), .A2(new_n1086), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(KEYINPUT53), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1961), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1078), .B1(new_n496), .B2(new_n1045), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1079), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1052), .B1(new_n1082), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT45), .B(new_n1045), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1076), .A2(new_n1050), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(new_n1081), .A3(new_n1052), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1089), .A2(new_n1098), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1088), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G171), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1052), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G305), .A2(G1981), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n588), .A2(new_n589), .A3(new_n847), .A4(new_n590), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT49), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(KEYINPUT49), .A3(new_n1112), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1110), .A2(new_n1115), .A3(G8), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1976), .ZN(new_n1118));
  NOR2_X1   g693(.A1(G288), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT52), .B1(G288), .B2(new_n1118), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1110), .A2(G8), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1051), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1123));
  INV_X1    g698(.A(G8), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n1119), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1117), .B(new_n1122), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1128), .A2(KEYINPUT112), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT55), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(G166), .B2(new_n1124), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(KEYINPUT112), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1051), .B1(new_n1076), .B2(new_n1050), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1099), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1971), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G2090), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1094), .A2(new_n1138), .A3(new_n1097), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1124), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1127), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1133), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1095), .B(new_n1045), .C1(new_n925), .C2(new_n494), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT113), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1077), .A2(new_n1079), .A3(new_n1090), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1138), .A3(new_n1052), .A4(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1146), .A2(new_n1137), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1142), .B1(new_n1147), .B2(new_n1124), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1141), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1090), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT114), .B(G2084), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1150), .A2(new_n1096), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(G1966), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1154));
  OAI21_X1  g729(.A(G286), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n805), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1094), .A2(new_n1097), .A3(new_n1151), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(new_n1158), .A3(G168), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1155), .A2(new_n1159), .A3(G8), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT51), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT51), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1162), .A3(G8), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1161), .A2(KEYINPUT62), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT62), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1109), .B(new_n1149), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(G288), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1117), .A2(new_n1118), .A3(new_n1167), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n1124), .B(new_n1123), .C1(new_n1168), .C2(new_n1112), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1140), .A2(new_n1133), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(new_n1127), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1127), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1124), .B(G286), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1148), .A2(new_n1170), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(KEYINPUT115), .B(KEYINPUT63), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1173), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT63), .B1(new_n1140), .B2(new_n1133), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT116), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1179), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT116), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(new_n1141), .A3(new_n1182), .A4(new_n1174), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1177), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1166), .A2(new_n1172), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1149), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT119), .ZN(new_n1188));
  XNOR2_X1  g763(.A(KEYINPUT58), .B(G1341), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1110), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(KEYINPUT119), .B1(new_n1123), .B2(new_n1189), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1099), .A2(new_n1039), .A3(new_n1134), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT59), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1194), .A2(new_n1195), .A3(new_n548), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT121), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1194), .A2(new_n548), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT120), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT120), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1199), .A2(new_n1203), .A3(KEYINPUT59), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1198), .A2(new_n1201), .A3(new_n1202), .A4(new_n1204), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1144), .A2(new_n1052), .A3(new_n1145), .ZN(new_n1206));
  INV_X1    g781(.A(G1956), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(KEYINPUT56), .B(G2072), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1099), .A2(new_n1134), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(KEYINPUT57), .B1(new_n572), .B2(new_n579), .ZN(new_n1211));
  AOI22_X1  g786(.A1(G299), .A2(KEYINPUT57), .B1(new_n1211), .B2(new_n566), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1208), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  AND2_X1   g788(.A1(new_n1213), .A2(KEYINPUT61), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1215), .A2(KEYINPUT118), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT118), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1217), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1214), .B1(new_n1219), .B2(new_n1212), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1212), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1215), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g797(.A(KEYINPUT61), .B1(new_n1222), .B2(new_n1213), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1150), .A2(new_n1096), .ZN(new_n1226));
  OAI221_X1 g801(.A(new_n1225), .B1(G2067), .B2(new_n1110), .C1(new_n1226), .C2(G1348), .ZN(new_n1227));
  OAI22_X1  g802(.A1(new_n1226), .A2(G1348), .B1(G2067), .B2(new_n1110), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1228), .A2(KEYINPUT60), .A3(new_n616), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1224), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1223), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1205), .A2(new_n1220), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1219), .A2(new_n1212), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1228), .A2(new_n616), .ZN(new_n1234));
  XNOR2_X1  g809(.A(new_n1234), .B(KEYINPUT117), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1213), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1187), .B1(new_n1232), .B2(new_n1236), .ZN(new_n1237));
  OR3_X1    g812(.A1(new_n1104), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1238));
  OAI21_X1  g813(.A(KEYINPUT124), .B1(new_n1104), .B2(G171), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1241));
  AND3_X1   g816(.A1(new_n1099), .A2(new_n1081), .A3(new_n1052), .ZN(new_n1242));
  NAND3_X1  g817(.A1(new_n1241), .A2(KEYINPUT53), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g818(.A(G301), .B1(new_n1243), .B2(new_n1103), .ZN(new_n1244));
  OAI21_X1  g819(.A(KEYINPUT54), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1245));
  AND2_X1   g820(.A1(new_n1103), .A2(G301), .ZN(new_n1246));
  AOI21_X1  g821(.A(KEYINPUT54), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1247), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g824(.A(new_n1185), .B1(new_n1237), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1061), .A2(new_n1043), .ZN(new_n1251));
  AOI21_X1  g826(.A(new_n1251), .B1(G1986), .B2(G290), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1053), .B1(new_n1252), .B2(new_n1057), .ZN(new_n1253));
  OAI21_X1  g828(.A(new_n1075), .B1(new_n1250), .B2(new_n1253), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1256));
  NOR2_X1   g830(.A1(G229), .A2(G227), .ZN(new_n1257));
  AND3_X1   g831(.A1(new_n687), .A2(new_n1257), .A3(G319), .ZN(new_n1258));
  NAND2_X1  g832(.A1(new_n1258), .A2(new_n952), .ZN(new_n1259));
  INV_X1    g833(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g834(.A(new_n1256), .B1(new_n1036), .B2(new_n1260), .ZN(new_n1261));
  AOI211_X1 g835(.A(KEYINPUT127), .B(new_n1259), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1262));
  NOR2_X1   g836(.A1(new_n1261), .A2(new_n1262), .ZN(G308));
  AOI21_X1  g837(.A(new_n1034), .B1(new_n1015), .B2(new_n1025), .ZN(new_n1264));
  INV_X1    g838(.A(new_n1035), .ZN(new_n1265));
  OAI21_X1  g839(.A(new_n1260), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g840(.A1(new_n1266), .A2(KEYINPUT127), .ZN(new_n1267));
  NAND3_X1  g841(.A1(new_n1036), .A2(new_n1256), .A3(new_n1260), .ZN(new_n1268));
  NAND2_X1  g842(.A1(new_n1267), .A2(new_n1268), .ZN(G225));
endmodule


