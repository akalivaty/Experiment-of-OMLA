

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732;

  XNOR2_X1 U371 ( .A(n361), .B(G107), .ZN(n493) );
  AND2_X1 U372 ( .A1(n652), .A2(n535), .ZN(n426) );
  INV_X1 U373 ( .A(G953), .ZN(n721) );
  NOR2_X1 U374 ( .A1(n609), .A2(n698), .ZN(n610) );
  XNOR2_X2 U375 ( .A(n436), .B(KEYINPUT0), .ZN(n529) );
  NOR2_X2 U376 ( .A1(n727), .A2(n731), .ZN(n365) );
  XNOR2_X2 U377 ( .A(KEYINPUT42), .B(n558), .ZN(n727) );
  XNOR2_X2 U378 ( .A(n426), .B(n425), .ZN(n571) );
  XNOR2_X2 U379 ( .A(KEYINPUT38), .B(n536), .ZN(n653) );
  XOR2_X2 U380 ( .A(n452), .B(n451), .Z(n551) );
  NOR2_X1 U381 ( .A1(n659), .A2(n656), .ZN(n364) );
  BUF_X1 U382 ( .A(n535), .Z(n594) );
  NAND2_X1 U383 ( .A1(n523), .A2(n522), .ZN(n630) );
  NAND2_X1 U384 ( .A1(n702), .A2(n714), .ZN(n670) );
  XNOR2_X1 U385 ( .A(n510), .B(KEYINPUT22), .ZN(n515) );
  XNOR2_X1 U386 ( .A(n364), .B(KEYINPUT41), .ZN(n667) );
  XNOR2_X1 U387 ( .A(n424), .B(n423), .ZN(n535) );
  XNOR2_X1 U388 ( .A(n403), .B(n402), .ZN(n666) );
  XNOR2_X1 U389 ( .A(n370), .B(G110), .ZN(n445) );
  XNOR2_X1 U390 ( .A(G146), .B(G125), .ZN(n444) );
  XNOR2_X1 U391 ( .A(n453), .B(n396), .ZN(n466) );
  XNOR2_X1 U392 ( .A(G134), .B(G131), .ZN(n396) );
  XNOR2_X1 U393 ( .A(n492), .B(KEYINPUT4), .ZN(n453) );
  AND2_X1 U394 ( .A1(n714), .A2(n391), .ZN(n389) );
  NAND2_X1 U395 ( .A1(n394), .A2(n392), .ZN(n391) );
  NAND2_X1 U396 ( .A1(n393), .A2(n603), .ZN(n392) );
  NAND2_X1 U397 ( .A1(n350), .A2(KEYINPUT71), .ZN(n394) );
  NAND2_X1 U398 ( .A1(n384), .A2(n383), .ZN(n534) );
  NOR2_X1 U399 ( .A1(n617), .A2(n351), .ZN(n383) );
  XNOR2_X1 U400 ( .A(n386), .B(n385), .ZN(n384) );
  XNOR2_X1 U401 ( .A(KEYINPUT10), .B(n444), .ZN(n712) );
  NOR2_X1 U402 ( .A1(G953), .A2(G237), .ZN(n481) );
  INV_X1 U403 ( .A(KEYINPUT51), .ZN(n379) );
  NOR2_X1 U404 ( .A1(n650), .A2(n379), .ZN(n378) );
  INV_X1 U405 ( .A(G116), .ZN(n361) );
  NAND2_X1 U406 ( .A1(n653), .A2(n652), .ZN(n659) );
  XNOR2_X1 U407 ( .A(n463), .B(G472), .ZN(n553) );
  XNOR2_X1 U408 ( .A(n448), .B(n369), .ZN(n368) );
  XNOR2_X1 U409 ( .A(n445), .B(KEYINPUT24), .ZN(n369) );
  XNOR2_X1 U410 ( .A(n447), .B(n446), .ZN(n499) );
  XNOR2_X1 U411 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n446) );
  XNOR2_X1 U412 ( .A(n363), .B(n486), .ZN(n684) );
  XNOR2_X1 U413 ( .A(n487), .B(n353), .ZN(n363) );
  XNOR2_X1 U414 ( .A(n466), .B(n465), .ZN(n713) );
  XOR2_X1 U415 ( .A(G101), .B(G104), .Z(n468) );
  XOR2_X1 U416 ( .A(KEYINPUT73), .B(G107), .Z(n471) );
  INV_X1 U417 ( .A(KEYINPUT65), .ZN(n397) );
  INV_X1 U418 ( .A(KEYINPUT85), .ZN(n402) );
  NAND2_X1 U419 ( .A1(n430), .A2(G952), .ZN(n403) );
  XNOR2_X1 U420 ( .A(n381), .B(n380), .ZN(n664) );
  OR2_X2 U421 ( .A1(n529), .A2(n509), .ZN(n510) );
  OR2_X1 U422 ( .A1(n678), .A2(G902), .ZN(n474) );
  NOR2_X1 U423 ( .A1(n515), .A2(n644), .ZN(n520) );
  XNOR2_X1 U424 ( .A(KEYINPUT6), .B(n553), .ZN(n562) );
  NOR2_X1 U425 ( .A1(G952), .A2(n721), .ZN(n698) );
  XNOR2_X1 U426 ( .A(n382), .B(KEYINPUT49), .ZN(n641) );
  NAND2_X1 U427 ( .A1(n519), .A2(n507), .ZN(n382) );
  INV_X1 U428 ( .A(n602), .ZN(n393) );
  OR2_X1 U429 ( .A1(G237), .A2(G902), .ZN(n420) );
  XNOR2_X1 U430 ( .A(n438), .B(n366), .ZN(n440) );
  XNOR2_X1 U431 ( .A(KEYINPUT20), .B(KEYINPUT88), .ZN(n366) );
  XOR2_X1 U432 ( .A(KEYINPUT5), .B(G137), .Z(n458) );
  XNOR2_X1 U433 ( .A(G116), .B(G119), .ZN(n454) );
  XOR2_X1 U434 ( .A(KEYINPUT70), .B(G146), .Z(n455) );
  XNOR2_X1 U435 ( .A(G101), .B(KEYINPUT3), .ZN(n409) );
  XNOR2_X1 U436 ( .A(n408), .B(n407), .ZN(n412) );
  XNOR2_X1 U437 ( .A(n493), .B(n406), .ZN(n408) );
  XNOR2_X1 U438 ( .A(KEYINPUT68), .B(KEYINPUT16), .ZN(n406) );
  INV_X1 U439 ( .A(KEYINPUT44), .ZN(n385) );
  INV_X1 U440 ( .A(G119), .ZN(n370) );
  XOR2_X1 U441 ( .A(G122), .B(G104), .Z(n485) );
  XNOR2_X1 U442 ( .A(G113), .B(G143), .ZN(n479) );
  XOR2_X1 U443 ( .A(KEYINPUT11), .B(KEYINPUT92), .Z(n483) );
  XOR2_X1 U444 ( .A(G137), .B(G140), .Z(n464) );
  XNOR2_X1 U445 ( .A(n428), .B(n404), .ZN(n430) );
  XNOR2_X1 U446 ( .A(n427), .B(KEYINPUT69), .ZN(n404) );
  NAND2_X1 U447 ( .A1(G234), .A2(G237), .ZN(n427) );
  NAND2_X1 U448 ( .A1(n376), .A2(n375), .ZN(n381) );
  AND2_X1 U449 ( .A1(n377), .A2(n358), .ZN(n376) );
  INV_X1 U450 ( .A(KEYINPUT112), .ZN(n380) );
  XNOR2_X1 U451 ( .A(KEYINPUT19), .B(KEYINPUT72), .ZN(n425) );
  NOR2_X1 U452 ( .A1(n729), .A2(n598), .ZN(n599) );
  XOR2_X1 U453 ( .A(KEYINPUT93), .B(KEYINPUT9), .Z(n491) );
  XNOR2_X1 U454 ( .A(G134), .B(G122), .ZN(n490) );
  XOR2_X1 U455 ( .A(KEYINPUT7), .B(KEYINPUT94), .Z(n496) );
  XNOR2_X1 U456 ( .A(n453), .B(n355), .ZN(n417) );
  NOR2_X1 U457 ( .A1(n571), .A2(n570), .ZN(n580) );
  XNOR2_X1 U458 ( .A(n489), .B(n488), .ZN(n523) );
  XNOR2_X1 U459 ( .A(n368), .B(n367), .ZN(n449) );
  AND2_X1 U460 ( .A1(n499), .A2(G221), .ZN(n367) );
  BUF_X1 U461 ( .A(n682), .Z(n694) );
  XNOR2_X1 U462 ( .A(G146), .B(G110), .ZN(n470) );
  AND2_X1 U463 ( .A1(n672), .A2(n354), .ZN(n372) );
  NOR2_X1 U464 ( .A1(n667), .A2(n570), .ZN(n558) );
  NAND2_X1 U465 ( .A1(n399), .A2(n644), .ZN(n636) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n399) );
  XNOR2_X1 U467 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n400) );
  XNOR2_X1 U468 ( .A(KEYINPUT90), .B(n526), .ZN(n619) );
  NOR2_X1 U469 ( .A1(n642), .A2(n529), .ZN(n524) );
  NOR2_X1 U470 ( .A1(n521), .A2(n562), .ZN(n617) );
  AND2_X1 U471 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U472 ( .A1(KEYINPUT2), .A2(n601), .ZN(n350) );
  AND2_X1 U473 ( .A1(n533), .A2(n532), .ZN(n351) );
  AND2_X1 U474 ( .A1(n520), .A2(n512), .ZN(n352) );
  XOR2_X1 U475 ( .A(n480), .B(n479), .Z(n353) );
  OR2_X1 U476 ( .A1(n668), .A2(n667), .ZN(n354) );
  XOR2_X1 U477 ( .A(n443), .B(n416), .Z(n355) );
  XOR2_X1 U478 ( .A(n665), .B(KEYINPUT52), .Z(n356) );
  AND2_X1 U479 ( .A1(n650), .A2(n379), .ZN(n357) );
  NOR2_X1 U480 ( .A1(n667), .A2(n378), .ZN(n358) );
  XOR2_X1 U481 ( .A(KEYINPUT15), .B(G902), .Z(n603) );
  XOR2_X1 U482 ( .A(n607), .B(n606), .Z(n359) );
  AND2_X1 U483 ( .A1(n350), .A2(n398), .ZN(n360) );
  NAND2_X1 U484 ( .A1(n670), .A2(n360), .ZN(n388) );
  NAND2_X1 U485 ( .A1(n362), .A2(n503), .ZN(n504) );
  XNOR2_X1 U486 ( .A(n478), .B(KEYINPUT34), .ZN(n362) );
  INV_X1 U487 ( .A(n444), .ZN(n443) );
  NAND2_X1 U488 ( .A1(n565), .A2(n594), .ZN(n401) );
  NAND2_X1 U489 ( .A1(n412), .A2(n413), .ZN(n414) );
  XNOR2_X1 U490 ( .A(n365), .B(n559), .ZN(n587) );
  NOR2_X1 U491 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U492 ( .A1(n371), .A2(n673), .ZN(n674) );
  NAND2_X1 U493 ( .A1(n373), .A2(n372), .ZN(n371) );
  NAND2_X1 U494 ( .A1(n356), .A2(n374), .ZN(n373) );
  INV_X1 U495 ( .A(n666), .ZN(n374) );
  OR2_X1 U496 ( .A1(n651), .A2(n379), .ZN(n375) );
  NAND2_X1 U497 ( .A1(n651), .A2(n357), .ZN(n377) );
  INV_X1 U498 ( .A(n519), .ZN(n640) );
  XNOR2_X1 U499 ( .A(n551), .B(KEYINPUT96), .ZN(n519) );
  NAND2_X1 U500 ( .A1(n730), .A2(n387), .ZN(n386) );
  NOR2_X1 U501 ( .A1(n352), .A2(n728), .ZN(n387) );
  XNOR2_X2 U502 ( .A(n518), .B(KEYINPUT32), .ZN(n730) );
  NAND2_X1 U503 ( .A1(n390), .A2(n388), .ZN(n395) );
  NAND2_X1 U504 ( .A1(n389), .A2(n702), .ZN(n390) );
  XNOR2_X2 U505 ( .A(G143), .B(G128), .ZN(n492) );
  XNOR2_X2 U506 ( .A(n534), .B(KEYINPUT45), .ZN(n702) );
  NOR2_X1 U507 ( .A1(n670), .A2(n602), .ZN(n673) );
  XNOR2_X2 U508 ( .A(n395), .B(n397), .ZN(n682) );
  INV_X1 U509 ( .A(KEYINPUT71), .ZN(n398) );
  XNOR2_X1 U510 ( .A(n608), .B(n359), .ZN(n609) );
  AND2_X2 U511 ( .A1(n600), .A2(n599), .ZN(n714) );
  NAND2_X1 U512 ( .A1(n435), .A2(n434), .ZN(n436) );
  INV_X1 U513 ( .A(n485), .ZN(n407) );
  XNOR2_X1 U514 ( .A(KEYINPUT98), .B(KEYINPUT33), .ZN(n476) );
  INV_X1 U515 ( .A(n732), .ZN(n598) );
  INV_X1 U516 ( .A(n464), .ZN(n465) );
  NAND2_X1 U517 ( .A1(n508), .A2(n639), .ZN(n509) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U519 ( .A(KEYINPUT82), .ZN(n421) );
  XNOR2_X1 U520 ( .A(n462), .B(n461), .ZN(n611) );
  BUF_X1 U521 ( .A(n705), .Z(n706) );
  XNOR2_X1 U522 ( .A(n713), .B(n469), .ZN(n473) );
  XNOR2_X1 U523 ( .A(n422), .B(n421), .ZN(n423) );
  INV_X1 U524 ( .A(n551), .ZN(n511) );
  XNOR2_X1 U525 ( .A(n450), .B(n449), .ZN(n693) );
  XNOR2_X1 U526 ( .A(n684), .B(n683), .ZN(n685) );
  INV_X1 U527 ( .A(n567), .ZN(n503) );
  NOR2_X1 U528 ( .A1(n642), .A2(n511), .ZN(n512) );
  XNOR2_X1 U529 ( .A(n504), .B(KEYINPUT35), .ZN(n728) );
  NAND2_X1 U530 ( .A1(G214), .A2(n420), .ZN(n405) );
  XOR2_X1 U531 ( .A(KEYINPUT83), .B(n405), .Z(n652) );
  INV_X1 U532 ( .A(n412), .ZN(n411) );
  XNOR2_X1 U533 ( .A(n409), .B(G113), .ZN(n459) );
  XNOR2_X1 U534 ( .A(n459), .B(n445), .ZN(n413) );
  INV_X1 U535 ( .A(n413), .ZN(n410) );
  NAND2_X1 U536 ( .A1(n411), .A2(n410), .ZN(n415) );
  NAND2_X1 U537 ( .A1(n415), .A2(n414), .ZN(n705) );
  XNOR2_X1 U538 ( .A(n705), .B(KEYINPUT17), .ZN(n419) );
  NAND2_X1 U539 ( .A1(G224), .A2(n721), .ZN(n416) );
  XOR2_X1 U540 ( .A(n417), .B(KEYINPUT18), .Z(n418) );
  XNOR2_X1 U541 ( .A(n418), .B(n419), .ZN(n604) );
  INV_X1 U542 ( .A(n603), .ZN(n437) );
  NAND2_X1 U543 ( .A1(n604), .A2(n437), .ZN(n424) );
  NAND2_X1 U544 ( .A1(G210), .A2(n420), .ZN(n422) );
  INV_X1 U545 ( .A(n571), .ZN(n435) );
  XOR2_X1 U546 ( .A(KEYINPUT84), .B(KEYINPUT14), .Z(n428) );
  AND2_X1 U547 ( .A1(n430), .A2(G953), .ZN(n429) );
  NAND2_X1 U548 ( .A1(G902), .A2(n429), .ZN(n540) );
  NOR2_X1 U549 ( .A1(G898), .A2(n540), .ZN(n432) );
  NOR2_X1 U550 ( .A1(n666), .A2(G953), .ZN(n431) );
  XNOR2_X1 U551 ( .A(n431), .B(KEYINPUT86), .ZN(n541) );
  NOR2_X1 U552 ( .A1(n432), .A2(n541), .ZN(n433) );
  XNOR2_X1 U553 ( .A(KEYINPUT87), .B(n433), .ZN(n434) );
  NAND2_X1 U554 ( .A1(n437), .A2(G234), .ZN(n438) );
  NAND2_X1 U555 ( .A1(n440), .A2(G221), .ZN(n439) );
  XOR2_X1 U556 ( .A(KEYINPUT21), .B(n439), .Z(n639) );
  INV_X1 U557 ( .A(n639), .ZN(n507) );
  XOR2_X1 U558 ( .A(KEYINPUT89), .B(KEYINPUT25), .Z(n442) );
  NAND2_X1 U559 ( .A1(G217), .A2(n440), .ZN(n441) );
  XNOR2_X1 U560 ( .A(n442), .B(n441), .ZN(n452) );
  XOR2_X1 U561 ( .A(KEYINPUT23), .B(n712), .Z(n450) );
  NAND2_X1 U562 ( .A1(n721), .A2(G234), .ZN(n447) );
  XNOR2_X1 U563 ( .A(G128), .B(n464), .ZN(n448) );
  NOR2_X1 U564 ( .A1(G902), .A2(n693), .ZN(n451) );
  NOR2_X1 U565 ( .A1(n507), .A2(n551), .ZN(n645) );
  XNOR2_X1 U566 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U567 ( .A(n466), .B(n456), .ZN(n462) );
  NAND2_X1 U568 ( .A1(n481), .A2(G210), .ZN(n457) );
  XNOR2_X1 U569 ( .A(n458), .B(n457), .ZN(n460) );
  NOR2_X1 U570 ( .A1(n611), .A2(G902), .ZN(n463) );
  AND2_X1 U571 ( .A1(n645), .A2(n562), .ZN(n475) );
  NAND2_X1 U572 ( .A1(G227), .A2(n721), .ZN(n467) );
  XNOR2_X1 U573 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U574 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U575 ( .A(n473), .B(n472), .ZN(n678) );
  XNOR2_X2 U576 ( .A(n474), .B(G469), .ZN(n557) );
  XNOR2_X1 U577 ( .A(n557), .B(KEYINPUT1), .ZN(n527) );
  AND2_X1 U578 ( .A1(n475), .A2(n527), .ZN(n477) );
  XNOR2_X1 U579 ( .A(n477), .B(n476), .ZN(n668) );
  NOR2_X1 U580 ( .A1(n529), .A2(n668), .ZN(n478) );
  XNOR2_X1 U581 ( .A(KEYINPUT13), .B(G475), .ZN(n489) );
  XOR2_X1 U582 ( .A(G140), .B(G131), .Z(n480) );
  NAND2_X1 U583 ( .A1(G214), .A2(n481), .ZN(n482) );
  XNOR2_X1 U584 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U585 ( .A(n484), .B(KEYINPUT12), .Z(n487) );
  XNOR2_X1 U586 ( .A(n485), .B(n712), .ZN(n486) );
  NOR2_X1 U587 ( .A1(G902), .A2(n684), .ZN(n488) );
  XNOR2_X1 U588 ( .A(n491), .B(n490), .ZN(n498) );
  INV_X1 U589 ( .A(n492), .ZN(n494) );
  XNOR2_X1 U590 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U591 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U592 ( .A(n498), .B(n497), .Z(n501) );
  NAND2_X1 U593 ( .A1(G217), .A2(n499), .ZN(n500) );
  XNOR2_X1 U594 ( .A(n501), .B(n500), .ZN(n691) );
  NOR2_X1 U595 ( .A1(G902), .A2(n691), .ZN(n502) );
  XNOR2_X1 U596 ( .A(G478), .B(n502), .ZN(n522) );
  INV_X1 U597 ( .A(n522), .ZN(n505) );
  NAND2_X1 U598 ( .A1(n523), .A2(n505), .ZN(n567) );
  NOR2_X1 U599 ( .A1(n505), .A2(n523), .ZN(n506) );
  XNOR2_X1 U600 ( .A(n506), .B(KEYINPUT95), .ZN(n656) );
  INV_X1 U601 ( .A(n656), .ZN(n508) );
  BUF_X1 U602 ( .A(n527), .Z(n644) );
  INV_X1 U603 ( .A(n553), .ZN(n642) );
  XOR2_X1 U604 ( .A(n562), .B(KEYINPUT74), .Z(n517) );
  NAND2_X1 U605 ( .A1(n519), .A2(n644), .ZN(n513) );
  XOR2_X1 U606 ( .A(KEYINPUT97), .B(n513), .Z(n514) );
  NOR2_X1 U607 ( .A1(n515), .A2(n514), .ZN(n516) );
  NAND2_X1 U608 ( .A1(n517), .A2(n516), .ZN(n518) );
  NAND2_X1 U609 ( .A1(n640), .A2(n520), .ZN(n521) );
  NOR2_X1 U610 ( .A1(n523), .A2(n522), .ZN(n581) );
  INV_X1 U611 ( .A(n581), .ZN(n633) );
  NAND2_X1 U612 ( .A1(n630), .A2(n633), .ZN(n533) );
  AND2_X1 U613 ( .A1(n557), .A2(n645), .ZN(n525) );
  NAND2_X1 U614 ( .A1(n525), .A2(n524), .ZN(n526) );
  AND2_X1 U615 ( .A1(n645), .A2(n527), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n642), .A2(n528), .ZN(n650) );
  NOR2_X1 U617 ( .A1(n650), .A2(n529), .ZN(n531) );
  XOR2_X1 U618 ( .A(KEYINPUT91), .B(KEYINPUT31), .Z(n530) );
  XNOR2_X1 U619 ( .A(n531), .B(n530), .ZN(n632) );
  NAND2_X1 U620 ( .A1(n619), .A2(n632), .ZN(n532) );
  INV_X1 U621 ( .A(n594), .ZN(n536) );
  INV_X1 U622 ( .A(n652), .ZN(n537) );
  NOR2_X1 U623 ( .A1(n537), .A2(n553), .ZN(n539) );
  XNOR2_X1 U624 ( .A(KEYINPUT101), .B(KEYINPUT30), .ZN(n538) );
  XNOR2_X1 U625 ( .A(n539), .B(n538), .ZN(n547) );
  NOR2_X1 U626 ( .A1(G900), .A2(n540), .ZN(n542) );
  NOR2_X1 U627 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U628 ( .A(n543), .B(KEYINPUT75), .ZN(n544) );
  NAND2_X1 U629 ( .A1(n544), .A2(n639), .ZN(n550) );
  NOR2_X1 U630 ( .A1(n551), .A2(n550), .ZN(n545) );
  NAND2_X1 U631 ( .A1(n557), .A2(n545), .ZN(n546) );
  NOR2_X1 U632 ( .A1(n547), .A2(n546), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n653), .A2(n566), .ZN(n548) );
  XOR2_X1 U634 ( .A(n548), .B(KEYINPUT39), .Z(n596) );
  NOR2_X1 U635 ( .A1(n630), .A2(n596), .ZN(n549) );
  XNOR2_X1 U636 ( .A(n549), .B(KEYINPUT40), .ZN(n731) );
  XOR2_X1 U637 ( .A(KEYINPUT28), .B(KEYINPUT102), .Z(n555) );
  XNOR2_X1 U638 ( .A(KEYINPUT67), .B(n550), .ZN(n552) );
  NAND2_X1 U639 ( .A1(n552), .A2(n551), .ZN(n560) );
  NOR2_X1 U640 ( .A1(n553), .A2(n560), .ZN(n554) );
  XOR2_X1 U641 ( .A(n555), .B(n554), .Z(n556) );
  NAND2_X1 U642 ( .A1(n557), .A2(n556), .ZN(n570) );
  XNOR2_X1 U643 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n559) );
  NOR2_X1 U644 ( .A1(n630), .A2(n560), .ZN(n561) );
  NAND2_X1 U645 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U646 ( .A(n563), .B(KEYINPUT99), .ZN(n564) );
  NAND2_X1 U647 ( .A1(n564), .A2(n652), .ZN(n591) );
  INV_X1 U648 ( .A(n591), .ZN(n565) );
  XNOR2_X1 U649 ( .A(n636), .B(KEYINPUT80), .ZN(n578) );
  INV_X1 U650 ( .A(n566), .ZN(n568) );
  NOR2_X1 U651 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U652 ( .A1(n569), .A2(n594), .ZN(n628) );
  AND2_X1 U653 ( .A1(n633), .A2(n630), .ZN(n658) );
  NAND2_X1 U654 ( .A1(n658), .A2(KEYINPUT76), .ZN(n572) );
  NAND2_X1 U655 ( .A1(n572), .A2(n580), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n573), .A2(KEYINPUT47), .ZN(n574) );
  NAND2_X1 U657 ( .A1(n628), .A2(n574), .ZN(n576) );
  NOR2_X1 U658 ( .A1(KEYINPUT76), .A2(n658), .ZN(n575) );
  NOR2_X1 U659 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U660 ( .A1(n578), .A2(n577), .ZN(n585) );
  INV_X1 U661 ( .A(n580), .ZN(n579) );
  NOR2_X1 U662 ( .A1(n630), .A2(n579), .ZN(n629) );
  NAND2_X1 U663 ( .A1(n581), .A2(n580), .ZN(n625) );
  NAND2_X1 U664 ( .A1(KEYINPUT76), .A2(n625), .ZN(n582) );
  NOR2_X1 U665 ( .A1(n629), .A2(n582), .ZN(n583) );
  NOR2_X1 U666 ( .A1(KEYINPUT47), .A2(n583), .ZN(n584) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(n590) );
  XNOR2_X1 U668 ( .A(KEYINPUT48), .B(KEYINPUT66), .ZN(n588) );
  XNOR2_X1 U669 ( .A(n588), .B(KEYINPUT79), .ZN(n589) );
  XNOR2_X1 U670 ( .A(n590), .B(n589), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n644), .A2(n591), .ZN(n592) );
  XNOR2_X1 U672 ( .A(n592), .B(KEYINPUT43), .ZN(n593) );
  NOR2_X1 U673 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U674 ( .A(KEYINPUT100), .B(n595), .ZN(n729) );
  OR2_X1 U675 ( .A1(n633), .A2(n596), .ZN(n597) );
  XNOR2_X1 U676 ( .A(n597), .B(KEYINPUT104), .ZN(n732) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT78), .ZN(n601) );
  XOR2_X1 U678 ( .A(KEYINPUT2), .B(KEYINPUT71), .Z(n602) );
  NAND2_X1 U679 ( .A1(G210), .A2(n682), .ZN(n608) );
  XOR2_X1 U680 ( .A(KEYINPUT116), .B(KEYINPUT54), .Z(n607) );
  BUF_X1 U681 ( .A(n604), .Z(n605) );
  XNOR2_X1 U682 ( .A(n605), .B(KEYINPUT55), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U684 ( .A(n611), .B(KEYINPUT62), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G472), .A2(n682), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X2 U687 ( .A1(n614), .A2(n698), .ZN(n616) );
  XNOR2_X1 U688 ( .A(KEYINPUT63), .B(KEYINPUT81), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n616), .B(n615), .ZN(G57) );
  XOR2_X1 U690 ( .A(G101), .B(n617), .Z(G3) );
  NOR2_X1 U691 ( .A1(n619), .A2(n630), .ZN(n618) );
  XOR2_X1 U692 ( .A(G104), .B(n618), .Z(G6) );
  NOR2_X1 U693 ( .A1(n619), .A2(n633), .ZN(n624) );
  XOR2_X1 U694 ( .A(KEYINPUT27), .B(KEYINPUT106), .Z(n621) );
  XNOR2_X1 U695 ( .A(G107), .B(KEYINPUT26), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U697 ( .A(KEYINPUT105), .B(n622), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n624), .B(n623), .ZN(G9) );
  XOR2_X1 U699 ( .A(n352), .B(G110), .Z(G12) );
  XNOR2_X1 U700 ( .A(KEYINPUT107), .B(KEYINPUT29), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U702 ( .A(G128), .B(n627), .ZN(G30) );
  XNOR2_X1 U703 ( .A(G143), .B(n628), .ZN(G45) );
  XOR2_X1 U704 ( .A(n629), .B(G146), .Z(G48) );
  NOR2_X1 U705 ( .A1(n630), .A2(n632), .ZN(n631) );
  XOR2_X1 U706 ( .A(G113), .B(n631), .Z(G15) );
  NOR2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U708 ( .A(KEYINPUT108), .B(n634), .Z(n635) );
  XNOR2_X1 U709 ( .A(G116), .B(n635), .ZN(G18) );
  XNOR2_X1 U710 ( .A(KEYINPUT37), .B(KEYINPUT109), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U712 ( .A(G125), .B(n638), .ZN(G27) );
  NOR2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U714 ( .A(KEYINPUT110), .B(n643), .Z(n648) );
  NOR2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U716 ( .A(KEYINPUT50), .B(n646), .ZN(n647) );
  NOR2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n649), .B(KEYINPUT111), .ZN(n651) );
  NOR2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U720 ( .A(KEYINPUT113), .B(n654), .Z(n655) );
  NOR2_X1 U721 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U722 ( .A(n657), .B(KEYINPUT114), .ZN(n661) );
  NOR2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U725 ( .A1(n668), .A2(n662), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n664), .A2(n663), .ZN(n665) );
  INV_X1 U727 ( .A(KEYINPUT2), .ZN(n669) );
  NOR2_X1 U728 ( .A1(KEYINPUT71), .A2(n669), .ZN(n671) );
  NAND2_X1 U729 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U730 ( .A(n674), .B(KEYINPUT115), .ZN(n675) );
  NOR2_X1 U731 ( .A1(G953), .A2(n675), .ZN(n676) );
  XNOR2_X1 U732 ( .A(KEYINPUT53), .B(n676), .ZN(G75) );
  NAND2_X1 U733 ( .A1(G469), .A2(n694), .ZN(n680) );
  XOR2_X1 U734 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n677) );
  XNOR2_X1 U735 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U736 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U737 ( .A1(n698), .A2(n681), .ZN(G54) );
  INV_X1 U738 ( .A(n698), .ZN(n688) );
  NAND2_X1 U739 ( .A1(G475), .A2(n682), .ZN(n686) );
  XOR2_X1 U740 ( .A(KEYINPUT59), .B(KEYINPUT117), .Z(n683) );
  XNOR2_X1 U741 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U742 ( .A(n689), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U743 ( .A1(G478), .A2(n694), .ZN(n690) );
  XNOR2_X1 U744 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U745 ( .A1(n698), .A2(n692), .ZN(G63) );
  XNOR2_X1 U746 ( .A(n693), .B(KEYINPUT118), .ZN(n696) );
  NAND2_X1 U747 ( .A1(n694), .A2(G217), .ZN(n695) );
  XNOR2_X1 U748 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U749 ( .A1(n698), .A2(n697), .ZN(G66) );
  XOR2_X1 U750 ( .A(KEYINPUT119), .B(KEYINPUT61), .Z(n700) );
  NAND2_X1 U751 ( .A1(G224), .A2(G953), .ZN(n699) );
  XNOR2_X1 U752 ( .A(n700), .B(n699), .ZN(n701) );
  NAND2_X1 U753 ( .A1(n701), .A2(G898), .ZN(n704) );
  NAND2_X1 U754 ( .A1(n702), .A2(n721), .ZN(n703) );
  NAND2_X1 U755 ( .A1(n704), .A2(n703), .ZN(n711) );
  XNOR2_X1 U756 ( .A(KEYINPUT120), .B(n706), .ZN(n708) );
  NOR2_X1 U757 ( .A1(n721), .A2(G898), .ZN(n707) );
  NOR2_X1 U758 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U759 ( .A(KEYINPUT121), .B(n709), .Z(n710) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(G69) );
  XOR2_X1 U761 ( .A(n713), .B(n712), .Z(n716) );
  XNOR2_X1 U762 ( .A(n716), .B(n714), .ZN(n715) );
  NOR2_X1 U763 ( .A1(G953), .A2(n715), .ZN(n724) );
  XNOR2_X1 U764 ( .A(n716), .B(G227), .ZN(n717) );
  XNOR2_X1 U765 ( .A(n717), .B(KEYINPUT122), .ZN(n718) );
  NAND2_X1 U766 ( .A1(n718), .A2(G900), .ZN(n719) );
  XNOR2_X1 U767 ( .A(KEYINPUT123), .B(n719), .ZN(n720) );
  NOR2_X1 U768 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U769 ( .A(n722), .B(KEYINPUT124), .ZN(n723) );
  NOR2_X1 U770 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U771 ( .A(KEYINPUT125), .B(n725), .ZN(G72) );
  XOR2_X1 U772 ( .A(G137), .B(KEYINPUT126), .Z(n726) );
  XNOR2_X1 U773 ( .A(n727), .B(n726), .ZN(G39) );
  XOR2_X1 U774 ( .A(n728), .B(G122), .Z(G24) );
  XOR2_X1 U775 ( .A(G140), .B(n729), .Z(G42) );
  XNOR2_X1 U776 ( .A(G119), .B(n730), .ZN(G21) );
  XOR2_X1 U777 ( .A(G131), .B(n731), .Z(G33) );
  XNOR2_X1 U778 ( .A(G134), .B(n732), .ZN(G36) );
endmodule

