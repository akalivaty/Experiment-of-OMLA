//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n449, new_n451, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n637, new_n638, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(new_n462));
  INV_X1    g037(.A(new_n456), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2106), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT70), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT70), .B1(new_n469), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(KEYINPUT71), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT3), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n480), .A2(G137), .A3(new_n467), .A4(new_n469), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n479), .ZN(new_n483));
  AND4_X1   g058(.A1(new_n482), .A2(new_n483), .A3(G101), .A4(new_n467), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n477), .B2(new_n479), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n485), .B2(G101), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n481), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n476), .A2(new_n487), .ZN(G160));
  NAND2_X1  g063(.A1(new_n480), .A2(new_n469), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(new_n467), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT73), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n489), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G136), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n468), .A2(G2104), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT70), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n504), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(G2105), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n480), .A2(new_n469), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n503), .A2(new_n505), .B1(new_n507), .B2(KEYINPUT4), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT74), .A2(G114), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT74), .A2(G114), .ZN(new_n510));
  OAI211_X1 g085(.A(KEYINPUT75), .B(G2105), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT74), .A2(G114), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT74), .A2(G114), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n467), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT75), .B1(G102), .B2(G2105), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n511), .B(G2104), .C1(new_n514), .C2(new_n516), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n480), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n508), .A2(new_n519), .ZN(G164));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(KEYINPUT76), .A2(KEYINPUT5), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G62), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n521), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT77), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT77), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT6), .B(G651), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n532), .A2(G543), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n533), .A2(G88), .B1(new_n534), .B2(G50), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  AND2_X1   g112(.A1(new_n533), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n532), .A2(G543), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n539), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n538), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n521), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n526), .A2(new_n532), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n548), .A2(new_n549), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n547), .A2(new_n551), .ZN(G171));
  AOI22_X1  g127(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n521), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT78), .B(G81), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n526), .A2(new_n532), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n532), .A2(G43), .A3(G543), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n557), .B1(new_n556), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n554), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT80), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n554), .B(new_n564), .C1(new_n560), .C2(new_n561), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n543), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n532), .A2(new_n574), .A3(G53), .A4(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(new_n525), .ZN(new_n578));
  AOI21_X1  g153(.A(G543), .B1(KEYINPUT76), .B2(KEYINPUT5), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n533), .A2(G91), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n576), .A2(new_n583), .A3(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  INV_X1    g161(.A(G168), .ZN(G286));
  NAND2_X1  g162(.A1(new_n533), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n534), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT81), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n524), .B2(new_n525), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT82), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n598), .B(G651), .C1(new_n593), .C2(new_n595), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G86), .ZN(new_n601));
  INV_X1    g176(.A(G48), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n548), .A2(new_n601), .B1(new_n543), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G305));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  INV_X1    g181(.A(G72), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n580), .A2(new_n606), .B1(new_n607), .B2(new_n523), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT83), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n610), .B1(new_n607), .B2(new_n523), .C1(new_n580), .C2(new_n606), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n609), .A2(G651), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT85), .B(G47), .Z(new_n616));
  AOI22_X1  g191(.A1(new_n533), .A2(G85), .B1(new_n534), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(G290));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n580), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G651), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT86), .B(KEYINPUT10), .Z(new_n623));
  NAND3_X1  g198(.A1(new_n533), .A2(G92), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n534), .A2(G54), .ZN(new_n625));
  INV_X1    g200(.A(new_n623), .ZN(new_n626));
  INV_X1    g201(.A(G92), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n548), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n622), .A2(new_n624), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(G171), .ZN(G284));
  OAI21_X1  g207(.A(new_n631), .B1(new_n630), .B2(G171), .ZN(G321));
  NAND2_X1  g208(.A1(G299), .A2(new_n630), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n630), .B2(G168), .ZN(G297));
  OAI21_X1  g210(.A(new_n634), .B1(new_n630), .B2(G168), .ZN(G280));
  INV_X1    g211(.A(new_n629), .ZN(new_n637));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n566), .B2(G868), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n503), .A2(new_n485), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT13), .Z(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT87), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n495), .A2(G135), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n490), .A2(G123), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n467), .A2(G111), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n646), .B2(new_n647), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n656), .ZN(G156));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  NOR2_X1   g250(.A1(G2072), .A2(G2078), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n442), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n673), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(KEYINPUT17), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n675), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n673), .B(new_n674), .C1(new_n442), .C2(new_n676), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT18), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n675), .A3(new_n673), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT89), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1961), .B(G1966), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT90), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n688), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n694), .B2(new_n693), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(new_n688), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n690), .A2(new_n692), .ZN(new_n701));
  MUX2_X1   g276(.A(new_n700), .B(new_n688), .S(new_n701), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT92), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n705), .B(new_n709), .ZN(G229));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n566), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(G19), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G1341), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(G1341), .ZN(new_n716));
  INV_X1    g291(.A(G2090), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n718), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT29), .Z(new_n721));
  OAI211_X1 g296(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n717), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT100), .B(KEYINPUT28), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n718), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n495), .A2(G140), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n490), .A2(G128), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT98), .B1(G104), .B2(G2105), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g305(.A1(KEYINPUT98), .A2(G104), .A3(G2105), .ZN(new_n731));
  OAI221_X1 g306(.A(G2104), .B1(G116), .B2(new_n467), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n727), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT99), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n727), .A2(new_n728), .A3(KEYINPUT99), .A4(new_n732), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n726), .B1(new_n737), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2067), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n723), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G11), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(G28), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n718), .B1(new_n742), .B2(G28), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n741), .B1(new_n743), .B2(new_n744), .C1(new_n654), .C2(new_n718), .ZN(new_n745));
  NOR2_X1   g320(.A1(G171), .A2(new_n711), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G5), .B2(new_n711), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n745), .B1(new_n748), .B2(G1961), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n637), .A2(new_n711), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G4), .B2(new_n711), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n718), .A2(G32), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n495), .A2(G141), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n490), .A2(G129), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI22_X1  g335(.A1(G105), .A2(new_n485), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n755), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n754), .B1(new_n763), .B2(new_n718), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n764), .B(new_n765), .Z(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n711), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n711), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n747), .A2(new_n767), .B1(G1966), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G1966), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n711), .A2(G20), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT23), .Z(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G299), .B2(G16), .ZN(new_n774));
  INV_X1    g349(.A(G1956), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR4_X1   g351(.A1(new_n753), .A2(new_n766), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n752), .A2(new_n750), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n718), .A2(G33), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n467), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n495), .A2(G139), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT25), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(new_n718), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G2072), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n718), .B1(new_n789), .B2(G34), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n789), .B2(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G160), .B2(G29), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G2084), .ZN(new_n793));
  NAND2_X1  g368(.A1(G164), .A2(G29), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G27), .B2(G29), .ZN(new_n795));
  INV_X1    g370(.A(G2078), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n778), .A2(new_n788), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n787), .A2(G2072), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n799), .B1(new_n796), .B2(new_n795), .C1(G2084), .C2(new_n792), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n777), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n722), .A2(new_n740), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G290), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G16), .B2(G24), .ZN(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G25), .A2(G29), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n495), .A2(G131), .ZN(new_n811));
  OR2_X1    g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n490), .A2(G119), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT93), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT93), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n810), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT94), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n807), .B2(new_n808), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n711), .A2(G23), .ZN(new_n824));
  INV_X1    g399(.A(G288), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(new_n711), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT33), .ZN(new_n827));
  INV_X1    g402(.A(G1976), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n711), .A2(G22), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT96), .Z(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G166), .B2(new_n711), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT97), .B(G1971), .Z(new_n833));
  XOR2_X1   g408(.A(new_n832), .B(new_n833), .Z(new_n834));
  NOR2_X1   g409(.A1(G6), .A2(G16), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n604), .B2(G16), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT32), .B(G1981), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT95), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n836), .B(new_n838), .Z(new_n839));
  NOR3_X1   g414(.A1(new_n829), .A2(new_n834), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT34), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n809), .B(new_n823), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n804), .B1(new_n845), .B2(new_n846), .ZN(G311));
  INV_X1    g422(.A(new_n846), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n803), .B1(new_n848), .B2(new_n849), .ZN(G150));
  NOR2_X1   g425(.A1(new_n629), .A2(new_n638), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n533), .A2(G93), .B1(new_n534), .B2(G55), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n521), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n563), .A2(new_n565), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(KEYINPUT101), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n853), .B(new_n858), .C1(new_n521), .C2(new_n854), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n562), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n852), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n863));
  AOI21_X1  g438(.A(G860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n857), .A2(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(G145));
  XNOR2_X1  g444(.A(new_n786), .B(KEYINPUT102), .ZN(new_n870));
  AOI21_X1  g445(.A(G164), .B1(new_n735), .B2(new_n736), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n735), .A2(G164), .A3(new_n736), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n762), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n875), .A2(new_n763), .A3(new_n871), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n870), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n816), .A2(new_n817), .ZN(new_n878));
  INV_X1    g453(.A(new_n814), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n645), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n495), .A2(G142), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n490), .A2(G130), .ZN(new_n883));
  OR2_X1    g458(.A1(G106), .A2(G2105), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n884), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n645), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n818), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n881), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n887), .B1(new_n881), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n763), .B1(new_n875), .B2(new_n871), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n872), .A2(new_n762), .A3(new_n873), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n786), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n877), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n877), .A2(new_n896), .ZN(new_n900));
  INV_X1    g475(.A(new_n892), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n892), .A2(new_n877), .A3(new_n896), .A4(KEYINPUT103), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n654), .B(G160), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(G162), .Z(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G37), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n897), .A2(new_n906), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n892), .B1(new_n896), .B2(new_n877), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT104), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n902), .A2(new_n912), .A3(new_n906), .A4(new_n897), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g491(.A(new_n861), .B(new_n640), .Z(new_n917));
  XNOR2_X1  g492(.A(new_n629), .B(G299), .ZN(new_n918));
  XNOR2_X1  g493(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT106), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(KEYINPUT41), .B2(new_n918), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n923), .B2(KEYINPUT106), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n918), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n917), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT42), .ZN(new_n930));
  XNOR2_X1  g505(.A(G290), .B(G288), .ZN(new_n931));
  XNOR2_X1  g506(.A(G303), .B(new_n604), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n805), .A2(G288), .ZN(new_n935));
  NOR2_X1   g510(.A1(G290), .A2(new_n825), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(KEYINPUT107), .B2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n925), .B(new_n927), .C1(KEYINPUT107), .C2(new_n940), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n930), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n930), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(G868), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n866), .A2(new_n630), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(G295));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n946), .ZN(G331));
  XNOR2_X1  g523(.A(G168), .B(G171), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n856), .A2(new_n949), .A3(new_n860), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n856), .B2(new_n860), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n924), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n926), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n956), .B2(new_n938), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n629), .A2(G299), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n629), .A2(G299), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n959), .B(KEYINPUT41), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n962), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n960), .A3(new_n919), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n959), .B1(new_n918), .B2(KEYINPUT41), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT109), .B1(new_n968), .B2(new_n952), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  OAI221_X1 g545(.A(new_n970), .B1(new_n950), .B2(new_n951), .C1(new_n967), .C2(new_n966), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n971), .A3(new_n954), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n972), .A2(new_n973), .A3(new_n939), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n972), .B2(new_n939), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n957), .B(new_n958), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n939), .B1(new_n953), .B2(new_n955), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n938), .B(new_n954), .C1(new_n924), .C2(new_n952), .ZN(new_n979));
  INV_X1    g554(.A(G37), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n976), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n977), .A2(new_n958), .A3(new_n980), .A4(new_n979), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n986), .B2(KEYINPUT111), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n957), .A2(new_n988), .A3(new_n958), .A4(new_n977), .ZN(new_n989));
  INV_X1    g564(.A(new_n975), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n972), .A2(new_n973), .A3(new_n939), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n987), .B(new_n989), .C1(new_n992), .C2(new_n958), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n985), .A2(new_n993), .ZN(G397));
  INV_X1    g569(.A(KEYINPUT62), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n508), .B2(new_n519), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G40), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n476), .A2(new_n487), .A3(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(KEYINPUT45), .B(new_n996), .C1(new_n508), .C2(new_n519), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1966), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(G2084), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(new_n996), .C1(new_n508), .C2(new_n519), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1006), .A2(new_n1007), .A3(new_n1001), .A4(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(G168), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  AOI21_X1  g587(.A(G168), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1011), .A2(new_n1016), .A3(G8), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1015), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n995), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT121), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(KEYINPUT62), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT114), .B(G1971), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1003), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1006), .A2(new_n717), .A3(new_n1001), .A4(new_n1009), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND3_X1   g604(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n517), .A2(new_n518), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n505), .B1(new_n472), .B2(new_n473), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(G160), .A3(G40), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT115), .B1(new_n1040), .B2(G8), .ZN(new_n1041));
  INV_X1    g616(.A(G125), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n501), .B2(new_n502), .ZN(new_n1043));
  INV_X1    g618(.A(new_n475), .ZN(new_n1044));
  OAI21_X1  g619(.A(G2105), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n483), .A2(G101), .A3(new_n467), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT72), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n485), .A2(new_n482), .A3(G101), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1045), .A2(G40), .A3(new_n481), .A4(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT115), .B(G8), .C1(new_n1050), .C2(new_n997), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1041), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G288), .A2(new_n828), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1054), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n828), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1056), .B(new_n1057), .C1(new_n1041), .C2(new_n1052), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n597), .A2(KEYINPUT116), .A3(new_n599), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G1981), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT49), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT49), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1062), .A3(G1981), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(new_n604), .A3(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1059), .A2(new_n1062), .A3(G1981), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1062), .B1(new_n1059), .B2(G1981), .ZN(new_n1066));
  OAI21_X1  g641(.A(G305), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1064), .B(new_n1067), .C1(new_n1041), .C2(new_n1052), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1034), .A2(new_n1055), .A3(new_n1058), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1006), .A2(new_n1001), .A3(new_n1009), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1072), .A2(new_n717), .B1(new_n1003), .B2(new_n1026), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT117), .B(new_n1032), .C1(new_n1073), .C2(new_n1025), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1003), .B2(G2078), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1006), .A2(new_n1001), .A3(new_n1009), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n767), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1003), .A2(new_n1076), .A3(G2078), .ZN(new_n1081));
  OAI21_X1  g656(.A(G171), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1069), .A2(new_n1075), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1020), .A2(new_n1024), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1050), .A2(new_n997), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(new_n1025), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1054), .B1(new_n1088), .B2(new_n1051), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1058), .B(new_n1068), .C1(new_n1085), .C2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G305), .A2(G1981), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G288), .A2(G1976), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1068), .B2(new_n1092), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1090), .A2(new_n1034), .B1(new_n1093), .B2(new_n1053), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1073), .A2(new_n1025), .A3(new_n1032), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1072), .A2(new_n1007), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G168), .A2(G8), .ZN(new_n1099));
  OR3_X1    g674(.A1(new_n1098), .A2(KEYINPUT118), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT118), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1095), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1032), .B1(new_n1073), .B2(new_n1025), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1097), .A2(new_n1102), .A3(KEYINPUT63), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1094), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n576), .B2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(G299), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1078), .A2(new_n775), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1078), .A2(new_n750), .ZN(new_n1117));
  INV_X1    g692(.A(G2067), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1087), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n629), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1113), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1113), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(new_n1116), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1112), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(KEYINPUT61), .A3(new_n1123), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT58), .B(G1341), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1003), .A2(G1996), .B1(new_n1087), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n566), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1135));
  AND2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1127), .B(new_n1131), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n629), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n637), .B1(new_n1120), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1139), .A2(new_n1141), .B1(new_n1140), .B2(new_n1120), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1124), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1050), .B(KEYINPUT123), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT53), .B1(new_n1145), .B2(G2078), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1145), .B2(G2078), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1144), .A2(new_n999), .A3(new_n1002), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(new_n1079), .A3(new_n1077), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G171), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT125), .ZN(new_n1151));
  OR3_X1    g726(.A1(new_n1080), .A2(G171), .A3(new_n1081), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1149), .A2(new_n1153), .A3(G171), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1151), .A2(KEYINPUT54), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1148), .A2(G301), .A3(new_n1079), .A4(new_n1077), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1082), .B2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1158), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1109), .A2(new_n1143), .A3(new_n1155), .A4(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1084), .A2(new_n1108), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n999), .A2(new_n1050), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n737), .A2(G2067), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n735), .A2(new_n1118), .A3(new_n736), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n762), .A2(G1996), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n999), .A2(G1996), .A3(new_n1050), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT112), .B1(new_n1168), .B2(new_n763), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1168), .A2(KEYINPUT112), .A3(new_n763), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1167), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT113), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1171), .A2(KEYINPUT113), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n818), .A2(new_n820), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n818), .A2(new_n820), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1162), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n805), .A2(new_n808), .ZN(new_n1177));
  NOR2_X1   g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1162), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AND4_X1   g754(.A1(new_n1172), .A2(new_n1173), .A3(new_n1176), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1161), .A2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1168), .B(KEYINPUT46), .Z(new_n1182));
  OAI21_X1  g757(.A(new_n1162), .B1(new_n1165), .B2(new_n762), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT47), .Z(new_n1185));
  NAND2_X1  g760(.A1(new_n1178), .A2(new_n1162), .ZN(new_n1186));
  XOR2_X1   g761(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1187));
  XNOR2_X1  g762(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  AND4_X1   g763(.A1(new_n1172), .A2(new_n1173), .A3(new_n1176), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1173), .A2(new_n1172), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1174), .B(KEYINPUT126), .Z(new_n1191));
  OAI21_X1  g766(.A(new_n1164), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g767(.A(new_n1185), .B(new_n1189), .C1(new_n1162), .C2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1181), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g769(.A1(G229), .A2(new_n465), .A3(G401), .A4(G227), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n983), .A2(new_n915), .A3(new_n1196), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


