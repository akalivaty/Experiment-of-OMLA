//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G77), .A2(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G97), .C2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT64), .Z(new_n225));
  NOR2_X1   g0025(.A1(new_n222), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n220), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI22_X1  g0032(.A1(new_n223), .A2(KEYINPUT1), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n225), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n217), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n213), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G97), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G87), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n212), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G223), .A3(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G222), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n252), .B1(new_n253), .B2(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  OAI211_X1 g0059(.A(G1), .B(G13), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n260), .A2(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G226), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n262), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G190), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(G200), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT9), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n219), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n202), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n229), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(KEYINPUT67), .A3(new_n277), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n219), .A2(G20), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n283), .B(new_n284), .C1(KEYINPUT67), .C2(new_n282), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n220), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(G20), .B2(new_n203), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n279), .B1(new_n285), .B2(new_n202), .C1(new_n282), .C2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n274), .A2(new_n275), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n273), .A2(new_n276), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n273), .A2(new_n295), .A3(new_n298), .A4(new_n276), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT14), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n251), .A2(G232), .A3(G1698), .ZN(new_n303));
  INV_X1    g0103(.A(G97), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n303), .B1(new_n258), .B2(new_n304), .C1(new_n255), .C2(new_n211), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n265), .B1(new_n305), .B2(new_n261), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n267), .A2(G238), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n310));
  OAI211_X1 g0110(.A(G169), .B(new_n302), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n306), .A2(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT13), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(G179), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n313), .B2(new_n314), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT70), .B(KEYINPUT14), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n311), .B(new_n315), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n207), .A2(G20), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n320), .B1(new_n287), .B2(new_n253), .C1(new_n290), .C2(new_n202), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n281), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT11), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n278), .A2(new_n207), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT12), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(KEYINPUT11), .A3(new_n281), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n281), .B1(new_n219), .B2(G20), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G68), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n324), .A2(new_n326), .A3(new_n327), .A4(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n313), .A2(new_n314), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(G200), .B1(new_n331), .B2(new_n332), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n313), .A2(G190), .A3(new_n314), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n319), .A2(new_n333), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n270), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(new_n293), .C1(G169), .C2(new_n270), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n267), .A2(G244), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n251), .A2(G232), .A3(new_n254), .ZN(new_n343));
  INV_X1    g0143(.A(G107), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(new_n251), .ZN(new_n345));
  AOI211_X1 g0145(.A(new_n265), .B(new_n341), .C1(new_n345), .C2(new_n261), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n338), .ZN(new_n347));
  INV_X1    g0147(.A(new_n286), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT15), .B(G87), .Z(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n287), .B2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n281), .B1(new_n253), .B2(new_n278), .ZN(new_n353));
  INV_X1    g0153(.A(new_n328), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n253), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n347), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n346), .A2(G169), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n300), .A2(new_n337), .A3(new_n340), .A4(new_n359), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n220), .B(G87), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT22), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(KEYINPUT82), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT84), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n220), .B2(G107), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT23), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT23), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n368), .B(new_n371), .C1(new_n220), .C2(G107), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n220), .A2(G33), .A3(G116), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT83), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n367), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n365), .B(G87), .C1(new_n362), .C2(new_n361), .ZN(new_n378));
  NAND3_X1  g0178(.A1(KEYINPUT83), .A2(G33), .A3(G116), .ZN(new_n379));
  AOI21_X1  g0179(.A(G20), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT85), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n220), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT85), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n370), .A2(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n367), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n386), .A3(KEYINPUT24), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT24), .ZN(new_n388));
  OAI211_X1 g0188(.A(KEYINPUT85), .B(new_n388), .C1(new_n377), .C2(new_n380), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n281), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n219), .A2(G33), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n282), .A2(new_n277), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT25), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n277), .B2(G107), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n278), .A2(KEYINPUT25), .A3(new_n344), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n393), .A2(G107), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n251), .A2(G257), .A3(G1698), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n251), .A2(G250), .A3(new_n254), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G294), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G45), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(G1), .ZN(new_n404));
  AND2_X1   g0204(.A1(KEYINPUT5), .A2(G41), .ZN(new_n405));
  NOR2_X1   g0205(.A1(KEYINPUT5), .A2(G41), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n260), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n402), .A2(new_n261), .B1(new_n409), .B2(G264), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT5), .B(G41), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(G274), .A3(new_n404), .ZN(new_n412));
  AOI21_X1  g0212(.A(G169), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n402), .A2(new_n261), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n409), .A2(G264), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(G179), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n398), .A2(new_n414), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT21), .ZN(new_n421));
  OAI211_X1 g0221(.A(G264), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT80), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n251), .A2(KEYINPUT80), .A3(G264), .A4(G1698), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n251), .A2(G257), .A3(new_n254), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n361), .A2(new_n362), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G303), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n429), .A2(KEYINPUT81), .A3(new_n261), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n407), .A2(G270), .A3(new_n260), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n431), .A2(KEYINPUT79), .A3(new_n412), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT79), .B1(new_n431), .B2(new_n412), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT81), .B1(new_n429), .B2(new_n261), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n430), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G283), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n220), .C1(G33), .C2(new_n304), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n212), .A2(G20), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n281), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT20), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n441), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n442), .A2(new_n443), .B1(new_n212), .B2(new_n278), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n393), .A2(G116), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G169), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n421), .B1(new_n436), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n430), .A2(new_n435), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n431), .A2(new_n412), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n431), .A2(KEYINPUT79), .A3(new_n412), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n449), .A2(G179), .A3(new_n446), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n429), .A2(new_n261), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT81), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n429), .A2(KEYINPUT81), .A3(new_n261), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n316), .B1(new_n444), .B2(new_n445), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(KEYINPUT21), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n420), .A2(new_n448), .A3(new_n455), .A4(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n277), .A2(G97), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n392), .B2(new_n304), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT74), .B1(new_n289), .B2(G77), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n344), .A2(KEYINPUT6), .A3(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n344), .A2(G97), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n304), .A2(G107), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(KEYINPUT6), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n467), .B1(new_n472), .B2(G20), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT7), .B1(new_n427), .B2(new_n220), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT7), .ZN(new_n475));
  NOR4_X1   g0275(.A1(new_n361), .A2(new_n362), .A3(new_n475), .A4(G20), .ZN(new_n476));
  OAI21_X1  g0276(.A(G107), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n289), .A2(KEYINPUT74), .A3(G77), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n466), .B1(new_n479), .B2(new_n281), .ZN(new_n480));
  OAI211_X1 g0280(.A(G244), .B(new_n254), .C1(new_n361), .C2(new_n362), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(KEYINPUT76), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(KEYINPUT76), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n251), .A2(G244), .A3(new_n254), .A4(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n483), .A2(new_n437), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n261), .ZN(new_n488));
  INV_X1    g0288(.A(G257), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n412), .B1(new_n408), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G169), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n487), .B2(new_n261), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G179), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n480), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT75), .ZN(new_n497));
  INV_X1    g0297(.A(new_n467), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n344), .A2(KEYINPUT6), .A3(G97), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n247), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n498), .B1(new_n501), .B2(new_n220), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT3), .A2(G33), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT3), .A2(G33), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n220), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n475), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n503), .A2(KEYINPUT7), .A3(new_n220), .A4(new_n504), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n344), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n282), .B1(new_n509), .B2(new_n478), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n497), .B1(new_n510), .B2(new_n466), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n480), .A2(KEYINPUT75), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G190), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n494), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G200), .B2(new_n494), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n496), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n350), .A2(new_n277), .ZN(new_n518));
  INV_X1    g0318(.A(G87), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n392), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n251), .A2(new_n220), .A3(G68), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT19), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n287), .B2(new_n304), .ZN(new_n523));
  XOR2_X1   g0323(.A(KEYINPUT78), .B(G87), .Z(new_n524));
  NOR3_X1   g0324(.A1(new_n524), .A2(G97), .A3(G107), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n258), .A2(new_n304), .ZN(new_n526));
  AOI21_X1  g0326(.A(G20), .B1(new_n526), .B2(KEYINPUT19), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n521), .B(new_n523), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  AOI211_X1 g0328(.A(new_n518), .B(new_n520), .C1(new_n528), .C2(new_n281), .ZN(new_n529));
  OAI211_X1 g0329(.A(G238), .B(new_n254), .C1(new_n361), .C2(new_n362), .ZN(new_n530));
  OAI211_X1 g0330(.A(G244), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT77), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT77), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n530), .A2(new_n531), .A3(new_n535), .A4(new_n532), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n261), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n404), .A2(G274), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n260), .B(G250), .C1(G1), .C2(new_n403), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n537), .A2(G190), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n541));
  INV_X1    g0341(.A(G200), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n529), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n316), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n518), .B1(new_n528), .B2(new_n281), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n393), .A2(new_n350), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n537), .A2(new_n338), .A3(new_n538), .A4(new_n539), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n417), .A2(new_n542), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n410), .A2(new_n514), .A3(new_n412), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n390), .A2(new_n554), .A3(new_n397), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n460), .A2(G200), .ZN(new_n556));
  INV_X1    g0356(.A(new_n446), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n556), .B(new_n557), .C1(new_n514), .C2(new_n460), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n517), .A2(new_n551), .A3(new_n555), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n506), .A2(KEYINPUT71), .A3(new_n507), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n507), .A2(KEYINPUT71), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(G68), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n216), .A2(new_n207), .ZN(new_n563));
  OAI21_X1  g0363(.A(G20), .B1(new_n563), .B2(new_n201), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n289), .A2(G159), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(KEYINPUT16), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT16), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n207), .B1(new_n506), .B2(new_n507), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n566), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n281), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n285), .A2(new_n348), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n278), .B2(new_n348), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT17), .ZN(new_n577));
  OAI211_X1 g0377(.A(G223), .B(new_n254), .C1(new_n361), .C2(new_n362), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT72), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n251), .A2(KEYINPUT72), .A3(G223), .A4(new_n254), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G87), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n251), .A2(G226), .A3(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n261), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n260), .A2(G232), .A3(new_n263), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT73), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT73), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n260), .A2(new_n588), .A3(G232), .A4(new_n263), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(new_n266), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G200), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n585), .A2(G190), .A3(new_n590), .A4(new_n266), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n576), .A2(new_n577), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n572), .A2(new_n592), .A3(new_n574), .A4(new_n593), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT17), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n585), .A2(G179), .A3(new_n590), .A4(new_n266), .ZN(new_n597));
  AOI221_X4 g0397(.A(new_n265), .B1(new_n587), .B2(new_n589), .C1(new_n584), .C2(new_n261), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(new_n316), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n575), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT18), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n575), .A2(new_n599), .A3(KEYINPUT18), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n594), .A2(new_n596), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n346), .A2(new_n542), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n355), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n346), .A2(G190), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NOR4_X1   g0409(.A1(new_n360), .A2(new_n463), .A3(new_n559), .A4(new_n609), .ZN(G372));
  INV_X1    g0410(.A(new_n340), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n319), .A2(new_n333), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n335), .A2(new_n336), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n359), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n594), .A2(new_n596), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n614), .A2(new_n615), .B1(new_n602), .B2(new_n603), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n616), .A2(KEYINPUT88), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n616), .A2(KEYINPUT88), .B1(new_n297), .B2(new_n299), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n360), .A2(new_n609), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT86), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n420), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n455), .A2(new_n462), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT21), .B1(new_n460), .B2(new_n461), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n398), .A2(KEYINPUT86), .A3(new_n414), .A4(new_n419), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n622), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT87), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n479), .A2(new_n281), .ZN(new_n630));
  INV_X1    g0430(.A(new_n466), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT75), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI211_X1 g0432(.A(new_n497), .B(new_n466), .C1(new_n479), .C2(new_n281), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n516), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n493), .A2(new_n495), .ZN(new_n635));
  INV_X1    g0435(.A(new_n480), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n637), .A3(new_n555), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n543), .A2(new_n550), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n622), .A2(new_n625), .A3(KEYINPUT87), .A4(new_n626), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n629), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n635), .A2(new_n511), .A3(new_n512), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n551), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n550), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n543), .A2(new_n496), .A3(new_n550), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(KEYINPUT26), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n620), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n619), .A2(new_n650), .ZN(G369));
  NAND3_X1  g0451(.A1(new_n448), .A2(new_n455), .A3(new_n462), .ZN(new_n652));
  INV_X1    g0452(.A(G13), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G20), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n219), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n652), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n398), .A2(new_n660), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n420), .A2(new_n555), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n662), .B(new_n664), .C1(new_n420), .C2(new_n661), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n558), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n625), .B1(new_n557), .B2(new_n661), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n652), .A2(new_n446), .A3(new_n660), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(G330), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n622), .A2(new_n626), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n661), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n665), .A2(new_n674), .A3(KEYINPUT89), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT89), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n662), .A2(new_n664), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n660), .B1(new_n622), .B2(new_n626), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n672), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n226), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n525), .A2(new_n212), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n686), .A3(G1), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n231), .B2(new_n684), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT92), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n460), .A2(new_n338), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT90), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n541), .A2(new_n692), .A3(new_n410), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n415), .A2(new_n416), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT90), .B1(new_n544), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n691), .A2(new_n693), .A3(new_n494), .A4(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT91), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n544), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n537), .A2(KEYINPUT91), .A3(new_n538), .A4(new_n539), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n700), .A2(new_n492), .A3(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n460), .A2(new_n338), .A3(new_n417), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n690), .B1(new_n698), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n693), .A2(new_n695), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n691), .A4(new_n494), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n696), .A2(new_n697), .B1(new_n702), .B2(new_n703), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT92), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n661), .B1(new_n708), .B2(new_n707), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n559), .A2(new_n463), .A3(new_n660), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n647), .A2(new_n643), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT94), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n551), .A2(KEYINPUT26), .A3(new_n644), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n647), .A2(KEYINPUT94), .A3(new_n643), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n640), .A2(new_n463), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n550), .B(KEYINPUT93), .Z(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n661), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n660), .B1(new_n642), .B2(new_n648), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n718), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n689), .B1(new_n734), .B2(G1), .ZN(G364));
  AOI21_X1  g0535(.A(new_n219), .B1(new_n654), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n683), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(G1), .B(G13), .C1(new_n220), .C2(G169), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT95), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n220), .A2(G190), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n542), .A2(G179), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n344), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n220), .A2(new_n514), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n745), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n427), .B(new_n747), .C1(new_n524), .C2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT96), .Z(new_n752));
  NAND3_X1  g0552(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n338), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G50), .A2(new_n756), .B1(new_n759), .B2(G58), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n744), .A2(new_n757), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n760), .B1(new_n253), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n744), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G159), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT32), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n220), .B1(new_n764), .B2(G190), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n304), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n763), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT97), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n754), .B2(new_n514), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n753), .A2(KEYINPUT97), .A3(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n752), .B(new_n771), .C1(new_n207), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n427), .B1(new_n762), .B2(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G322), .A2(new_n759), .B1(new_n766), .B2(G329), .ZN(new_n779));
  INV_X1    g0579(.A(G303), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n780), .B2(new_n749), .ZN(new_n781));
  INV_X1    g0581(.A(new_n775), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n778), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n755), .B(KEYINPUT98), .ZN(new_n785));
  INV_X1    g0585(.A(new_n769), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n785), .A2(G326), .B1(G294), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT99), .ZN(new_n788));
  INV_X1    g0588(.A(G283), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n784), .B(new_n788), .C1(new_n789), .C2(new_n746), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n743), .B1(new_n776), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n742), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n246), .A2(G45), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n682), .A2(new_n251), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(G45), .C2(new_n231), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n226), .A2(G355), .A3(new_n251), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(G116), .C2(new_n226), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n791), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n794), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n738), .B(new_n801), .C1(new_n671), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n671), .A2(G330), .ZN(new_n804));
  INV_X1    g0604(.A(new_n738), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n671), .A2(G330), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(G396));
  INV_X1    g0608(.A(KEYINPUT101), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n358), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n358), .A2(new_n809), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n811), .A2(new_n812), .B1(new_n607), .B2(new_n606), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n649), .A2(new_n661), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n355), .A2(new_n660), .ZN(new_n815));
  INV_X1    g0615(.A(new_n812), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n608), .B(new_n815), .C1(new_n816), .C2(new_n810), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n359), .B2(new_n661), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n814), .B1(new_n730), .B2(new_n818), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(new_n718), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n718), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n820), .A2(new_n805), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G107), .A2(new_n750), .B1(new_n766), .B2(G311), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n212), .B2(new_n762), .C1(new_n824), .C2(new_n758), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n770), .B(new_n825), .C1(G303), .C2(new_n756), .ZN(new_n826));
  INV_X1    g0626(.A(new_n746), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G87), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n782), .A2(G283), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n826), .A2(new_n427), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n746), .A2(new_n207), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n756), .A2(G137), .B1(new_n761), .B2(G159), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n759), .A2(G143), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n288), .C2(new_n775), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT34), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n251), .B1(new_n765), .B2(new_n838), .C1(new_n202), .C2(new_n749), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G58), .B2(new_n786), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n836), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n830), .B1(new_n831), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n742), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n742), .A2(new_n792), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n738), .B1(new_n845), .B2(G77), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT100), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n843), .B(new_n847), .C1(new_n818), .C2(new_n793), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n822), .A2(new_n848), .ZN(G384));
  NAND2_X1  g0649(.A1(new_n333), .A2(new_n660), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n337), .A2(KEYINPUT103), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n337), .B2(KEYINPUT103), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n813), .A2(new_n815), .B1(new_n358), .B2(new_n660), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n715), .B(new_n661), .C1(new_n708), .C2(new_n707), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT107), .B1(new_n716), .B2(new_n857), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n413), .B(new_n418), .C1(new_n390), .C2(new_n397), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n652), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n640), .A2(new_n860), .A3(new_n558), .A4(new_n661), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n712), .B1(new_n861), .B2(KEYINPUT31), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT107), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n862), .A2(new_n863), .A3(new_n856), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n855), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT109), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n658), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n575), .B1(new_n599), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n870), .A3(new_n595), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT106), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT106), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n869), .A2(new_n873), .A3(new_n870), .A4(new_n595), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n568), .A2(new_n281), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT16), .B1(new_n562), .B2(new_n567), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n574), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT104), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT104), .B(new_n574), .C1(new_n876), .C2(new_n877), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n597), .B(new_n658), .C1(new_n598), .C2(new_n316), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n595), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n875), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n868), .A3(new_n881), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n602), .A2(new_n603), .ZN(new_n888));
  AOI211_X1 g0688(.A(KEYINPUT105), .B(new_n887), .C1(new_n615), .C2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n595), .A2(KEYINPUT17), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n595), .A2(KEYINPUT17), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n575), .A2(new_n599), .A3(KEYINPUT18), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT18), .B1(new_n575), .B2(new_n599), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n891), .A2(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n887), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(KEYINPUT38), .B(new_n886), .C1(new_n889), .C2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n604), .A2(new_n576), .A3(new_n658), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n870), .B1(new_n869), .B2(new_n595), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n872), .B2(new_n874), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n716), .A2(KEYINPUT107), .A3(new_n857), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n863), .B1(new_n862), .B2(new_n856), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(KEYINPUT109), .A3(new_n855), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n867), .A2(KEYINPUT40), .A3(new_n904), .A4(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT108), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n818), .B1(new_n851), .B2(new_n852), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n905), .B2(new_n906), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n886), .B1(new_n889), .B2(new_n897), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n899), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n898), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI211_X1 g0718(.A(KEYINPUT108), .B(KEYINPUT40), .C1(new_n912), .C2(new_n915), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n909), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n907), .A2(new_n620), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n920), .B(new_n921), .Z(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(G330), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n888), .A2(new_n868), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n816), .A2(new_n660), .A3(new_n810), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n853), .B1(new_n814), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n924), .B1(new_n927), .B2(new_n915), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n612), .A2(new_n660), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n914), .B2(new_n898), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n898), .A2(new_n903), .A3(new_n930), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n929), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n732), .A2(new_n729), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n620), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n619), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n935), .B(new_n938), .Z(new_n939));
  XNOR2_X1  g0739(.A(new_n923), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n219), .B2(new_n654), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n212), .B1(new_n472), .B2(KEYINPUT35), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n942), .B(new_n230), .C1(KEYINPUT35), .C2(new_n472), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT36), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n563), .A2(new_n231), .A3(new_n253), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT102), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n207), .A2(G50), .ZN(new_n947));
  OAI211_X1 g0747(.A(G1), .B(new_n653), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n941), .A2(new_n944), .A3(new_n948), .ZN(G367));
  NOR2_X1   g0749(.A1(new_n749), .A2(new_n212), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n950), .A2(KEYINPUT46), .B1(new_n344), .B2(new_n769), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n251), .B(new_n951), .C1(KEYINPUT46), .C2(new_n950), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n759), .A2(G303), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G311), .A2(new_n785), .B1(new_n782), .B2(G294), .ZN(new_n954));
  INV_X1    g0754(.A(G317), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n762), .A2(new_n789), .B1(new_n765), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n746), .A2(new_n304), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n746), .A2(new_n253), .ZN(new_n960));
  AOI22_X1  g0760(.A1(G150), .A2(new_n759), .B1(new_n750), .B2(G58), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n202), .B2(new_n762), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n960), .B(new_n962), .C1(G137), .C2(new_n766), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n785), .A2(G143), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n207), .C2(new_n769), .ZN(new_n965));
  INV_X1    g0765(.A(G159), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n251), .B1(new_n775), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n959), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n805), .B1(new_n969), .B2(new_n742), .ZN(new_n970));
  INV_X1    g0770(.A(new_n797), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n795), .B1(new_n226), .B2(new_n351), .C1(new_n242), .C2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n529), .A2(new_n661), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n551), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n550), .B2(new_n973), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(new_n802), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n970), .A2(new_n972), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n517), .B1(new_n513), .B2(new_n661), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n644), .A2(new_n660), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n672), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n982), .A2(new_n665), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n637), .B1(new_n982), .B2(new_n420), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n661), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT110), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n991), .A3(new_n988), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n975), .B(KEYINPUT43), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n990), .A2(new_n992), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n984), .B(new_n994), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  AND3_X1   g0797(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n996), .B1(new_n990), .B2(new_n992), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n983), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n680), .A2(new_n981), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n680), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n680), .B2(new_n981), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n675), .A2(new_n679), .A3(KEYINPUT44), .A4(new_n982), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n667), .B(new_n804), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n734), .A2(new_n1011), .A3(KEYINPUT111), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT111), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n718), .A2(new_n1012), .A3(new_n729), .A4(new_n732), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1004), .A2(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n733), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n683), .B(KEYINPUT41), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n736), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n978), .B1(new_n1001), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(G387));
  AOI22_X1  g0823(.A1(new_n785), .A2(G322), .B1(G303), .B2(new_n761), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n955), .B2(new_n758), .C1(new_n777), .C2(new_n775), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT112), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n750), .A2(G294), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n786), .A2(G283), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n766), .A2(G326), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n251), .B1(new_n827), .B2(G116), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n749), .A2(new_n253), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G150), .B2(new_n766), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n202), .B2(new_n758), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G68), .B2(new_n761), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n427), .B(new_n957), .C1(G159), .C2(new_n756), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n782), .A2(new_n348), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n786), .A2(new_n350), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n743), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n286), .A2(G50), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(G68), .A2(G77), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n686), .A2(new_n1049), .A3(new_n403), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n971), .B1(new_n239), .B2(G45), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n686), .A2(new_n682), .A3(new_n427), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n682), .A2(new_n344), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n794), .B(new_n742), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1047), .A2(new_n805), .A3(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT113), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n664), .B(new_n794), .C1(new_n420), .C2(new_n661), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1058), .A2(new_n1059), .B1(new_n737), .B2(new_n1012), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n734), .A2(new_n1012), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n683), .A3(new_n1015), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(G393));
  NOR2_X1   g0863(.A1(new_n1016), .A2(new_n672), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1006), .A2(new_n1010), .A3(new_n672), .ZN(new_n1065));
  OR3_X1    g0865(.A1(new_n1064), .A2(new_n1065), .A3(new_n736), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n982), .A2(new_n794), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT114), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n795), .B1(new_n304), .B2(new_n226), .C1(new_n249), .C2(new_n971), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(KEYINPUT114), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G68), .A2(new_n750), .B1(new_n766), .B2(G143), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n786), .A2(G77), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n286), .C2(new_n762), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G50), .B2(new_n782), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n288), .A2(new_n755), .B1(new_n758), .B2(new_n966), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1074), .A2(new_n251), .A3(new_n828), .A4(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n427), .B1(new_n212), .B2(new_n769), .C1(new_n775), .C2(new_n780), .ZN(new_n1078));
  INV_X1    g0878(.A(G322), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n762), .A2(new_n824), .B1(new_n765), .B2(new_n1079), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n747), .B(new_n1080), .C1(G283), .C2(new_n750), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n955), .A2(new_n755), .B1(new_n758), .B2(new_n777), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT52), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1077), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT115), .Z(new_n1086));
  AOI21_X1  g0886(.A(new_n805), .B1(new_n1086), .B2(new_n742), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n684), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT116), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1015), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1090), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1066), .B(new_n1088), .C1(new_n1092), .C2(new_n1093), .ZN(G390));
  NAND2_X1  g0894(.A1(new_n818), .A2(G330), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n853), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n717), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n929), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n904), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n727), .A2(new_n661), .A3(new_n813), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n853), .B1(new_n1102), .B2(new_n926), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n814), .A2(new_n926), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n929), .B1(new_n1105), .B2(new_n1097), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n898), .ZN(new_n1107));
  OAI21_X1  g0907(.A(KEYINPUT105), .B1(new_n604), .B2(new_n887), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n895), .A2(new_n890), .A3(new_n896), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT38), .B1(new_n1110), .B2(new_n886), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT39), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n932), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1099), .B(new_n1104), .C1(new_n1106), .C2(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n853), .B(new_n1095), .C1(new_n905), .C2(new_n906), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n925), .B1(new_n730), .B2(new_n813), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1100), .B1(new_n1117), .B2(new_n853), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n931), .A2(new_n933), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1114), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n907), .A2(G330), .A3(new_n620), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n937), .A2(new_n619), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1097), .B1(new_n1096), .B2(new_n717), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1105), .B1(new_n1115), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1102), .A2(new_n926), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1095), .B1(new_n905), .B2(new_n906), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n1098), .C1(new_n1127), .C2(new_n1097), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1123), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1121), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1121), .A2(new_n1129), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n683), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n845), .A2(new_n348), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n758), .A2(new_n212), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n762), .A2(new_n304), .B1(new_n519), .B2(new_n749), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(G294), .C2(new_n766), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n251), .B(new_n831), .C1(G283), .C2(new_n756), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n782), .A2(G107), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1136), .A2(new_n1072), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n750), .A2(G150), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n755), .A2(new_n1142), .B1(new_n769), .B2(new_n966), .ZN(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n251), .B1(new_n765), .B2(new_n1144), .C1(new_n838), .C2(new_n758), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT54), .B(G143), .Z(new_n1147));
  AOI22_X1  g0947(.A1(new_n782), .A2(G137), .B1(new_n761), .B2(new_n1147), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1148), .A2(KEYINPUT117), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(KEYINPUT117), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1146), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n746), .A2(new_n202), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1139), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n738), .B1(new_n1154), .B2(new_n743), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1133), .B(new_n1155), .C1(new_n1119), .C2(new_n792), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n1121), .B2(new_n737), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT119), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1132), .B1(new_n1159), .B2(new_n1160), .ZN(G378));
  NAND2_X1  g0961(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1123), .B1(new_n1121), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n909), .B(G330), .C1(new_n918), .C2(new_n919), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n293), .A2(new_n868), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n300), .B2(new_n340), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1166), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n611), .B(new_n1169), .C1(new_n297), .C2(new_n299), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT55), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1168), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT55), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT56), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1173), .A2(new_n1174), .A3(KEYINPUT56), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n928), .A2(new_n934), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n928), .B2(new_n934), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1165), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1164), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1163), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n683), .B1(new_n1185), .B2(KEYINPUT57), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT57), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1187), .B(new_n1163), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1177), .A2(new_n792), .A3(new_n1178), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n844), .A2(new_n202), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n746), .A2(new_n216), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G283), .B2(new_n766), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n344), .B2(new_n758), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1039), .B(new_n1194), .C1(new_n350), .C2(new_n761), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n427), .A2(new_n259), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n769), .A2(new_n207), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(G116), .C2(new_n756), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1195), .B(new_n1198), .C1(new_n304), .C2(new_n775), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT58), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n258), .A2(new_n259), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT120), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(new_n202), .A3(new_n1196), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(G159), .B2(new_n827), .ZN(new_n1204));
  INV_X1    g1004(.A(G124), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1204), .B1(new_n1205), .B2(new_n765), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT121), .Z(new_n1207));
  OAI22_X1  g1007(.A1(new_n755), .A2(new_n1144), .B1(new_n769), .B2(new_n288), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1147), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(new_n749), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G137), .C2(new_n761), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n1142), .B2(new_n758), .C1(new_n838), .C2(new_n775), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT59), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1200), .B(new_n1203), .C1(new_n1207), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n805), .B1(new_n1214), .B2(new_n742), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1190), .A2(new_n1191), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n737), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1189), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(G375));
  NOR2_X1   g1022(.A1(new_n749), .A2(new_n304), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n762), .A2(new_n344), .B1(new_n765), .B2(new_n780), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G283), .C2(new_n759), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n251), .B(new_n960), .C1(G294), .C2(new_n756), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n782), .A2(G116), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n1045), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n775), .A2(new_n1209), .B1(new_n838), .B2(new_n755), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G137), .B2(new_n759), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT123), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n769), .A2(new_n202), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n749), .A2(new_n966), .B1(new_n765), .B2(new_n1142), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(G150), .C2(new_n761), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(new_n251), .A3(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1228), .B1(new_n1235), .B2(new_n1192), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1236), .A2(new_n742), .B1(new_n207), .B2(new_n844), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n738), .B(new_n1237), .C1(new_n1097), .C2(new_n793), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1162), .B2(new_n737), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1125), .A2(new_n1123), .A3(new_n1128), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT122), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1125), .A2(new_n1123), .A3(KEYINPUT122), .A4(new_n1128), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1129), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1241), .B1(new_n1246), .B2(new_n1019), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1247), .A2(KEYINPUT124), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(KEYINPUT124), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(G381));
  NAND2_X1  g1050(.A1(new_n1132), .A2(new_n1157), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G375), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G384), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1248), .A2(new_n1253), .A3(new_n1022), .A4(new_n1249), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(G390), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1252), .A2(new_n1255), .A3(new_n1258), .ZN(G407));
  NAND2_X1  g1059(.A1(new_n1252), .A2(new_n659), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(G407), .A2(G213), .A3(new_n1260), .ZN(G409));
  OAI211_X1 g1061(.A(G378), .B(new_n1219), .C1(new_n1186), .C2(new_n1188), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1185), .A2(new_n1019), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1219), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1251), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n659), .A2(G213), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1242), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT60), .B1(new_n1273), .B2(new_n1123), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n684), .B(new_n1271), .C1(new_n1272), .C2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1253), .B1(new_n1275), .B2(new_n1241), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1271), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n683), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(G384), .A3(new_n1240), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n659), .A2(G213), .A3(G2897), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1276), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1280), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1269), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT126), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1267), .A2(new_n1268), .A3(new_n1287), .A4(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1288), .A2(KEYINPUT126), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1262), .A2(new_n1266), .B1(G213), .B2(new_n659), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1291), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(new_n1287), .A3(new_n1294), .A4(new_n1289), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1285), .A2(new_n1292), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G390), .A2(new_n1022), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT125), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G393), .A2(G396), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1257), .A3(new_n1299), .ZN(new_n1300));
  OR2_X1    g1100(.A1(G390), .A2(new_n1022), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1297), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1256), .B1(new_n1297), .B2(KEYINPUT125), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1304), .A2(new_n1297), .A3(new_n1301), .A4(new_n1299), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1296), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1283), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1281), .ZN(new_n1309));
  OAI21_X1  g1109(.A(KEYINPUT63), .B1(new_n1309), .B2(new_n1293), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1293), .A2(new_n1287), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1267), .A2(new_n1268), .A3(new_n1287), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1306), .B1(new_n1313), .B2(KEYINPUT63), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1312), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1307), .A2(new_n1316), .ZN(G405));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1306), .A2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1262), .B1(new_n1221), .B2(new_n1251), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1287), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1262), .B(new_n1286), .C1(new_n1221), .C2(new_n1251), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1319), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1306), .B(new_n1318), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1323), .B1(new_n1324), .B2(new_n1325), .ZN(G402));
endmodule


