

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X2 U323 ( .A(n310), .B(n309), .ZN(n557) );
  XNOR2_X1 U324 ( .A(n441), .B(KEYINPUT55), .ZN(n442) );
  XOR2_X1 U325 ( .A(n336), .B(n301), .Z(n291) );
  XOR2_X1 U326 ( .A(n329), .B(KEYINPUT45), .Z(n292) );
  AND2_X1 U327 ( .A1(n354), .A2(n353), .ZN(n293) );
  XOR2_X1 U328 ( .A(KEYINPUT9), .B(G92GAT), .Z(n294) );
  XNOR2_X1 U329 ( .A(n334), .B(KEYINPUT75), .ZN(n335) );
  XNOR2_X1 U330 ( .A(n435), .B(n335), .ZN(n337) );
  INV_X1 U331 ( .A(n375), .ZN(n353) );
  XNOR2_X1 U332 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U333 ( .A(n343), .B(n342), .ZN(n346) );
  NOR2_X1 U334 ( .A1(n425), .A2(n544), .ZN(n569) );
  XNOR2_X1 U335 ( .A(n384), .B(KEYINPUT48), .ZN(n545) );
  XNOR2_X1 U336 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U337 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT64), .B(KEYINPUT80), .Z(n296) );
  XNOR2_X1 U339 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n310) );
  XOR2_X1 U341 ( .A(G29GAT), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U342 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n366) );
  XNOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n299), .B(KEYINPUT81), .ZN(n393) );
  XNOR2_X1 U346 ( .A(n366), .B(n393), .ZN(n308) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .Z(n336) );
  XNOR2_X1 U348 ( .A(G134GAT), .B(G218GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n294), .B(n300), .ZN(n301) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n291), .B(n302), .ZN(n303) );
  XOR2_X1 U352 ( .A(n303), .B(KEYINPUT11), .Z(n306) );
  XNOR2_X1 U353 ( .A(G50GAT), .B(KEYINPUT79), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n304), .B(G162GAT), .ZN(n436) );
  XNOR2_X1 U355 ( .A(n436), .B(KEYINPUT66), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  INV_X1 U358 ( .A(n557), .ZN(n459) );
  XOR2_X1 U359 ( .A(G8GAT), .B(G183GAT), .Z(n385) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G155GAT), .Z(n427) );
  XOR2_X1 U361 ( .A(n385), .B(n427), .Z(n312) );
  NAND2_X1 U362 ( .A1(G231GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U364 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n314) );
  XNOR2_X1 U365 ( .A(KEYINPUT12), .B(KEYINPUT82), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U367 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G127GAT), .Z(n455) );
  XOR2_X1 U369 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n318) );
  XNOR2_X1 U370 ( .A(KEYINPUT85), .B(KEYINPUT83), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n455), .B(n319), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U374 ( .A(G64GAT), .B(G78GAT), .Z(n323) );
  XNOR2_X1 U375 ( .A(G71GAT), .B(G211GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U377 ( .A(n325), .B(n324), .Z(n327) );
  XOR2_X1 U378 ( .A(KEYINPUT73), .B(G1GAT), .Z(n365) );
  XOR2_X1 U379 ( .A(KEYINPUT13), .B(G57GAT), .Z(n344) );
  XNOR2_X1 U380 ( .A(n365), .B(n344), .ZN(n326) );
  XOR2_X1 U381 ( .A(n327), .B(n326), .Z(n554) );
  INV_X1 U382 ( .A(n554), .ZN(n581) );
  XNOR2_X1 U383 ( .A(n557), .B(KEYINPUT36), .ZN(n328) );
  XNOR2_X1 U384 ( .A(KEYINPUT103), .B(n328), .ZN(n585) );
  NOR2_X1 U385 ( .A1(n581), .A2(n585), .ZN(n330) );
  XNOR2_X1 U386 ( .A(KEYINPUT65), .B(KEYINPUT114), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n292), .ZN(n354) );
  XOR2_X1 U388 ( .A(KEYINPUT74), .B(KEYINPUT77), .Z(n332) );
  XNOR2_X1 U389 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n347) );
  XNOR2_X1 U391 ( .A(G106GAT), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n333), .B(G148GAT), .ZN(n435) );
  AND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n343) );
  XOR2_X1 U395 ( .A(G120GAT), .B(G71GAT), .Z(n454) );
  XOR2_X1 U396 ( .A(G64GAT), .B(G92GAT), .Z(n339) );
  XNOR2_X1 U397 ( .A(G176GAT), .B(G204GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n388) );
  XOR2_X1 U399 ( .A(n454), .B(n388), .Z(n341) );
  INV_X1 U400 ( .A(KEYINPUT32), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n344), .B(KEYINPUT76), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n348) );
  NAND2_X1 U403 ( .A1(n347), .A2(n348), .ZN(n352) );
  INV_X1 U404 ( .A(n347), .ZN(n350) );
  INV_X1 U405 ( .A(n348), .ZN(n349) );
  NAND2_X1 U406 ( .A1(n350), .A2(n349), .ZN(n351) );
  NAND2_X1 U407 ( .A1(n352), .A2(n351), .ZN(n375) );
  XOR2_X1 U408 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n356) );
  XNOR2_X1 U409 ( .A(G8GAT), .B(KEYINPUT69), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n374) );
  XOR2_X1 U411 ( .A(G197GAT), .B(G22GAT), .Z(n358) );
  XNOR2_X1 U412 ( .A(G50GAT), .B(G36GAT), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U414 ( .A(G113GAT), .B(G15GAT), .Z(n360) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(G141GAT), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U417 ( .A(n362), .B(n361), .Z(n372) );
  XOR2_X1 U418 ( .A(KEYINPUT72), .B(KEYINPUT68), .Z(n364) );
  XNOR2_X1 U419 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n370) );
  XOR2_X1 U421 ( .A(n366), .B(n365), .Z(n368) );
  NAND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(n548) );
  INV_X1 U427 ( .A(n548), .ZN(n572) );
  NAND2_X1 U428 ( .A1(n293), .A2(n572), .ZN(n383) );
  XOR2_X1 U429 ( .A(n375), .B(KEYINPUT41), .Z(n507) );
  NAND2_X1 U430 ( .A1(n507), .A2(n548), .ZN(n377) );
  XNOR2_X1 U431 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n379) );
  NOR2_X1 U433 ( .A1(n554), .A2(n557), .ZN(n378) );
  NAND2_X1 U434 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n380), .B(KEYINPUT47), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n381), .B(KEYINPUT113), .ZN(n382) );
  NAND2_X1 U437 ( .A1(n383), .A2(n382), .ZN(n384) );
  XOR2_X1 U438 ( .A(KEYINPUT97), .B(n385), .Z(n387) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n389) );
  XOR2_X1 U441 ( .A(n389), .B(n388), .Z(n395) );
  XOR2_X1 U442 ( .A(KEYINPUT91), .B(G218GAT), .Z(n391) );
  XNOR2_X1 U443 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U445 ( .A(G197GAT), .B(n392), .Z(n431) );
  XNOR2_X1 U446 ( .A(n431), .B(n393), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U448 ( .A(KEYINPUT17), .B(KEYINPUT88), .Z(n397) );
  XNOR2_X1 U449 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U451 ( .A(G169GAT), .B(n398), .ZN(n449) );
  XNOR2_X1 U452 ( .A(n399), .B(n449), .ZN(n522) );
  NAND2_X1 U453 ( .A1(n545), .A2(n522), .ZN(n401) );
  XOR2_X1 U454 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n425) );
  XOR2_X1 U456 ( .A(G57GAT), .B(G148GAT), .Z(n403) );
  XNOR2_X1 U457 ( .A(G127GAT), .B(G120GAT), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U459 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n405) );
  XNOR2_X1 U460 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U462 ( .A(n407), .B(n406), .Z(n414) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G155GAT), .Z(n411) );
  XOR2_X1 U464 ( .A(KEYINPUT0), .B(KEYINPUT87), .Z(n409) );
  XNOR2_X1 U465 ( .A(G113GAT), .B(G134GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n452) );
  XNOR2_X1 U467 ( .A(n452), .B(G162GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(G29GAT), .B(n412), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n424) );
  XOR2_X1 U471 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n416) );
  XNOR2_X1 U472 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n422) );
  XOR2_X1 U474 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n418) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n426) );
  XOR2_X1 U477 ( .A(n426), .B(KEYINPUT4), .Z(n420) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U480 ( .A(n422), .B(n421), .Z(n423) );
  XOR2_X1 U481 ( .A(n424), .B(n423), .Z(n475) );
  INV_X1 U482 ( .A(n475), .ZN(n544) );
  XOR2_X1 U483 ( .A(n426), .B(G204GAT), .Z(n429) );
  XNOR2_X1 U484 ( .A(n427), .B(KEYINPUT24), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n440) );
  XOR2_X1 U487 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n433) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U490 ( .A(n434), .B(KEYINPUT90), .Z(n438) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n473) );
  NAND2_X1 U494 ( .A1(n569), .A2(n473), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(KEYINPUT118), .ZN(n458) );
  XOR2_X1 U496 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n444) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U499 ( .A(n445), .B(G176GAT), .Z(n451) );
  XOR2_X1 U500 ( .A(G183GAT), .B(G99GAT), .Z(n447) );
  XNOR2_X1 U501 ( .A(G43GAT), .B(G190GAT), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n453) );
  XOR2_X1 U505 ( .A(n453), .B(n452), .Z(n457) );
  XNOR2_X1 U506 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U507 ( .A(n457), .B(n456), .Z(n534) );
  INV_X1 U508 ( .A(n534), .ZN(n524) );
  NAND2_X1 U509 ( .A1(n458), .A2(n524), .ZN(n566) );
  NOR2_X1 U510 ( .A1(n459), .A2(n566), .ZN(n463) );
  XNOR2_X1 U511 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n461) );
  INV_X1 U512 ( .A(G190GAT), .ZN(n460) );
  NAND2_X1 U513 ( .A1(n548), .A2(n353), .ZN(n464) );
  XNOR2_X1 U514 ( .A(n464), .B(KEYINPUT78), .ZN(n494) );
  NOR2_X1 U515 ( .A1(n581), .A2(n557), .ZN(n465) );
  XNOR2_X1 U516 ( .A(n465), .B(KEYINPUT16), .ZN(n482) );
  XOR2_X1 U517 ( .A(n522), .B(KEYINPUT98), .Z(n466) );
  XOR2_X1 U518 ( .A(KEYINPUT27), .B(n466), .Z(n472) );
  NOR2_X1 U519 ( .A1(n473), .A2(n524), .ZN(n467) );
  XNOR2_X1 U520 ( .A(n467), .B(KEYINPUT26), .ZN(n570) );
  NAND2_X1 U521 ( .A1(n472), .A2(n570), .ZN(n547) );
  NAND2_X1 U522 ( .A1(n524), .A2(n522), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n473), .A2(n468), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT25), .B(n469), .Z(n470) );
  NAND2_X1 U525 ( .A1(n547), .A2(n470), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n471), .A2(n475), .ZN(n481) );
  INV_X1 U527 ( .A(n472), .ZN(n477) );
  XOR2_X1 U528 ( .A(n473), .B(KEYINPUT67), .Z(n474) );
  XOR2_X1 U529 ( .A(KEYINPUT28), .B(n474), .Z(n526) );
  OR2_X1 U530 ( .A1(n475), .A2(n526), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n532) );
  XNOR2_X1 U532 ( .A(KEYINPUT99), .B(n532), .ZN(n478) );
  NOR2_X1 U533 ( .A1(n524), .A2(n478), .ZN(n479) );
  XOR2_X1 U534 ( .A(KEYINPUT100), .B(n479), .Z(n480) );
  NAND2_X1 U535 ( .A1(n481), .A2(n480), .ZN(n491) );
  NAND2_X1 U536 ( .A1(n482), .A2(n491), .ZN(n509) );
  NOR2_X1 U537 ( .A1(n494), .A2(n509), .ZN(n488) );
  NAND2_X1 U538 ( .A1(n544), .A2(n488), .ZN(n483) );
  XNOR2_X1 U539 ( .A(n483), .B(KEYINPUT34), .ZN(n484) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n488), .A2(n522), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U544 ( .A1(n488), .A2(n524), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  XOR2_X1 U546 ( .A(G22GAT), .B(KEYINPUT101), .Z(n490) );
  NAND2_X1 U547 ( .A1(n488), .A2(n526), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .Z(n497) );
  NAND2_X1 U550 ( .A1(n581), .A2(n491), .ZN(n492) );
  NOR2_X1 U551 ( .A1(n585), .A2(n492), .ZN(n493) );
  XNOR2_X1 U552 ( .A(KEYINPUT37), .B(n493), .ZN(n520) );
  NOR2_X1 U553 ( .A1(n520), .A2(n494), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n495), .B(KEYINPUT38), .ZN(n504) );
  NAND2_X1 U555 ( .A1(n504), .A2(n544), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U557 ( .A(KEYINPUT102), .B(n498), .ZN(G1328GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n500) );
  NAND2_X1 U559 ( .A1(n522), .A2(n504), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n504), .A2(n524), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n504), .A2(n526), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n505), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n511) );
  INV_X1 U569 ( .A(n507), .ZN(n560) );
  NOR2_X1 U570 ( .A1(n548), .A2(n560), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n508), .B(KEYINPUT107), .ZN(n519) );
  NOR2_X1 U572 ( .A1(n519), .A2(n509), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n515), .A2(n544), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n512), .Z(G1332GAT) );
  NAND2_X1 U576 ( .A1(n515), .A2(n522), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n515), .A2(n524), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n526), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n518), .Z(G1335GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n527), .A2(n544), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n527), .A2(n522), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n527), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n531) );
  XOR2_X1 U592 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n529) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n545), .A2(n532), .ZN(n533) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n541), .A2(n548), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U601 ( .A1(n541), .A2(n507), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n539) );
  NAND2_X1 U604 ( .A1(n541), .A2(n554), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n557), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n548), .A2(n556), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n553) );
  XOR2_X1 U615 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U616 ( .A1(n556), .A2(n507), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n556), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n572), .A2(n566), .ZN(n559) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n559), .Z(G1348GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n566), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n562) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(KEYINPUT56), .B(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n581), .A2(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT123), .B(n571), .Z(n584) );
  NOR2_X1 U636 ( .A1(n572), .A2(n584), .ZN(n577) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT124), .B(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n353), .A2(n584), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

