//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT26), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  AND3_X1   g006(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT68), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT68), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n214), .A3(new_n211), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT27), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n223), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT28), .A4(new_n220), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT67), .A3(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n213), .A2(new_n215), .A3(new_n224), .A4(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G134gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G127gat), .ZN(new_n230));
  INV_X1    g029(.A(G127gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G134gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT69), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n230), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n234), .B(new_n236), .C1(KEYINPUT1), .C2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n237), .A2(KEYINPUT70), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n241));
  OR2_X1    g040(.A1(G113gat), .A2(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(G113gat), .A2(G120gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n239), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247));
  NAND3_X1  g046(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT23), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n252), .B(new_n254), .C1(new_n208), .C2(new_n209), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n247), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  NOR3_X1   g055(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n248), .ZN(new_n259));
  NAND3_X1  g058(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT24), .B1(new_n211), .B2(new_n261), .ZN(new_n262));
  AOI211_X1 g061(.A(new_n257), .B(new_n259), .C1(new_n260), .C2(new_n262), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n208), .A2(new_n209), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n254), .A4(new_n252), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n256), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n228), .A2(new_n246), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n246), .B1(new_n228), .B2(new_n266), .ZN(new_n268));
  INV_X1    g067(.A(G227gat), .ZN(new_n269));
  INV_X1    g068(.A(G233gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n267), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n202), .B1(new_n273), .B2(KEYINPUT33), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n228), .A2(new_n266), .ZN(new_n275));
  INV_X1    g074(.A(new_n246), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n228), .A2(new_n266), .A3(new_n246), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n271), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT33), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(KEYINPUT71), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G15gat), .B(G43gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n284), .B1(new_n279), .B2(KEYINPUT32), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n274), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n277), .A2(new_n278), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT34), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(new_n288), .A3(new_n272), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n287), .B2(new_n272), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n279), .B(KEYINPUT32), .C1(new_n280), .C2(new_n284), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n292), .B1(new_n293), .B2(new_n286), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G141gat), .B(G148gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(KEYINPUT2), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n299), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n303), .B(new_n302), .C1(new_n298), .C2(KEYINPUT2), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT22), .ZN(new_n310));
  INV_X1    g109(.A(G211gat), .ZN(new_n311));
  INV_X1    g110(.A(G218gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(KEYINPUT29), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n308), .B1(new_n317), .B2(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT78), .ZN(new_n319));
  INV_X1    g118(.A(new_n308), .ZN(new_n320));
  INV_X1    g119(.A(new_n315), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n314), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n320), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n306), .A2(new_n307), .A3(new_n325), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n323), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n330), .A2(new_n316), .B1(G228gat), .B2(G233gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n319), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n329), .A2(KEYINPUT79), .A3(new_n323), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n322), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n326), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n332), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT31), .B(G50gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT77), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n340), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n332), .B(new_n342), .C1(new_n333), .C2(new_n337), .ZN(new_n343));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(G22gat), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n341), .B2(new_n343), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(KEYINPUT75), .B(KEYINPUT30), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n275), .A2(new_n323), .ZN(new_n351));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n228), .B2(new_n266), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n322), .A3(new_n355), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n275), .A2(new_n323), .B1(G226gat), .B2(G233gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n316), .B1(new_n357), .B2(new_n354), .ZN(new_n358));
  XNOR2_X1  g157(.A(G8gat), .B(G36gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(G64gat), .ZN(new_n360));
  INV_X1    g159(.A(G92gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n356), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT74), .A4(new_n362), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n350), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n356), .A2(new_n358), .ZN(new_n368));
  INV_X1    g167(.A(new_n362), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(new_n363), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n297), .A2(new_n348), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT35), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT76), .B1(new_n246), .B2(new_n308), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n320), .A2(new_n377), .A3(new_n238), .A4(new_n245), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT4), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT5), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n308), .A2(KEYINPUT3), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n246), .A3(new_n329), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n246), .A2(new_n308), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n379), .B(new_n382), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n376), .A2(new_n378), .B1(KEYINPUT4), .B2(new_n380), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n276), .A2(KEYINPUT4), .A3(new_n320), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n384), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT5), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n376), .A2(new_n378), .B1(new_n308), .B2(new_n246), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n380), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n388), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT0), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G57gat), .ZN(new_n398));
  INV_X1    g197(.A(G85gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n388), .B(new_n400), .C1(new_n392), .C2(new_n394), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(KEYINPUT6), .A3(new_n401), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OR3_X1    g207(.A1(new_n374), .A2(new_n375), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n375), .B1(new_n374), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n322), .B1(new_n353), .B2(new_n355), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n357), .A2(new_n316), .A3(new_n354), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT37), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT37), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n356), .A2(new_n358), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n369), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT38), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT38), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n414), .A2(new_n419), .A3(new_n369), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n365), .A2(new_n366), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n422), .A3(new_n406), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n348), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT39), .ZN(new_n425));
  INV_X1    g224(.A(new_n379), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n387), .B1(new_n384), .B2(KEYINPUT4), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n425), .B(new_n381), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n380), .B1(new_n429), .B2(new_n379), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n393), .A2(new_n380), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT39), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n428), .B(new_n400), .C1(new_n430), .C2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT40), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n381), .B1(new_n426), .B2(new_n427), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT39), .A3(new_n431), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n437), .A2(KEYINPUT40), .A3(new_n400), .A4(new_n428), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n435), .A2(new_n402), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n439), .B(new_n440), .C1(new_n367), .C2(new_n372), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n435), .A2(new_n402), .A3(new_n438), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT81), .B1(new_n373), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n424), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n346), .A2(new_n347), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n367), .A2(new_n372), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n446), .B2(new_n408), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n286), .A2(new_n293), .ZN(new_n448));
  INV_X1    g247(.A(new_n292), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT36), .A3(new_n294), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n450), .B2(new_n294), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT73), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n452), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n454), .B(new_n456), .C1(new_n295), .C2(new_n296), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n447), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n444), .B1(new_n459), .B2(KEYINPUT80), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT80), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n447), .B(new_n461), .C1(new_n455), .C2(new_n458), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n411), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G113gat), .B(G141gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT11), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(G169gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G197gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n466), .B(new_n204), .ZN(new_n469));
  INV_X1    g268(.A(G197gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n468), .A2(new_n471), .A3(KEYINPUT12), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT12), .B1(new_n468), .B2(new_n471), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G22gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G15gat), .ZN(new_n477));
  INV_X1    g276(.A(G15gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G22gat), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT16), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(G1gat), .ZN(new_n481));
  AOI21_X1  g280(.A(G1gat), .B1(new_n477), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n481), .B1(new_n482), .B2(KEYINPUT83), .ZN(new_n483));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n484), .A2(new_n485), .A3(G1gat), .ZN(new_n486));
  OAI21_X1  g285(.A(G8gat), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(KEYINPUT84), .B(G8gat), .C1(new_n483), .C2(new_n486), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n482), .ZN(new_n492));
  INV_X1    g291(.A(G8gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n481), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(KEYINPUT85), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G29gat), .ZN(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT14), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(G29gat), .B2(G36gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(G43gat), .A2(G50gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(G43gat), .A2(G50gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n508), .A3(new_n505), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n503), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT82), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n503), .A2(new_n507), .A3(KEYINPUT82), .A4(new_n509), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n503), .A2(new_n507), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n512), .A2(KEYINPUT17), .A3(new_n513), .A4(new_n514), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n491), .A3(new_n495), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(KEYINPUT86), .A2(KEYINPUT18), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n521), .B(KEYINPUT13), .Z(new_n525));
  INV_X1    g324(.A(new_n515), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n491), .A2(new_n526), .A3(new_n495), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n526), .B1(new_n491), .B2(new_n495), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n523), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n516), .A2(new_n520), .A3(new_n521), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n475), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n522), .A2(new_n523), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n535), .A2(new_n474), .A3(new_n530), .A4(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G176gat), .ZN(new_n540));
  INV_X1    g339(.A(G204gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT7), .B1(new_n399), .B2(new_n361), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT7), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(G85gat), .A3(G92gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n543), .A2(new_n545), .B1(new_n399), .B2(new_n361), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(KEYINPUT93), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(KEYINPUT93), .B2(new_n548), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G99gat), .ZN(new_n552));
  INV_X1    g351(.A(G106gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n548), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT87), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G57gat), .ZN(new_n566));
  INV_X1    g365(.A(G64gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G57gat), .A2(G64gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n559), .A2(KEYINPUT87), .A3(new_n560), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n563), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT90), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT89), .B1(new_n566), .B2(KEYINPUT88), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT89), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n576), .A3(G57gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n577), .A3(G64gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n565), .A3(new_n561), .ZN(new_n579));
  AOI21_X1  g378(.A(G64gat), .B1(new_n574), .B2(new_n577), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n572), .B(new_n573), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n574), .A2(new_n577), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n567), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n584), .A2(new_n578), .A3(new_n565), .A4(new_n561), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n573), .B1(new_n585), .B2(new_n572), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n558), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT10), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n572), .B1(new_n579), .B2(new_n580), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n556), .A2(KEYINPUT97), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n554), .A2(new_n592), .A3(new_n548), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n551), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT98), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n551), .A2(new_n597), .A3(new_n594), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n590), .A2(new_n596), .A3(new_n557), .A4(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n587), .A2(new_n588), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n582), .B2(new_n586), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n558), .A2(new_n588), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n589), .A2(KEYINPUT90), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(KEYINPUT91), .A3(new_n581), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n587), .B2(new_n599), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n542), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n608), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n600), .B2(new_n606), .ZN(new_n614));
  INV_X1    g413(.A(new_n542), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n614), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n538), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  NAND3_X1  g422(.A1(new_n602), .A2(KEYINPUT21), .A3(new_n605), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n491), .A3(new_n495), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(G183gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n625), .A2(G183gat), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  INV_X1    g429(.A(new_n623), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT21), .B1(new_n604), .B2(new_n581), .ZN(new_n633));
  XNOR2_X1  g432(.A(G127gat), .B(G155gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n633), .A2(new_n635), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n311), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n636), .A2(new_n637), .A3(G211gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n629), .A2(new_n632), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n629), .B2(new_n632), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G190gat), .B(G218gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n518), .A2(new_n519), .A3(new_n558), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n555), .A2(new_n557), .ZN(new_n648));
  AND2_X1   g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n648), .A2(new_n515), .B1(KEYINPUT41), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n646), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G134gat), .B(G162gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT92), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  NAND3_X1  g455(.A1(new_n647), .A2(new_n646), .A3(new_n650), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n652), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT94), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n657), .B1(new_n651), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n647), .A2(new_n650), .A3(KEYINPUT94), .A4(new_n646), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n656), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI211_X1 g464(.A(KEYINPUT95), .B(new_n656), .C1(new_n661), .C2(new_n662), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n658), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n620), .B1(new_n644), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n629), .A2(new_n632), .ZN(new_n669));
  INV_X1    g468(.A(new_n641), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n629), .A2(new_n632), .A3(new_n641), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n667), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(KEYINPUT96), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n463), .A2(new_n619), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n408), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n446), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT99), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n683));
  OAI22_X1  g482(.A1(new_n681), .A2(new_n493), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT42), .B1(new_n681), .B2(new_n682), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n684), .A2(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(new_n677), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n455), .A2(new_n458), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n677), .A2(new_n478), .A3(new_n297), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT100), .ZN(G1326gat));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n445), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  NOR2_X1   g495(.A1(new_n619), .A2(new_n673), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n463), .A2(new_n674), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n497), .A3(new_n408), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n463), .B2(new_n674), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n409), .B(new_n410), .C1(new_n459), .C2(new_n444), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n667), .ZN(new_n705));
  AOI211_X1 g504(.A(KEYINPUT101), .B(new_n698), .C1(new_n702), .C2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n459), .A2(KEYINPUT80), .ZN(new_n708));
  INV_X1    g507(.A(new_n444), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n462), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n411), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n674), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n705), .B1(new_n712), .B2(new_n704), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n707), .B1(new_n713), .B2(new_n697), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n706), .A2(new_n714), .A3(new_n407), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n701), .B1(new_n715), .B2(new_n497), .ZN(G1328gat));
  NOR2_X1   g515(.A1(new_n706), .A2(new_n714), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n498), .B1(new_n717), .B2(new_n446), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n719));
  AOI21_X1  g518(.A(G36gat), .B1(new_n719), .B2(KEYINPUT46), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n699), .A2(new_n446), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n719), .A2(KEYINPUT46), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT103), .B1(new_n718), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n706), .A2(new_n714), .A3(new_n373), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n723), .B(new_n726), .C1(new_n727), .C2(new_n498), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(new_n699), .ZN(new_n730));
  INV_X1    g529(.A(new_n297), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n730), .A2(G43gat), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n697), .ZN(new_n734));
  OAI21_X1  g533(.A(G43gat), .B1(new_n734), .B2(new_n689), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n735), .A3(KEYINPUT47), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n717), .A2(new_n688), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n732), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g538(.A1(new_n699), .A2(KEYINPUT105), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n699), .A2(KEYINPUT105), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n348), .A2(G50gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G50gat), .B1(new_n734), .B2(new_n348), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(new_n744), .A3(KEYINPUT48), .ZN(new_n745));
  INV_X1    g544(.A(new_n743), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n717), .A2(new_n445), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(G50gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n749));
  OAI21_X1  g548(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(G1331gat));
  INV_X1    g549(.A(new_n617), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n676), .A2(new_n537), .A3(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(new_n703), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n408), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n446), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT49), .B(G64gat), .Z(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT106), .ZN(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n753), .A2(new_n761), .A3(new_n297), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n753), .A2(new_n688), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(new_n761), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g564(.A1(new_n753), .A2(new_n445), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g566(.A1(new_n673), .A2(new_n537), .A3(new_n751), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n713), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n407), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n673), .A2(new_n537), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n703), .A2(new_n667), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT51), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n751), .A2(new_n407), .A3(G85gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT107), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n773), .B2(new_n775), .ZN(G1336gat));
  INV_X1    g575(.A(new_n769), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n361), .B1(new_n777), .B2(new_n446), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n783));
  OR3_X1    g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n772), .A2(new_n780), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n373), .A2(new_n751), .A3(G92gat), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n778), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  INV_X1    g589(.A(new_n788), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n773), .B2(new_n791), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n789), .A2(new_n790), .B1(new_n778), .B2(new_n792), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n769), .B2(new_n689), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n773), .A2(new_n751), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n297), .A2(new_n552), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(G1338gat));
  AOI21_X1  g596(.A(new_n553), .B1(new_n777), .B2(new_n445), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n445), .A2(new_n553), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n751), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n798), .B1(new_n787), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n795), .B2(new_n799), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n801), .A2(new_n802), .B1(new_n798), .B2(new_n803), .ZN(G1339gat));
  NAND3_X1  g603(.A1(new_n600), .A2(new_n606), .A3(new_n613), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n609), .A2(KEYINPUT54), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n542), .B1(new_n614), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n616), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT55), .B1(new_n806), .B2(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n468), .A2(new_n471), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n528), .A2(new_n529), .A3(new_n525), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n521), .B1(new_n516), .B2(new_n520), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n536), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n667), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n600), .A2(new_n606), .A3(new_n613), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n614), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n607), .A2(new_n608), .A3(new_n807), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n615), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n820), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n537), .A2(new_n826), .A3(new_n810), .A4(new_n809), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n536), .B(new_n816), .C1(new_n612), .C2(new_n616), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT111), .B(new_n819), .C1(new_n829), .C2(new_n667), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n831));
  INV_X1    g630(.A(new_n819), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n667), .B1(new_n827), .B2(new_n828), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n834), .A3(new_n644), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n537), .A2(new_n617), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n668), .A2(new_n675), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n348), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT112), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n446), .A2(new_n407), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n297), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n538), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n838), .A2(new_n408), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n374), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n538), .A2(G113gat), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT113), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n848), .ZN(G1340gat));
  OAI21_X1  g648(.A(G120gat), .B1(new_n842), .B2(new_n751), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n751), .A2(G120gat), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT114), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(G1341gat));
  OAI21_X1  g653(.A(G127gat), .B1(new_n842), .B2(new_n644), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n845), .A2(new_n231), .A3(new_n673), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  NAND3_X1  g656(.A1(new_n845), .A2(new_n229), .A3(new_n667), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT56), .Z(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n842), .B2(new_n674), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1343gat));
  AOI21_X1  g660(.A(new_n348), .B1(new_n835), .B2(new_n837), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT116), .B1(new_n823), .B2(new_n825), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n806), .A2(new_n866), .A3(new_n808), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n820), .A3(new_n867), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n868), .A2(new_n537), .A3(new_n811), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n828), .B(KEYINPUT115), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n674), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n673), .B1(new_n871), .B2(new_n819), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n668), .A2(new_n675), .A3(new_n836), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n445), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT57), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n688), .A2(new_n407), .A3(new_n446), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n864), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G141gat), .B1(new_n877), .B2(new_n538), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n689), .A2(new_n445), .A3(new_n373), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n844), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n838), .A2(KEYINPUT119), .A3(new_n408), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n538), .A2(G141gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n878), .A2(new_n879), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n828), .B(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n868), .A2(new_n537), .A3(new_n811), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n667), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n644), .B1(new_n890), .B2(new_n832), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n348), .B1(new_n891), .B2(new_n837), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n876), .B1(new_n892), .B2(new_n863), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT57), .B(new_n348), .C1(new_n835), .C2(new_n837), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT117), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n864), .A2(new_n875), .A3(new_n896), .A4(new_n876), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n897), .A3(new_n537), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(G141gat), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n898), .B2(G141gat), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n882), .A2(KEYINPUT120), .A3(new_n883), .A4(new_n884), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n886), .B1(new_n906), .B2(new_n879), .ZN(G1344gat));
  NAND3_X1  g706(.A1(new_n895), .A2(new_n897), .A3(new_n617), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(G148gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n908), .A2(KEYINPUT121), .A3(new_n909), .A4(G148gat), .ZN(new_n913));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n892), .A2(new_n863), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n915), .B(new_n617), .C1(new_n863), .C2(new_n862), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n917), .B2(new_n876), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n912), .B(new_n913), .C1(new_n909), .C2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n882), .A2(new_n883), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n914), .A3(new_n617), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n922), .ZN(G1345gat));
  NAND2_X1  g722(.A1(new_n895), .A2(new_n897), .ZN(new_n924));
  OAI21_X1  g723(.A(G155gat), .B1(new_n924), .B2(new_n644), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n300), .A3(new_n673), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n924), .B2(new_n674), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n921), .A2(new_n301), .A3(new_n667), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n408), .A2(new_n373), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n840), .A2(new_n297), .A3(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(new_n204), .A3(new_n538), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n408), .B1(new_n835), .B2(new_n837), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n731), .A2(new_n445), .A3(new_n373), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT122), .Z(new_n937));
  AOI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n537), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n933), .A2(new_n938), .ZN(G1348gat));
  OAI21_X1  g738(.A(G176gat), .B1(new_n932), .B2(new_n751), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n205), .A3(new_n617), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1349gat));
  OAI21_X1  g741(.A(G183gat), .B1(new_n932), .B2(new_n644), .ZN(new_n943));
  AND2_X1   g742(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n944));
  INV_X1    g743(.A(new_n936), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n945), .A2(new_n217), .A3(new_n219), .A4(new_n673), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n937), .A2(new_n220), .A3(new_n667), .ZN(new_n950));
  OAI21_X1  g749(.A(G190gat), .B1(new_n932), .B2(new_n674), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(KEYINPUT61), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n953), .B(G190gat), .C1(new_n932), .C2(new_n674), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n950), .B1(new_n952), .B2(new_n955), .ZN(G1351gat));
  NOR3_X1   g755(.A1(new_n688), .A2(new_n348), .A3(new_n373), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n934), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n470), .A3(new_n537), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n689), .A2(new_n931), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n915), .B(new_n962), .C1(new_n863), .C2(new_n862), .ZN(new_n963));
  OAI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n538), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n960), .A2(new_n964), .ZN(G1352gat));
  NAND3_X1  g764(.A1(new_n958), .A2(new_n541), .A3(new_n617), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT62), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n541), .B1(new_n917), .B2(new_n962), .ZN(new_n969));
  OR3_X1    g768(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1353gat));
  OAI21_X1  g771(.A(G211gat), .B1(new_n963), .B2(new_n644), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(KEYINPUT126), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n958), .A2(new_n311), .A3(new_n673), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n977), .B(new_n978), .C1(KEYINPUT126), .C2(new_n976), .ZN(G1354gat));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n674), .B1(new_n963), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n981), .B1(new_n980), .B2(new_n963), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G218gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n958), .A2(new_n312), .A3(new_n667), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


