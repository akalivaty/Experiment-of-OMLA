//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n585, new_n587, new_n588,
    new_n589, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n644, new_n645, new_n647,
    new_n648, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1243, new_n1244, new_n1245;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(KEYINPUT67), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  NAND3_X1  g048(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G137), .B1(G101), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n470), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G100), .ZN(new_n481));
  NAND2_X1  g056(.A1(G112), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n463), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n475), .A2(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n480), .B1(new_n473), .B2(new_n474), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n483), .B(new_n484), .C1(G124), .C2(new_n485), .ZN(G162));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n473), .B2(new_n474), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT69), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n463), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT4), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n473), .B2(new_n474), .ZN(new_n496));
  AND2_X1   g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n480), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(G138), .A3(new_n480), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n494), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XOR2_X1   g086(.A(KEYINPUT71), .B(G88), .Z(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n507), .B2(new_n508), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(KEYINPUT72), .A2(G75), .A3(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(G651), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n521), .A2(new_n522), .ZN(new_n527));
  AND3_X1   g102(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(G543), .B1(KEYINPUT70), .B2(KEYINPUT5), .ZN(new_n529));
  OAI21_X1  g104(.A(G62), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(KEYINPUT73), .A3(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n516), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(KEYINPUT74), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  AOI211_X1 g110(.A(new_n535), .B(new_n516), .C1(new_n526), .C2(new_n532), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  NAND2_X1  g113(.A1(new_n507), .A2(new_n508), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(KEYINPUT6), .A2(G651), .ZN(new_n544));
  NOR2_X1   g119(.A1(KEYINPUT6), .A2(G651), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n528), .A2(new_n529), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G89), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(G543), .B1(new_n544), .B2(new_n545), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g127(.A(KEYINPUT75), .B(G543), .C1(new_n544), .C2(new_n545), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G51), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n549), .A2(new_n555), .ZN(G286));
  INV_X1    g131(.A(G286), .ZN(G168));
  AOI22_X1  g132(.A1(new_n554), .A2(G52), .B1(G90), .B2(new_n511), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n559));
  INV_X1    g134(.A(G64), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n507), .B2(new_n508), .ZN(new_n561));
  NAND2_X1  g136(.A1(G77), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n559), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n528), .A2(new_n529), .ZN(new_n565));
  OAI211_X1 g140(.A(KEYINPUT76), .B(new_n562), .C1(new_n565), .C2(new_n560), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n566), .A3(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n558), .A2(new_n567), .ZN(G301));
  INV_X1    g143(.A(G301), .ZN(G171));
  NAND2_X1  g144(.A1(new_n509), .A2(new_n510), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT75), .B1(new_n570), .B2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n553), .ZN(new_n572));
  OAI21_X1  g147(.A(G43), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G651), .ZN(new_n574));
  OAI21_X1  g149(.A(G56), .B1(new_n528), .B2(new_n529), .ZN(new_n575));
  NAND2_X1  g150(.A1(G68), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  XOR2_X1   g153(.A(KEYINPUT77), .B(G81), .Z(new_n579));
  NOR2_X1   g154(.A1(new_n546), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n573), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G860), .ZN(G153));
  AND3_X1   g159(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G36), .ZN(G176));
  NAND2_X1  g161(.A1(G1), .A2(G3), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT78), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT8), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G188));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n591));
  INV_X1    g166(.A(G65), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n507), .B2(new_n508), .ZN(new_n593));
  NAND2_X1  g168(.A1(G78), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n591), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g171(.A(KEYINPUT79), .B(new_n594), .C1(new_n565), .C2(new_n592), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n596), .A2(new_n597), .A3(G651), .ZN(new_n598));
  INV_X1    g173(.A(G53), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT9), .B1(new_n550), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT9), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n570), .A2(new_n601), .A3(G53), .A4(G543), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n600), .A2(new_n602), .B1(G91), .B2(new_n511), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n598), .A2(new_n603), .ZN(G299));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n605));
  INV_X1    g180(.A(G87), .ZN(new_n606));
  INV_X1    g181(.A(G49), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n546), .A2(new_n606), .B1(new_n550), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G74), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n574), .B1(new_n565), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n605), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n511), .A2(G87), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n539), .B2(G74), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n514), .A2(G49), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n612), .A2(KEYINPUT80), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(G288));
  AOI22_X1  g192(.A1(new_n511), .A2(G86), .B1(new_n514), .B2(G48), .ZN(new_n618));
  INV_X1    g193(.A(G61), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n507), .B2(new_n508), .ZN(new_n620));
  AND2_X1   g195(.A1(G73), .A2(G543), .ZN(new_n621));
  OAI21_X1  g196(.A(G651), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(G305));
  NAND2_X1  g198(.A1(new_n554), .A2(G47), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT81), .B(G85), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n511), .A2(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n539), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n626), .C1(new_n574), .C2(new_n627), .ZN(G290));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n629));
  INV_X1    g204(.A(G92), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n546), .B2(new_n630), .ZN(new_n631));
  NAND4_X1  g206(.A1(new_n539), .A2(new_n570), .A3(KEYINPUT10), .A4(G92), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(G54), .B1(new_n571), .B2(new_n572), .ZN(new_n634));
  NAND2_X1  g209(.A1(G79), .A2(G543), .ZN(new_n635));
  INV_X1    g210(.A(G66), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n565), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G651), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  MUX2_X1   g214(.A(new_n639), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g215(.A(new_n639), .B(G301), .S(G868), .Z(G321));
  MUX2_X1   g216(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g217(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g218(.A(new_n639), .ZN(new_n644));
  INV_X1    g219(.A(G559), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(G860), .ZN(G148));
  NOR2_X1   g221(.A1(new_n582), .A2(G868), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n639), .A2(G559), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n647), .B1(new_n648), .B2(G868), .ZN(G323));
  XNOR2_X1  g224(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n653), .B(new_n654), .C1(G111), .C2(new_n480), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n485), .A2(G123), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n475), .A2(G135), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n480), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT12), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT13), .ZN(new_n663));
  INV_X1    g238(.A(G2100), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n660), .A2(new_n665), .A3(new_n666), .ZN(G156));
  INV_X1    g242(.A(KEYINPUT14), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT15), .B(G2435), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2438), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2427), .ZN(new_n671));
  INV_X1    g246(.A(G2430), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2451), .B(G2454), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT16), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2443), .B(G2446), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1341), .B(G1348), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n674), .A2(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(G14), .A3(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G401));
  XNOR2_X1  g259(.A(G2072), .B(G2078), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2084), .B(G2090), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2067), .B(G2678), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT83), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT18), .ZN(new_n693));
  INV_X1    g268(.A(new_n685), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(new_n691), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n693), .B1(new_n695), .B2(new_n688), .ZN(new_n696));
  OR4_X1    g271(.A1(new_n693), .A2(new_n694), .A3(new_n691), .A4(new_n688), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n690), .A2(new_n692), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(new_n694), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(new_n688), .C1(new_n692), .C2(new_n687), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(new_n659), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(new_n664), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G227));
  XNOR2_X1  g279(.A(G1961), .B(G1966), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT86), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT86), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1956), .B(G2474), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT85), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1971), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT19), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n707), .A3(new_n706), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n713), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n714), .A2(KEYINPUT20), .A3(new_n713), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n715), .B1(new_n713), .B2(new_n711), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(G1991), .B(G1996), .ZN(new_n723));
  XNOR2_X1  g298(.A(G1981), .B(G1986), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n722), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(G229));
  NAND2_X1  g304(.A1(G303), .A2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G22), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT91), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G1971), .ZN(new_n735));
  INV_X1    g310(.A(G1971), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n730), .A2(new_n736), .A3(new_n733), .ZN(new_n737));
  NOR2_X1   g312(.A1(G6), .A2(G16), .ZN(new_n738));
  INV_X1    g313(.A(G305), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT32), .B(G1981), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n740), .B(new_n741), .Z(new_n742));
  NOR2_X1   g317(.A1(G16), .A2(G23), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT90), .Z(new_n744));
  NOR2_X1   g319(.A1(new_n608), .A2(new_n610), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n744), .B1(new_n746), .B2(new_n731), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT33), .B(G1976), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n747), .B(new_n748), .Z(new_n749));
  NAND4_X1  g324(.A1(new_n735), .A2(new_n737), .A3(new_n742), .A4(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(KEYINPUT34), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(KEYINPUT34), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n731), .A2(G24), .ZN(new_n753));
  XOR2_X1   g328(.A(G290), .B(KEYINPUT89), .Z(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(new_n731), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1986), .Z(new_n756));
  XOR2_X1   g331(.A(KEYINPUT87), .B(G29), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G25), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n475), .A2(G131), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n485), .A2(G119), .ZN(new_n760));
  AND2_X1   g335(.A1(G107), .A2(G2105), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G95), .B2(new_n480), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n759), .B(new_n760), .C1(new_n463), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT88), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(new_n757), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT35), .B(G1991), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n751), .A2(new_n752), .A3(new_n756), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT36), .ZN(new_n769));
  INV_X1    g344(.A(new_n757), .ZN(new_n770));
  NAND2_X1  g345(.A1(G162), .A2(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(G35), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT29), .ZN(new_n774));
  INV_X1    g349(.A(G2090), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G168), .A2(new_n731), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n731), .B2(G21), .ZN(new_n778));
  INV_X1    g353(.A(G1966), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n658), .A2(new_n757), .ZN(new_n782));
  OR2_X1    g357(.A1(KEYINPUT30), .A2(G28), .ZN(new_n783));
  NAND2_X1  g358(.A1(KEYINPUT30), .A2(G28), .ZN(new_n784));
  AOI21_X1  g359(.A(G29), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT31), .B(G11), .Z(new_n786));
  NOR3_X1   g361(.A1(new_n782), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n776), .A2(new_n780), .A3(new_n781), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n770), .A2(G27), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G164), .B2(new_n770), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n774), .B2(new_n775), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT25), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n475), .A2(G139), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n796), .B(new_n797), .C1(new_n480), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G29), .ZN(new_n801));
  NOR2_X1   g376(.A1(G29), .A2(G33), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT92), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G2072), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n731), .A2(G20), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT23), .Z(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G299), .B2(G16), .ZN(new_n808));
  INV_X1    g383(.A(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(KEYINPUT24), .A2(G34), .ZN(new_n811));
  AND2_X1   g386(.A1(KEYINPUT24), .A2(G34), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n757), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G29), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n478), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT94), .ZN(new_n816));
  INV_X1    g391(.A(G2084), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n805), .A2(new_n810), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n814), .A2(G32), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n485), .A2(G129), .ZN(new_n821));
  NAND3_X1  g396(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT95), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT26), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n475), .A2(G141), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n821), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n823), .A2(new_n824), .B1(G105), .B2(new_n476), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n820), .B1(new_n830), .B2(new_n814), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT27), .B(G1996), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT96), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n757), .A2(G26), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT28), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n475), .A2(G140), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n485), .A2(G128), .ZN(new_n838));
  MUX2_X1   g413(.A(G104), .B(G116), .S(G2105), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G2104), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n836), .B1(new_n841), .B2(G29), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G2067), .ZN(new_n843));
  NOR2_X1   g418(.A1(G4), .A2(G16), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n644), .B2(G16), .ZN(new_n845));
  INV_X1    g420(.A(G1348), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(G16), .A2(G19), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n583), .B2(G16), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(G1341), .Z(new_n850));
  NAND4_X1  g425(.A1(new_n834), .A2(new_n843), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n731), .A2(G5), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(G171), .B2(new_n731), .ZN(new_n853));
  INV_X1    g428(.A(G1961), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n816), .B2(new_n817), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n794), .A2(new_n819), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n769), .A2(new_n860), .ZN(G311));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n769), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n769), .B2(new_n860), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(G150));
  NAND2_X1  g440(.A1(new_n644), .A2(G559), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n580), .B1(new_n554), .B2(G43), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT100), .B1(new_n868), .B2(new_n578), .ZN(new_n869));
  INV_X1    g444(.A(G43), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n552), .B2(new_n553), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  NOR4_X1   g447(.A1(new_n871), .A2(new_n577), .A3(new_n580), .A4(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G55), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n552), .B2(new_n553), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n539), .A2(G67), .ZN(new_n876));
  NAND2_X1  g451(.A1(G80), .A2(G543), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n574), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT99), .B(G93), .Z(new_n879));
  NOR2_X1   g454(.A1(new_n546), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n875), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n869), .A2(new_n873), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n875), .A2(new_n880), .ZN(new_n883));
  INV_X1    g458(.A(new_n878), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n582), .A2(new_n872), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n868), .A2(KEYINPUT100), .A3(new_n578), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n867), .B(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n890), .A2(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(KEYINPUT39), .ZN(new_n892));
  XNOR2_X1  g467(.A(KEYINPUT101), .B(G860), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n881), .A2(new_n893), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(G145));
  OR2_X1    g472(.A1(new_n763), .A2(new_n662), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n475), .A2(G142), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n485), .A2(G130), .ZN(new_n900));
  MUX2_X1   g475(.A(G106), .B(G118), .S(G2105), .Z(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G2104), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n763), .A2(new_n662), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n898), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n503), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n498), .A2(new_n494), .A3(new_n502), .A4(KEYINPUT102), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n841), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n841), .B1(new_n909), .B2(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n830), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n829), .A3(new_n911), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n916), .A3(new_n799), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT103), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n829), .B1(new_n915), .B2(new_n911), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n912), .A2(new_n830), .A3(new_n913), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n800), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n914), .A2(new_n916), .A3(new_n923), .A4(new_n799), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n907), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G162), .B(G160), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(new_n658), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n907), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT104), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(new_n918), .A3(new_n924), .A4(new_n922), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n926), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(KEYINPUT105), .B(G37), .Z(new_n936));
  AND2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n919), .A2(new_n925), .B1(new_n931), .B2(new_n932), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n929), .B1(new_n938), .B2(new_n934), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g517(.A1(new_n885), .A2(G868), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n889), .B(new_n648), .ZN(new_n944));
  NAND2_X1  g519(.A1(G299), .A2(new_n639), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n554), .A2(G54), .B1(new_n637), .B2(G651), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n598), .A3(new_n603), .A4(new_n633), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n947), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n949), .A2(KEYINPUT107), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n950), .A2(KEYINPUT107), .A3(new_n952), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n944), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n950), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n944), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT42), .ZN(new_n960));
  XNOR2_X1  g535(.A(G290), .B(new_n746), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n513), .A2(new_n515), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT73), .B1(new_n531), .B2(G651), .ZN(new_n964));
  AOI211_X1 g539(.A(new_n525), .B(new_n574), .C1(new_n527), .C2(new_n530), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n535), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n533), .A2(KEYINPUT74), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n739), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n739), .B1(new_n967), .B2(new_n968), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(G305), .B1(new_n534), .B2(new_n536), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(new_n961), .A3(new_n969), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n960), .B(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n943), .B1(new_n976), .B2(G868), .ZN(G295));
  AOI21_X1  g552(.A(new_n943), .B1(new_n976), .B2(G868), .ZN(G331));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g554(.A1(G301), .A2(G286), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n558), .A2(new_n549), .A3(new_n555), .A4(new_n567), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n882), .A2(new_n982), .A3(new_n888), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n881), .B1(new_n869), .B2(new_n873), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n886), .A2(new_n885), .A3(new_n887), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n984), .A2(new_n985), .B1(new_n980), .B2(new_n981), .ZN(new_n986));
  OAI22_X1  g561(.A1(new_n983), .A2(new_n986), .B1(new_n953), .B2(new_n954), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n982), .B1(new_n882), .B2(new_n888), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n984), .A2(new_n985), .A3(new_n980), .A4(new_n981), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n957), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n973), .A2(new_n961), .A3(new_n969), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n961), .B1(new_n973), .B2(new_n969), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n949), .A2(KEYINPUT107), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n950), .A2(new_n952), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n950), .A2(KEYINPUT107), .A3(new_n952), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n998), .A2(new_n999), .B1(new_n988), .B2(new_n989), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n988), .A2(new_n957), .A3(new_n989), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT108), .B1(new_n1002), .B2(new_n975), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n975), .A2(new_n987), .A3(KEYINPUT108), .A4(new_n990), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n995), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(KEYINPUT43), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n945), .A2(new_n947), .A3(new_n952), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n957), .B2(KEYINPUT41), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n988), .B2(new_n989), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n994), .B1(new_n1011), .B2(new_n1001), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n936), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n991), .B2(new_n994), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1013), .B1(new_n1015), .B2(new_n1004), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1008), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1004), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1020), .B2(new_n995), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(new_n1007), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n979), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT110), .ZN(new_n1024));
  INV_X1    g599(.A(G37), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n1002), .B2(new_n975), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1015), .B2(new_n1004), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT109), .B1(new_n1027), .B2(new_n1017), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(new_n1008), .A3(new_n1018), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n979), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n979), .B1(new_n1027), .B2(new_n1017), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(new_n1031), .A3(new_n1033), .ZN(G397));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n909), .A2(new_n910), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(G1384), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n470), .A2(G40), .A3(new_n471), .A4(new_n477), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1040), .A2(G1996), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n841), .A2(G2067), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n841), .A2(G2067), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n1041), .A2(new_n829), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1039), .A2(G1996), .A3(new_n829), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT111), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n763), .B(new_n766), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G290), .B(G1986), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1039), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1038), .ZN(new_n1053));
  INV_X1    g628(.A(G1384), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n503), .A2(KEYINPUT50), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT50), .B1(new_n503), .B2(new_n1054), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1053), .B(new_n775), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n503), .A2(new_n1054), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1038), .B1(new_n1059), .B2(new_n1035), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n909), .A2(KEYINPUT45), .A3(new_n1054), .A4(new_n910), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1971), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n967), .A2(new_n968), .A3(G8), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n967), .A2(new_n968), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT113), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT112), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1063), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1059), .A2(new_n1038), .ZN(new_n1077));
  INV_X1    g652(.A(G1981), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n622), .B2(KEYINPUT116), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G305), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n618), .B(new_n622), .C1(KEYINPUT116), .C2(new_n1078), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(KEYINPUT49), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1077), .A2(G8), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT49), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n745), .A2(G1976), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(G8), .C1(new_n1059), .C2(new_n1038), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1083), .A2(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1976), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n611), .A2(new_n1090), .A3(new_n615), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1088), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT114), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1094), .A3(new_n1088), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1087), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT115), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1087), .A2(new_n1093), .A3(new_n1098), .A4(new_n1095), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1089), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1076), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1102), .A2(G1976), .A3(G288), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G305), .A2(G1981), .ZN(new_n1104));
  OAI211_X1 g679(.A(G8), .B(new_n1077), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1063), .A2(new_n1073), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G8), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1059), .B2(new_n1035), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n503), .A2(KEYINPUT117), .A3(KEYINPUT45), .A4(new_n1054), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1060), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n779), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1056), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n503), .A2(KEYINPUT50), .A3(new_n1054), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1038), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n817), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1109), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G168), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1076), .A2(new_n1108), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT63), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1120), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1124), .B(new_n1125), .C1(new_n1126), .C2(new_n1063), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(KEYINPUT118), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1106), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G8), .ZN(new_n1132));
  NAND2_X1  g707(.A1(G286), .A2(G8), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT51), .B1(new_n1119), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1132), .A2(new_n1135), .A3(KEYINPUT51), .A4(new_n1133), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1119), .A2(G286), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n854), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1143), .A2(G2078), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1113), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1060), .A2(new_n1061), .A3(new_n791), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1147), .A2(new_n1143), .ZN(new_n1148));
  OAI21_X1  g723(.A(G171), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1143), .ZN(new_n1150));
  AND4_X1   g725(.A1(G40), .A2(new_n477), .A3(new_n468), .A4(new_n1144), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1037), .A2(new_n1061), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(new_n1152), .A3(new_n1142), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1149), .B1(G171), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n1155));
  OR3_X1    g730(.A1(new_n1146), .A2(new_n1148), .A3(G171), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1153), .B2(G171), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1154), .A2(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1076), .A2(new_n1108), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1140), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1141), .A2(new_n809), .ZN(new_n1162));
  XNOR2_X1  g737(.A(G299), .B(KEYINPUT57), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(KEYINPUT56), .B(G2072), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1060), .A2(new_n1061), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1164), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(new_n1168), .B2(KEYINPUT121), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1170), .A2(KEYINPUT121), .A3(new_n1163), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1161), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1163), .B(KEYINPUT119), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1170), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(KEYINPUT61), .A3(new_n1167), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1059), .A2(new_n1038), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT58), .B(G1341), .Z(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT120), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1176), .A2(G1996), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1180), .A2(KEYINPUT59), .A3(new_n583), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT59), .B1(new_n1180), .B2(new_n583), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1172), .A2(new_n1175), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(G2067), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1177), .A2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(KEYINPUT60), .B(new_n1186), .C1(new_n1117), .C2(G1348), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT122), .B1(new_n1187), .B2(new_n644), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1141), .A2(new_n846), .B1(new_n1185), .B2(new_n1177), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1189), .A2(new_n1190), .A3(KEYINPUT60), .A4(new_n639), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1187), .A2(new_n644), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1188), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1189), .A2(KEYINPUT60), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(KEYINPUT123), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1193), .A2(new_n1197), .A3(new_n1194), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1184), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1189), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1200), .A2(new_n1167), .A3(new_n644), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1174), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1160), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1130), .A2(new_n1203), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1076), .A2(new_n1108), .A3(new_n1149), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1137), .A2(new_n1206), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  AND2_X1   g783(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1206), .B1(new_n1209), .B2(new_n1137), .ZN(new_n1210));
  OAI21_X1  g785(.A(KEYINPUT125), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1140), .A2(KEYINPUT62), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1212), .A2(new_n1213), .A3(new_n1207), .A4(new_n1205), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1052), .B1(new_n1204), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1217), .A2(KEYINPUT46), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1217), .A2(KEYINPUT46), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1218), .B1(new_n1041), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1044), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1039), .B1(new_n829), .B2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g797(.A(new_n1220), .B(new_n1222), .C1(new_n1041), .C2(new_n1218), .ZN(new_n1223));
  XOR2_X1   g798(.A(new_n1223), .B(KEYINPUT47), .Z(new_n1224));
  NAND3_X1  g799(.A1(new_n1048), .A2(new_n764), .A3(new_n766), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1040), .B1(new_n1225), .B2(new_n1042), .ZN(new_n1226));
  NOR3_X1   g801(.A1(new_n1040), .A2(G1986), .A3(G290), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1227), .B(KEYINPUT48), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n1050), .A2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g804(.A1(new_n1224), .A2(new_n1226), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1216), .A2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g806(.A1(new_n703), .A2(G319), .A3(new_n683), .ZN(new_n1233));
  AOI21_X1  g807(.A(new_n1233), .B1(new_n727), .B2(new_n726), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n935), .A2(new_n936), .ZN(new_n1235));
  OAI21_X1  g809(.A(new_n1234), .B1(new_n1235), .B2(new_n939), .ZN(new_n1236));
  AOI22_X1  g810(.A1(new_n1021), .A2(new_n1007), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1237));
  AOI211_X1 g811(.A(KEYINPUT127), .B(new_n1236), .C1(new_n1237), .C2(new_n1028), .ZN(new_n1238));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1239));
  INV_X1    g813(.A(new_n1236), .ZN(new_n1240));
  AOI21_X1  g814(.A(new_n1239), .B1(new_n1029), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g815(.A1(new_n1238), .A2(new_n1241), .ZN(G308));
  OAI21_X1  g816(.A(new_n1240), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1243));
  NAND2_X1  g817(.A1(new_n1243), .A2(KEYINPUT127), .ZN(new_n1244));
  NAND3_X1  g818(.A1(new_n1029), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1245));
  NAND2_X1  g819(.A1(new_n1244), .A2(new_n1245), .ZN(G225));
endmodule


