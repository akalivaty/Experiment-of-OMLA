//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G77), .A2(G244), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G68), .A2(G238), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n205), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n208), .B(new_n222), .C1(new_n225), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n223), .ZN(new_n251));
  OR2_X1    g0051(.A1(new_n251), .A2(KEYINPUT69), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(KEYINPUT69), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G50), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n258));
  OAI21_X1  g0058(.A(G20), .B1(new_n228), .B2(G50), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT68), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n263), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n251), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n257), .B1(G50), .B2(new_n258), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT73), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n266), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G222), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n279), .C1(new_n280), .C2(new_n278), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n284), .C1(G77), .C2(new_n277), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n283), .A2(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G226), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n285), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G200), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n273), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT10), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n293), .B2(KEYINPUT74), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n270), .A2(new_n271), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n294), .A2(new_n297), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n273), .A2(new_n293), .A3(new_n301), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n296), .B1(new_n303), .B2(new_n299), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n292), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n270), .B(new_n307), .C1(G179), .C2(new_n292), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G50), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n262), .A2(new_n311), .B1(new_n224), .B2(G68), .ZN(new_n312));
  INV_X1    g0112(.A(G77), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n266), .A2(new_n313), .A3(G20), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n251), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT11), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT71), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n269), .A2(new_n258), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n258), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT71), .B1(new_n319), .B2(new_n251), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G68), .A3(new_n254), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n227), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT12), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n316), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT75), .ZN(new_n326));
  INV_X1    g0126(.A(G226), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n278), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n233), .A2(G1698), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G97), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n326), .B1(new_n334), .B2(new_n283), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(new_n333), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT75), .A3(new_n284), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n288), .B1(new_n290), .B2(G238), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT13), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n335), .A2(new_n337), .A3(new_n341), .A4(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n325), .B1(new_n343), .B2(G200), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(G190), .A3(new_n342), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT76), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n340), .A2(KEYINPUT76), .A3(G190), .A4(new_n342), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT77), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT77), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n344), .A2(new_n347), .A3(new_n351), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n306), .B1(new_n340), .B2(new_n342), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT14), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n340), .A2(G179), .A3(new_n342), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n355), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n325), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n264), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n262), .A2(KEYINPUT70), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT70), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n261), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  XOR2_X1   g0166(.A(KEYINPUT15), .B(G87), .Z(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n267), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n368), .C1(new_n224), .C2(new_n313), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n251), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n319), .A2(new_n313), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n321), .A2(G77), .A3(new_n254), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G238), .A2(G1698), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n277), .B(new_n374), .C1(new_n233), .C2(G1698), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n284), .C1(G107), .C2(new_n277), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n290), .A2(G244), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n289), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n306), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT72), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n378), .A2(G179), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n373), .A2(new_n379), .A3(KEYINPUT72), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n378), .A2(G200), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n378), .A2(new_n298), .ZN(new_n388));
  OR3_X1    g0188(.A1(new_n387), .A2(new_n373), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n361), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n330), .A2(new_n331), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n392), .B2(new_n224), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n224), .A4(new_n276), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G159), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n262), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G58), .A2(G68), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n224), .B1(new_n228), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n275), .A2(new_n224), .A3(new_n276), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n394), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n401), .B1(new_n409), .B2(G68), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT16), .A3(new_n399), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n405), .A2(new_n251), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n280), .A2(new_n278), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n327), .A2(G1698), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(new_n330), .C2(new_n331), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n288), .B1(new_n417), .B2(new_n284), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n283), .A2(G232), .A3(new_n286), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G200), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G190), .B2(new_n421), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n256), .A2(new_n265), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n258), .B2(new_n265), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n412), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n269), .B1(new_n403), .B2(new_n404), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n426), .B1(new_n431), .B2(new_n411), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(KEYINPUT17), .A3(new_n424), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n412), .A2(new_n427), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n306), .B1(new_n418), .B2(new_n420), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n283), .B1(new_n415), .B2(new_n416), .ZN(new_n436));
  INV_X1    g0236(.A(G179), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n436), .A2(new_n437), .A3(new_n419), .A4(new_n288), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT18), .B1(new_n434), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  AOI211_X1 g0242(.A(new_n442), .B(new_n439), .C1(new_n412), .C2(new_n427), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n430), .B(new_n433), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n310), .A2(new_n391), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n258), .A2(G97), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n266), .A2(G1), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n319), .A2(new_n251), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n450), .B2(G97), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G97), .A2(G107), .ZN(new_n455));
  NAND2_X1  g0255(.A1(KEYINPUT6), .A2(G107), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n203), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(G97), .A2(G107), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n452), .B(new_n453), .C1(new_n458), .C2(new_n202), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n224), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n262), .A2(new_n313), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n409), .A2(G107), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n269), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT79), .ZN(new_n466));
  AOI211_X1 g0266(.A(new_n466), .B(new_n269), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n451), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(G244), .B1(new_n330), .B2(new_n331), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n469), .A2(new_n470), .B1(G33), .B2(G283), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .A4(new_n278), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n277), .A2(G250), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n278), .B1(new_n474), .B2(KEYINPUT4), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT80), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n392), .A2(new_n211), .ZN(new_n477));
  OAI21_X1  g0277(.A(G1698), .B1(new_n477), .B2(new_n470), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n471), .A4(new_n472), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n480), .A3(new_n284), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(G274), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n483), .B1(new_n485), .B2(new_n484), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n488), .A2(new_n283), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n487), .B1(new_n489), .B2(G257), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n306), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n481), .A2(new_n437), .A3(new_n490), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n468), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(G200), .ZN(new_n495));
  INV_X1    g0295(.A(new_n451), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n497));
  INV_X1    g0297(.A(G107), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n408), .B2(new_n394), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n499), .A2(new_n460), .A3(new_n461), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n466), .B1(new_n500), .B2(new_n269), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n496), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n481), .A2(G190), .A3(new_n490), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n495), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n494), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n449), .B1(new_n318), .B2(new_n320), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G116), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n319), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(G20), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n251), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT85), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n251), .A2(new_n513), .A3(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(G20), .B1(G33), .B2(G283), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G33), .B2(new_n212), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT20), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n251), .A2(new_n513), .A3(new_n510), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n513), .B1(new_n251), .B2(new_n510), .ZN(new_n520));
  OAI211_X1 g0320(.A(KEYINPUT20), .B(new_n517), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n507), .B(new_n509), .C1(new_n518), .C2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n488), .A2(G270), .A3(new_n283), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT84), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n488), .A2(KEYINPUT84), .A3(G270), .A4(new_n283), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n487), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G264), .A2(G1698), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n277), .B(new_n529), .C1(new_n213), .C2(G1698), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(new_n284), .C1(G303), .C2(new_n277), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n306), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n523), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n531), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT20), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n521), .B1(G116), .B2(new_n506), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n528), .A2(G190), .A3(new_n531), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n537), .A2(new_n509), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n523), .A2(G179), .A3(new_n531), .A4(new_n528), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n523), .A2(KEYINPUT21), .A3(new_n532), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n535), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n547), .B(KEYINPUT83), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n277), .A2(G238), .A3(new_n278), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n266), .B2(new_n508), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n284), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n253), .A2(G45), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(KEYINPUT81), .A3(G250), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT81), .ZN(new_n554));
  AOI21_X1  g0354(.A(G274), .B1(new_n554), .B2(G250), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(new_n552), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT82), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n556), .A2(new_n557), .A3(new_n283), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n557), .B1(new_n556), .B2(new_n283), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n277), .A2(new_n224), .A3(G68), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n333), .A2(new_n224), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n563), .B(KEYINPUT19), .C1(new_n203), .C2(G87), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n333), .A2(G20), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n562), .B(new_n564), .C1(KEYINPUT19), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n251), .ZN(new_n567));
  INV_X1    g0367(.A(new_n367), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n319), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n450), .A2(new_n367), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n561), .A2(G179), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(G169), .B1(new_n551), .B2(new_n560), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n551), .A2(new_n560), .A3(G190), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n450), .A2(G87), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n567), .A2(new_n575), .A3(new_n569), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n422), .B1(new_n551), .B2(new_n560), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n572), .A2(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n546), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n213), .A2(G1698), .ZN(new_n581));
  OAI221_X1 g0381(.A(new_n581), .B1(G250), .B2(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G294), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n284), .A2(new_n584), .B1(new_n489), .B2(G264), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n585), .A2(new_n486), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G190), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n224), .B(G87), .C1(new_n330), .C2(new_n331), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT22), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n224), .A2(G33), .A3(G116), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n224), .A2(G107), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n591), .B(KEYINPUT23), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g0393(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n594), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n589), .A2(new_n596), .A3(new_n590), .A4(new_n592), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n251), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n450), .A2(G107), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n258), .A2(G107), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n600), .B(KEYINPUT25), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n587), .A2(new_n598), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n586), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT87), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n585), .A2(G179), .A3(new_n486), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n605), .B(new_n606), .C1(new_n586), .C2(new_n306), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n306), .B1(new_n585), .B2(new_n486), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n584), .A2(new_n284), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n489), .A2(G264), .ZN(new_n610));
  AND4_X1   g0410(.A1(G179), .A2(new_n609), .A3(new_n610), .A4(new_n486), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT87), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n602), .A2(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n505), .A2(new_n580), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n447), .A2(new_n616), .ZN(G372));
  OAI21_X1  g0417(.A(new_n614), .B1(new_n608), .B2(new_n611), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n535), .A2(new_n544), .A3(new_n545), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n619), .A2(KEYINPUT90), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(KEYINPUT90), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT89), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n561), .A2(G200), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT88), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n574), .A2(new_n576), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT88), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n578), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n561), .A2(new_n306), .ZN(new_n630));
  OAI221_X1 g0430(.A(new_n630), .B1(G179), .B2(new_n561), .C1(new_n570), .C2(new_n571), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n494), .A2(new_n504), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n602), .A2(new_n604), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n623), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n629), .A2(new_n631), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n602), .A2(new_n604), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n505), .A2(new_n635), .A3(KEYINPUT89), .A4(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n622), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n629), .A2(new_n631), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n639), .A2(KEYINPUT26), .A3(new_n494), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n494), .B2(new_n579), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n631), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n447), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n434), .A2(KEYINPUT18), .A3(new_n440), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n442), .B1(new_n432), .B2(new_n439), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n353), .A2(new_n386), .B1(new_n325), .B2(new_n359), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n430), .A2(new_n433), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n305), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n308), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n645), .A2(new_n654), .ZN(G369));
  INV_X1    g0455(.A(G13), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G20), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n253), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G343), .ZN(new_n663));
  XOR2_X1   g0463(.A(new_n663), .B(KEYINPUT91), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n523), .ZN(new_n665));
  OR3_X1    g0465(.A1(new_n620), .A2(new_n621), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n665), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n546), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  INV_X1    g0469(.A(new_n615), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n664), .A2(new_n614), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n613), .A2(new_n614), .ZN(new_n672));
  INV_X1    g0472(.A(new_n664), .ZN(new_n673));
  OAI22_X1  g0473(.A1(new_n670), .A2(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n619), .A2(new_n673), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n615), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n618), .A2(new_n664), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n681), .ZN(G399));
  NAND3_X1  g0482(.A1(new_n202), .A2(new_n210), .A3(new_n508), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT92), .ZN(new_n684));
  INV_X1    g0484(.A(new_n206), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n684), .A2(new_n253), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n230), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g0488(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n688), .B(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT26), .B1(new_n639), .B2(new_n494), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n494), .A2(new_n579), .A3(KEYINPUT26), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n631), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n619), .B1(new_n614), .B2(new_n613), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n694), .A2(new_n632), .A3(new_n633), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n673), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n664), .B1(new_n638), .B2(new_n643), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT95), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n699), .B1(new_n701), .B2(new_n698), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n505), .A2(new_n580), .A3(new_n615), .A4(new_n673), .ZN(new_n703));
  INV_X1    g0503(.A(new_n491), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n528), .A2(G179), .A3(new_n531), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n561), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n704), .A2(new_n706), .A3(KEYINPUT30), .A4(new_n585), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n561), .A2(new_n705), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n481), .A2(new_n490), .A3(new_n585), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(G179), .B1(new_n481), .B2(new_n490), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n561), .A3(new_n536), .A4(new_n603), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n707), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n714), .A2(new_n715), .A3(new_n664), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n714), .B2(new_n664), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n703), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT94), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT94), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n721), .A3(G330), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n702), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n690), .B1(new_n725), .B2(G1), .ZN(G364));
  NAND2_X1  g0526(.A1(new_n657), .A2(G45), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n727), .A2(KEYINPUT96), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(KEYINPUT96), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G1), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n686), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n669), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G330), .B2(new_n668), .ZN(new_n733));
  INV_X1    g0533(.A(new_n731), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n223), .B1(G20), .B2(new_n306), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n224), .A2(new_n437), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n422), .A2(G190), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G317), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT33), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n741), .A2(KEYINPUT33), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n224), .A2(G190), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(new_n437), .A3(new_n422), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G329), .ZN(new_n748));
  INV_X1    g0548(.A(G283), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n224), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n738), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n744), .B(new_n748), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n737), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n753), .A2(new_n298), .A3(G200), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n752), .B1(G322), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT98), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n298), .A2(new_n422), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n756), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n737), .A2(new_n757), .A3(KEYINPUT98), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G326), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n298), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n224), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G294), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n757), .A2(new_n750), .ZN(new_n767));
  INV_X1    g0567(.A(G303), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n745), .A2(G179), .A3(new_n422), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n277), .B(new_n769), .C1(G311), .C2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n755), .A2(new_n762), .A3(new_n766), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n767), .A2(new_n210), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n751), .A2(new_n498), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n774), .B(new_n775), .C1(new_n761), .C2(G50), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n770), .A2(new_n313), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n764), .A2(new_n212), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n777), .B(new_n778), .C1(G58), .C2(new_n754), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n392), .B1(new_n740), .B2(G68), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n746), .A2(new_n397), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n776), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n736), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  OR3_X1    g0584(.A1(KEYINPUT97), .A2(G13), .A3(G33), .ZN(new_n785));
  OAI21_X1  g0585(.A(KEYINPUT97), .B1(G13), .B2(G33), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n735), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n248), .A2(G45), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n685), .A2(new_n277), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(G45), .C2(new_n229), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n685), .A2(new_n392), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G355), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n793), .B(new_n795), .C1(G116), .C2(new_n206), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n734), .B(new_n784), .C1(new_n790), .C2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT99), .Z(new_n798));
  INV_X1    g0598(.A(new_n789), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n668), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n733), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  NAND2_X1  g0602(.A1(new_n664), .A2(new_n373), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n385), .A2(new_n803), .A3(new_n389), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT103), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n385), .A2(new_n803), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT103), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n385), .A2(new_n803), .A3(new_n807), .A4(new_n389), .ZN(new_n808));
  AND3_X1   g0608(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n664), .B(new_n809), .C1(new_n638), .C2(new_n643), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n701), .B2(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n813), .A2(new_n723), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n723), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n734), .A3(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n761), .A2(G303), .B1(G283), .B2(new_n740), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n508), .B2(new_n770), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT100), .Z(new_n819));
  NAND2_X1  g0619(.A1(new_n747), .A2(G311), .ZN(new_n820));
  INV_X1    g0620(.A(new_n754), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n821), .A2(new_n822), .B1(new_n751), .B2(new_n210), .ZN(new_n823));
  INV_X1    g0623(.A(new_n767), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n778), .B(new_n823), .C1(G107), .C2(new_n824), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n819), .A2(new_n392), .A3(new_n820), .A4(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT102), .B(G143), .Z(new_n827));
  AOI22_X1  g0627(.A1(new_n754), .A2(new_n827), .B1(G159), .B2(new_n771), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n761), .A2(G137), .B1(G150), .B2(new_n740), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT34), .Z(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G50), .B2(new_n824), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n834), .B1(new_n226), .B2(new_n764), .C1(new_n227), .C2(new_n751), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n277), .B1(new_n746), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n826), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n734), .B1(new_n838), .B2(new_n735), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n788), .A2(new_n736), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(G77), .B2(new_n840), .C1(new_n788), .C2(new_n812), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n816), .A2(new_n841), .ZN(G384));
  NAND2_X1  g0642(.A1(new_n664), .A2(new_n325), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n353), .A2(new_n360), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(new_n353), .B2(new_n360), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n718), .B(new_n812), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n434), .A2(new_n662), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n430), .A2(new_n433), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n648), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n412), .A2(new_n424), .A3(new_n427), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n412), .A2(new_n427), .B1(new_n439), .B2(new_n661), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT16), .B1(new_n410), .B2(new_n399), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n227), .B1(new_n408), .B2(new_n394), .ZN(new_n855));
  NOR4_X1   g0655(.A1(new_n855), .A2(new_n404), .A3(new_n398), .A4(new_n401), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n854), .A2(new_n856), .A3(new_n269), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n857), .A2(new_n426), .B1(new_n440), .B2(new_n662), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n428), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n847), .B1(new_n850), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n403), .A2(KEYINPUT104), .A3(new_n404), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n404), .A2(KEYINPUT104), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n410), .A2(new_n399), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n251), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n661), .B1(new_n866), .B2(new_n427), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n441), .A2(new_n443), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(new_n650), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n435), .A2(new_n438), .A3(new_n662), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n866), .B2(new_n427), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n851), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n860), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n862), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n846), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI221_X4 g0678(.A(new_n847), .B1(new_n872), .B2(new_n860), .C1(new_n444), .C2(new_n867), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n869), .B2(new_n873), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n877), .B1(new_n846), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT109), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT109), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n884), .B(new_n877), .C1(new_n846), .C2(new_n881), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n878), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n718), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n446), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n886), .B(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(G330), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n867), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n849), .B2(new_n648), .ZN(new_n893));
  INV_X1    g0693(.A(new_n873), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n847), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n874), .ZN(new_n896));
  INV_X1    g0696(.A(new_n843), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n361), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n353), .A2(new_n360), .A3(new_n843), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n385), .A2(new_n664), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n896), .B(new_n900), .C1(new_n810), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n868), .A2(new_n661), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT105), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT105), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT39), .B1(new_n879), .B2(new_n880), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n862), .A2(new_n909), .A3(new_n874), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(KEYINPUT107), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT107), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n862), .A2(new_n874), .A3(new_n912), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n359), .A2(new_n325), .A3(new_n673), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT106), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT108), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n919), .A3(new_n913), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n915), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n905), .A2(new_n907), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT95), .B1(new_n644), .B2(new_n673), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT95), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n924), .B(new_n664), .C1(new_n638), .C2(new_n643), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n698), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n699), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n446), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n653), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n922), .B(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT110), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n891), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(KEYINPUT110), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n932), .B1(new_n253), .B2(new_n657), .C1(new_n933), .C2(new_n891), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n457), .A2(new_n459), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n508), .B1(new_n935), .B2(KEYINPUT35), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(new_n225), .C1(KEYINPUT35), .C2(new_n935), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n400), .A2(G77), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n229), .A2(new_n939), .B1(G50), .B2(new_n227), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(G1), .A3(new_n656), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n747), .A2(G137), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n943), .B1(new_n227), .B2(new_n764), .C1(new_n397), .C2(new_n739), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n761), .A2(new_n827), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n277), .B1(new_n821), .B2(new_n260), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n767), .A2(new_n226), .ZN(new_n947));
  NOR4_X1   g0747(.A1(new_n944), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n948), .B1(new_n311), .B2(new_n770), .C1(new_n313), .C2(new_n751), .ZN(new_n949));
  INV_X1    g0749(.A(new_n761), .ZN(new_n950));
  XOR2_X1   g0750(.A(KEYINPUT111), .B(G311), .Z(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n764), .A2(new_n498), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n392), .B1(new_n746), .B2(new_n741), .C1(new_n749), .C2(new_n770), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(G303), .C2(new_n754), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n824), .A2(G116), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT46), .ZN(new_n958));
  INV_X1    g0758(.A(new_n751), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(G97), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n740), .A2(G294), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n956), .A2(new_n958), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n949), .B1(new_n953), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n735), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n673), .A2(new_n576), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n635), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n966), .A2(new_n631), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n789), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n792), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n790), .B1(new_n206), .B2(new_n568), .C1(new_n240), .C2(new_n970), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n965), .A2(new_n731), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n505), .B1(new_n502), .B2(new_n673), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n494), .A2(new_n673), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n680), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT44), .Z(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n974), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n681), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT45), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n675), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n977), .A2(new_n981), .A3(new_n675), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n678), .B1(new_n674), .B2(new_n677), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n669), .B(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n725), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n686), .B(KEYINPUT41), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n730), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n967), .A2(new_n968), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n983), .A2(new_n978), .ZN(new_n996));
  INV_X1    g0796(.A(new_n678), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n978), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT42), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n973), .A2(new_n672), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n664), .B1(new_n1000), .B2(new_n494), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n996), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n996), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n995), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n983), .A3(new_n978), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(new_n994), .A3(new_n1004), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n972), .B1(new_n992), .B2(new_n1011), .ZN(G387));
  NAND2_X1  g0812(.A1(new_n724), .A2(new_n989), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n702), .A2(new_n723), .A3(new_n988), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n686), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n674), .A2(new_n799), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n970), .B1(new_n236), .B2(G45), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n684), .B2(new_n794), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n362), .A2(new_n311), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n227), .A2(new_n313), .ZN(new_n1021));
  NOR4_X1   g0821(.A1(new_n1020), .A2(G45), .A3(new_n1021), .A4(new_n684), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1018), .A2(new_n1022), .B1(G107), .B2(new_n206), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n790), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n731), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n568), .A2(new_n764), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n265), .A2(new_n740), .B1(G150), .B2(new_n747), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n824), .A2(G77), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n311), .C2(new_n821), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1026), .B(new_n1029), .C1(G68), .C2(new_n771), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n761), .A2(G159), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1030), .A2(new_n277), .A3(new_n960), .A4(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n761), .A2(G322), .B1(G303), .B2(new_n771), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n741), .B2(new_n821), .C1(new_n739), .C2(new_n952), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT48), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n749), .B2(new_n764), .C1(new_n822), .C2(new_n767), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT49), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n959), .A2(G116), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n747), .A2(G326), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1038), .A2(new_n392), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1032), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1016), .B(new_n1025), .C1(new_n1043), .C2(new_n735), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n988), .B2(new_n730), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1015), .A2(new_n1045), .ZN(G393));
  NOR2_X1   g0846(.A1(new_n764), .A2(new_n313), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n761), .A2(G150), .B1(G159), .B2(new_n754), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(new_n362), .C2(new_n771), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n392), .B1(new_n747), .B2(new_n827), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n227), .B2(new_n767), .C1(new_n210), .C2(new_n751), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT112), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1050), .B(new_n1053), .C1(new_n311), .C2(new_n739), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT113), .Z(new_n1055));
  AOI22_X1  g0855(.A1(new_n761), .A2(G317), .B1(G311), .B2(new_n754), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT52), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n775), .B1(G294), .B2(new_n771), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n392), .C1(new_n768), .C2(new_n739), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n747), .A2(G322), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n765), .A2(G116), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n824), .A2(G283), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n736), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n790), .B1(new_n212), .B2(new_n206), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n244), .B2(new_n792), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1065), .A2(new_n734), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n799), .B2(new_n978), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n730), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n986), .B2(new_n1070), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n977), .A2(new_n675), .A3(new_n981), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n675), .B1(new_n977), .B2(new_n981), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n725), .A2(new_n1074), .A3(new_n988), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n686), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n986), .B2(new_n1014), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1071), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G390));
  AOI21_X1  g0879(.A(new_n901), .B1(new_n700), .B2(new_n812), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n844), .A2(new_n845), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n917), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n911), .A2(new_n919), .A3(new_n913), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n919), .B1(new_n911), .B2(new_n913), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n720), .A2(new_n722), .A3(new_n812), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n1081), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1081), .A2(new_n719), .A3(new_n809), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT114), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n696), .A2(new_n809), .B1(new_n385), .B2(new_n664), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n918), .B(new_n876), .C1(new_n1092), .C2(new_n900), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1085), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1085), .B2(new_n1094), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n888), .A2(G330), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n654), .B(new_n1099), .C1(new_n702), .C2(new_n446), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n720), .A2(new_n722), .A3(new_n812), .A4(new_n900), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1092), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1081), .B1(new_n719), .B2(new_n809), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1088), .B1(new_n1086), .B2(new_n1081), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n1080), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1076), .B1(new_n1098), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1085), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n915), .A2(new_n920), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1093), .B1(new_n1111), .B2(new_n1082), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1110), .B1(new_n1112), .B2(new_n1096), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n446), .A2(new_n890), .A3(new_n887), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n928), .A2(new_n653), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1106), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1109), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1098), .A2(new_n730), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n731), .B1(new_n265), .B2(new_n840), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n824), .A2(G150), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT53), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n392), .B(new_n1122), .C1(G128), .C2(new_n761), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n765), .A2(G159), .B1(new_n740), .B2(G137), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n770), .B2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT115), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G125), .B2(new_n747), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n311), .B2(new_n751), .C1(new_n836), .C2(new_n821), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT116), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n774), .A2(new_n277), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT117), .Z(new_n1133));
  AOI211_X1 g0933(.A(new_n1047), .B(new_n1133), .C1(G294), .C2(new_n747), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n950), .A2(new_n749), .B1(new_n508), .B2(new_n821), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G68), .B2(new_n959), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n212), .B2(new_n770), .C1(new_n498), .C2(new_n739), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1131), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1120), .B1(new_n1139), .B2(new_n735), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1111), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n788), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1118), .A2(new_n1119), .A3(new_n1142), .ZN(G378));
  INV_X1    g0943(.A(KEYINPUT57), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1100), .B1(new_n1098), .B2(new_n1108), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n878), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n885), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n900), .A2(new_n896), .A3(new_n718), .A4(new_n812), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n884), .B1(new_n1148), .B2(new_n877), .ZN(new_n1149));
  OAI211_X1 g0949(.A(G330), .B(new_n1146), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1151));
  NAND2_X1  g0951(.A1(new_n309), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1151), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n305), .A2(new_n308), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n270), .A2(new_n662), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1152), .A2(new_n270), .A3(new_n662), .A4(new_n1154), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1150), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n886), .B2(G330), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n922), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n906), .B1(new_n902), .B2(new_n903), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1150), .A2(new_n1159), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n886), .A2(G330), .A3(new_n1161), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n921), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1163), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1144), .B1(new_n1145), .B2(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1163), .A2(new_n1169), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1115), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(KEYINPUT57), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1171), .A2(new_n686), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n311), .B1(new_n330), .B2(G41), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n739), .A2(new_n836), .ZN(new_n1177));
  INV_X1    g0977(.A(G128), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n821), .A2(new_n1178), .B1(new_n767), .B2(new_n1125), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT119), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1177), .B(new_n1180), .C1(G137), .C2(new_n771), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n260), .B2(new_n764), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G125), .B2(new_n761), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT59), .Z(new_n1184));
  AOI21_X1  g0984(.A(G33), .B1(new_n959), .B2(G159), .ZN(new_n1185));
  INV_X1    g0985(.A(G41), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n747), .A2(G124), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT120), .Z(new_n1189));
  OAI21_X1  g0989(.A(new_n1176), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n950), .A2(new_n508), .B1(new_n227), .B2(new_n764), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT118), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT118), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(new_n392), .A3(new_n1028), .A4(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n746), .A2(new_n749), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n821), .A2(new_n498), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n751), .A2(new_n226), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n568), .A2(new_n770), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n212), .B2(new_n739), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(new_n1194), .A2(G41), .A3(new_n1195), .A4(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT58), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n735), .B1(new_n1190), .B2(new_n1202), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n731), .C1(G50), .C2(new_n840), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1161), .B2(new_n787), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1172), .B2(new_n730), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1175), .A2(new_n1206), .ZN(G375));
  NOR2_X1   g1007(.A1(new_n739), .A2(new_n1125), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n277), .B1(new_n746), .B2(new_n1178), .C1(new_n260), .C2(new_n770), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1197), .B(new_n1209), .C1(G159), .C2(new_n824), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n950), .A2(KEYINPUT123), .A3(new_n836), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT123), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n761), .B2(G132), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1210), .B1(new_n311), .B2(new_n764), .C1(new_n1211), .C2(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1208), .B(new_n1214), .C1(G137), .C2(new_n754), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n392), .B1(new_n751), .B2(new_n313), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT122), .Z(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n749), .B2(new_n821), .C1(new_n822), .C2(new_n950), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n739), .A2(new_n508), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n770), .A2(new_n498), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1026), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n212), .B2(new_n767), .C1(new_n768), .C2(new_n746), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n735), .B1(new_n1215), .B2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n731), .C1(G68), .C2(new_n840), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1081), .B2(new_n787), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n730), .B(KEYINPUT121), .Z(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1106), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n991), .B1(new_n1115), .B2(new_n1106), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1229), .B2(new_n1108), .ZN(G381));
  NOR2_X1   g1030(.A1(G375), .A2(G378), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1078), .B(new_n972), .C1(new_n992), .C2(new_n1011), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1015), .A2(new_n801), .A3(new_n1045), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1232), .A2(G384), .A3(G381), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(G407));
  INV_X1    g1035(.A(G343), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1231), .B1(new_n1236), .B2(new_n1234), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(G213), .ZN(G409));
  NAND2_X1  g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1233), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1232), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n724), .B1(new_n1074), .B2(new_n988), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n991), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1070), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1005), .A2(new_n1006), .A3(new_n995), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n994), .B1(new_n1009), .B2(new_n1004), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1078), .B1(new_n1249), .B2(new_n972), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1241), .B1(new_n1242), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n1232), .A3(new_n1240), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT125), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1255), .B(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(G213), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1258), .A2(G343), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1175), .A2(G378), .A3(new_n1206), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1119), .A2(new_n1142), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1117), .B2(new_n1109), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1227), .B1(new_n1173), .B2(new_n991), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(new_n1170), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1264), .B2(new_n1205), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1259), .B1(new_n1260), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1115), .B2(new_n1106), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n1107), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n686), .A4(new_n1116), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1270), .A2(G384), .A3(new_n1228), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G384), .B1(new_n1270), .B2(new_n1228), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1259), .A2(G2897), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT124), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1270), .A2(new_n1228), .ZN(new_n1278));
  INV_X1    g1078(.A(G384), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1270), .A2(G384), .A3(new_n1228), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(KEYINPUT124), .A3(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1277), .A2(new_n1282), .A3(new_n1274), .ZN(new_n1283));
  OR3_X1    g1083(.A1(new_n1266), .A2(new_n1275), .A3(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1277), .A2(new_n1282), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1266), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1285), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1257), .A2(new_n1284), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1260), .A2(new_n1265), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1259), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1285), .A4(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1252), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1266), .A2(new_n1275), .A3(new_n1283), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1292), .B1(new_n1266), .B2(new_n1285), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1251), .A2(KEYINPUT126), .A3(new_n1254), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT126), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1300));
  OR2_X1    g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1290), .B1(new_n1298), .B2(new_n1301), .ZN(G405));
  NAND2_X1  g1102(.A1(G375), .A2(new_n1262), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1260), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1285), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G375), .A2(KEYINPUT127), .A3(new_n1262), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1273), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1308), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1260), .A2(new_n1304), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G378), .B1(new_n1175), .B2(new_n1206), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1307), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1273), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1301), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1312), .A2(new_n1319), .ZN(G402));
endmodule


