

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XOR2_X1 U325 ( .A(n394), .B(n393), .Z(n467) );
  XNOR2_X1 U326 ( .A(KEYINPUT122), .B(KEYINPUT55), .ZN(n436) );
  NOR2_X1 U327 ( .A1(n523), .A2(n463), .ZN(n460) );
  XNOR2_X1 U328 ( .A(n303), .B(n352), .ZN(n304) );
  XNOR2_X1 U329 ( .A(n305), .B(n304), .ZN(n309) );
  XNOR2_X1 U330 ( .A(KEYINPUT107), .B(KEYINPUT37), .ZN(n495) );
  XNOR2_X1 U331 ( .A(n437), .B(n436), .ZN(n455) );
  XNOR2_X1 U332 ( .A(n496), .B(n495), .ZN(n522) );
  XOR2_X1 U333 ( .A(n454), .B(n453), .Z(n536) );
  INV_X1 U334 ( .A(KEYINPUT40), .ZN(n504) );
  XNOR2_X1 U335 ( .A(n456), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U336 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U337 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XNOR2_X1 U338 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n310) );
  XOR2_X1 U339 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n294) );
  NAND2_X1 U340 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U342 ( .A(n295), .B(KEYINPUT75), .Z(n301) );
  XNOR2_X1 U343 ( .A(G176GAT), .B(G204GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(G64GAT), .B(G92GAT), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n377) );
  INV_X1 U346 ( .A(n377), .ZN(n376) );
  XOR2_X1 U347 ( .A(G78GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n425) );
  XNOR2_X1 U350 ( .A(n376), .B(n425), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U352 ( .A(G120GAT), .B(G71GAT), .Z(n438) );
  XOR2_X1 U353 ( .A(G99GAT), .B(G85GAT), .Z(n331) );
  XOR2_X1 U354 ( .A(n438), .B(n331), .Z(n303) );
  XNOR2_X1 U355 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n302), .B(KEYINPUT13), .ZN(n352) );
  XOR2_X1 U357 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n307) );
  XNOR2_X1 U358 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n580) );
  XNOR2_X1 U361 ( .A(n310), .B(n580), .ZN(n555) );
  XOR2_X1 U362 ( .A(G113GAT), .B(G197GAT), .Z(n312) );
  XNOR2_X1 U363 ( .A(G141GAT), .B(G22GAT), .ZN(n311) );
  XOR2_X1 U364 ( .A(n312), .B(n311), .Z(n327) );
  XOR2_X1 U365 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U368 ( .A(G36GAT), .B(G50GAT), .Z(n316) );
  XOR2_X1 U369 ( .A(G169GAT), .B(G8GAT), .Z(n387) );
  XOR2_X1 U370 ( .A(G15GAT), .B(G1GAT), .Z(n349) );
  XNOR2_X1 U371 ( .A(n387), .B(n349), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U373 ( .A(n318), .B(n317), .Z(n320) );
  NAND2_X1 U374 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U376 ( .A(n321), .B(KEYINPUT68), .Z(n325) );
  XOR2_X1 U377 ( .A(G29GAT), .B(G43GAT), .Z(n323) );
  XNOR2_X1 U378 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n334) );
  XNOR2_X1 U380 ( .A(n334), .B(KEYINPUT69), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n537) );
  NAND2_X1 U383 ( .A1(n555), .A2(n537), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n328), .B(KEYINPUT46), .ZN(n366) );
  XOR2_X1 U385 ( .A(KEYINPUT78), .B(KEYINPUT10), .Z(n330) );
  XNOR2_X1 U386 ( .A(KEYINPUT11), .B(KEYINPUT66), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n345) );
  XOR2_X1 U388 ( .A(G36GAT), .B(G190GAT), .Z(n382) );
  XOR2_X1 U389 ( .A(n331), .B(n382), .Z(n333) );
  XNOR2_X1 U390 ( .A(G218GAT), .B(G106GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U392 ( .A(G134GAT), .B(n334), .Z(n336) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U395 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U396 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XOR2_X1 U397 ( .A(KEYINPUT9), .B(KEYINPUT79), .Z(n340) );
  XNOR2_X1 U398 ( .A(G92GAT), .B(KEYINPUT80), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n422), .B(n341), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n548) );
  INV_X1 U403 ( .A(n548), .ZN(n561) );
  XOR2_X1 U404 ( .A(G78GAT), .B(G211GAT), .Z(n347) );
  XNOR2_X1 U405 ( .A(G183GAT), .B(G127GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U407 ( .A(n348), .B(G71GAT), .Z(n351) );
  XNOR2_X1 U408 ( .A(G8GAT), .B(n349), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n356) );
  XOR2_X1 U410 ( .A(G22GAT), .B(G155GAT), .Z(n423) );
  XOR2_X1 U411 ( .A(n352), .B(n423), .Z(n354) );
  NAND2_X1 U412 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U414 ( .A(n356), .B(n355), .Z(n364) );
  XOR2_X1 U415 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n358) );
  XNOR2_X1 U416 ( .A(G64GAT), .B(KEYINPUT83), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n360) );
  XNOR2_X1 U419 ( .A(KEYINPUT81), .B(KEYINPUT15), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U422 ( .A(n364), .B(n363), .Z(n543) );
  INV_X1 U423 ( .A(n543), .ZN(n584) );
  AND2_X1 U424 ( .A1(n561), .A2(n584), .ZN(n365) );
  AND2_X1 U425 ( .A1(n366), .A2(n365), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n367), .B(KEYINPUT47), .ZN(n373) );
  XOR2_X1 U427 ( .A(KEYINPUT36), .B(n548), .Z(n587) );
  NOR2_X1 U428 ( .A1(n584), .A2(n587), .ZN(n369) );
  XNOR2_X1 U429 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n371) );
  INV_X1 U431 ( .A(n537), .ZN(n575) );
  AND2_X1 U432 ( .A1(n575), .A2(n580), .ZN(n370) );
  NAND2_X1 U433 ( .A1(n371), .A2(n370), .ZN(n372) );
  NAND2_X1 U434 ( .A1(n373), .A2(n372), .ZN(n374) );
  XNOR2_X1 U435 ( .A(KEYINPUT48), .B(n374), .ZN(n531) );
  INV_X1 U436 ( .A(KEYINPUT97), .ZN(n375) );
  NAND2_X1 U437 ( .A1(n376), .A2(n375), .ZN(n379) );
  NAND2_X1 U438 ( .A1(KEYINPUT97), .A2(n377), .ZN(n378) );
  NAND2_X1 U439 ( .A1(n379), .A2(n378), .ZN(n381) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n383) );
  XOR2_X1 U442 ( .A(n383), .B(n382), .Z(n389) );
  XOR2_X1 U443 ( .A(KEYINPUT92), .B(G218GAT), .Z(n385) );
  XNOR2_X1 U444 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(G197GAT), .B(n386), .Z(n433) );
  XNOR2_X1 U447 ( .A(n387), .B(n433), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n394) );
  XOR2_X1 U449 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n391) );
  XNOR2_X1 U450 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U452 ( .A(KEYINPUT18), .B(n392), .ZN(n452) );
  INV_X1 U453 ( .A(n452), .ZN(n393) );
  NAND2_X1 U454 ( .A1(n531), .A2(n467), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n395), .B(KEYINPUT54), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n396), .B(KEYINPUT121), .ZN(n419) );
  XOR2_X1 U457 ( .A(G57GAT), .B(G155GAT), .Z(n398) );
  XNOR2_X1 U458 ( .A(G1GAT), .B(G120GAT), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U460 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n400) );
  XNOR2_X1 U461 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U463 ( .A(n402), .B(n401), .Z(n407) );
  XOR2_X1 U464 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n404) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U467 ( .A(KEYINPUT4), .B(n405), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n412) );
  XNOR2_X1 U469 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n408), .B(KEYINPUT2), .ZN(n421) );
  XOR2_X1 U471 ( .A(G85GAT), .B(n421), .Z(n410) );
  XNOR2_X1 U472 ( .A(G148GAT), .B(G162GAT), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U474 ( .A(n412), .B(n411), .Z(n418) );
  INV_X1 U475 ( .A(G113GAT), .ZN(n416) );
  XOR2_X1 U476 ( .A(KEYINPUT86), .B(G134GAT), .Z(n414) );
  XNOR2_X1 U477 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n442) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(n442), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n523) );
  NAND2_X1 U482 ( .A1(n419), .A2(n523), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n420), .B(KEYINPUT65), .ZN(n574) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n429) );
  XOR2_X1 U486 ( .A(n425), .B(KEYINPUT22), .Z(n427) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U489 ( .A(n429), .B(n428), .Z(n435) );
  XOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n431) );
  XNOR2_X1 U491 ( .A(KEYINPUT93), .B(G204GAT), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n470) );
  NAND2_X1 U495 ( .A1(n574), .A2(n470), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(KEYINPUT91), .ZN(n440) );
  AND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U499 ( .A(n441), .B(G99GAT), .Z(n444) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U502 ( .A(KEYINPUT90), .B(G176GAT), .Z(n446) );
  XNOR2_X1 U503 ( .A(G15GAT), .B(G190GAT), .ZN(n445) );
  XOR2_X1 U504 ( .A(n446), .B(n445), .Z(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n450) );
  XNOR2_X1 U507 ( .A(G169GAT), .B(KEYINPUT89), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U509 ( .A(n452), .B(n451), .Z(n453) );
  INV_X1 U510 ( .A(n536), .ZN(n468) );
  NAND2_X1 U511 ( .A1(n455), .A2(n468), .ZN(n570) );
  NOR2_X1 U512 ( .A1(n570), .A2(n561), .ZN(n458) );
  INV_X1 U513 ( .A(G190GAT), .ZN(n456) );
  INV_X1 U514 ( .A(n467), .ZN(n485) );
  XOR2_X1 U515 ( .A(n485), .B(KEYINPUT98), .Z(n459) );
  XOR2_X1 U516 ( .A(n459), .B(KEYINPUT27), .Z(n463) );
  XOR2_X1 U517 ( .A(KEYINPUT99), .B(n460), .Z(n532) );
  XOR2_X1 U518 ( .A(n470), .B(KEYINPUT67), .Z(n461) );
  XNOR2_X1 U519 ( .A(KEYINPUT28), .B(n461), .ZN(n534) );
  AND2_X1 U520 ( .A1(n534), .A2(n536), .ZN(n462) );
  AND2_X1 U521 ( .A1(n532), .A2(n462), .ZN(n477) );
  INV_X1 U522 ( .A(n463), .ZN(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n468), .A2(n470), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n465), .B(n464), .ZN(n573) );
  NAND2_X1 U526 ( .A1(n466), .A2(n573), .ZN(n473) );
  NAND2_X1 U527 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n471) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n471), .Z(n472) );
  NAND2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n474), .A2(n523), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n475), .B(KEYINPUT101), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n477), .A2(n476), .ZN(n494) );
  NOR2_X1 U534 ( .A1(n584), .A2(n548), .ZN(n479) );
  XNOR2_X1 U535 ( .A(KEYINPUT16), .B(KEYINPUT85), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n494), .A2(n480), .ZN(n481) );
  XOR2_X1 U538 ( .A(KEYINPUT102), .B(n481), .Z(n509) );
  NAND2_X1 U539 ( .A1(n537), .A2(n580), .ZN(n497) );
  NOR2_X1 U540 ( .A1(n509), .A2(n497), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT103), .ZN(n490) );
  NOR2_X1 U542 ( .A1(n523), .A2(n490), .ZN(n483) );
  XOR2_X1 U543 ( .A(KEYINPUT34), .B(n483), .Z(n484) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U545 ( .A1(n485), .A2(n490), .ZN(n486) );
  XOR2_X1 U546 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  NOR2_X1 U547 ( .A1(n536), .A2(n490), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT35), .B(KEYINPUT104), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n489), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n534), .A2(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1327GAT) );
  OR2_X1 U554 ( .A1(n543), .A2(n587), .ZN(n493) );
  OR2_X1 U555 ( .A1(n494), .A2(n493), .ZN(n496) );
  NOR2_X1 U556 ( .A1(n497), .A2(n522), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT38), .B(n498), .Z(n499) );
  XNOR2_X1 U558 ( .A(KEYINPUT108), .B(n499), .ZN(n507) );
  NOR2_X1 U559 ( .A1(n523), .A2(n507), .ZN(n501) );
  XNOR2_X1 U560 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n485), .A2(n507), .ZN(n503) );
  XOR2_X1 U564 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  NOR2_X1 U565 ( .A1(n507), .A2(n536), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NOR2_X1 U567 ( .A1(n534), .A2(n507), .ZN(n508) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  NAND2_X1 U569 ( .A1(n575), .A2(n555), .ZN(n521) );
  NOR2_X1 U570 ( .A1(n521), .A2(n509), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n510), .B(KEYINPUT109), .ZN(n518) );
  NOR2_X1 U572 ( .A1(n523), .A2(n518), .ZN(n511) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n485), .A2(n518), .ZN(n513) );
  XOR2_X1 U576 ( .A(KEYINPUT110), .B(n513), .Z(n514) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n536), .A2(n518), .ZN(n516) );
  XNOR2_X1 U579 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(n517), .ZN(G1334GAT) );
  NOR2_X1 U582 ( .A1(n534), .A2(n518), .ZN(n520) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  OR2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U586 ( .A1(n523), .A2(n528), .ZN(n524) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n524), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n485), .A2(n528), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1337GAT) );
  NOR2_X1 U591 ( .A1(n536), .A2(n528), .ZN(n527) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n534), .A2(n528), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n529), .Z(n530) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(KEYINPUT115), .ZN(n552) );
  NAND2_X1 U598 ( .A1(n552), .A2(n534), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n549) );
  NAND2_X1 U600 ( .A1(n537), .A2(n549), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n540) );
  NAND2_X1 U603 ( .A1(n549), .A2(n555), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT116), .Z(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n543), .A2(n549), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n545) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n573), .A2(n552), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n575), .A2(n560), .ZN(n553) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n553), .Z(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT120), .B(n554), .ZN(G1344GAT) );
  INV_X1 U619 ( .A(n555), .ZN(n567) );
  NOR2_X1 U620 ( .A1(n567), .A2(n560), .ZN(n557) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n584), .A2(n560), .ZN(n559) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NOR2_X1 U628 ( .A1(n570), .A2(n575), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT123), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n566) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n567), .A2(n570), .ZN(n568) );
  XOR2_X1 U635 ( .A(n569), .B(n568), .Z(G1349GAT) );
  NOR2_X1 U636 ( .A1(n584), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1350GAT) );
  XNOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT59), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n586) );
  NOR2_X1 U641 ( .A1(n575), .A2(n586), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n586), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n586), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

