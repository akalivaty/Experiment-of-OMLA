//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT27), .Z(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n191), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT69), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT2), .B(G113), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n200), .A2(new_n204), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT66), .A2(G137), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT66), .A2(G137), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .A4(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT11), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n215), .A2(new_n217), .B1(new_n218), .B2(G137), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(G137), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n210), .B(new_n213), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n220), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n218), .A2(G137), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n227), .A2(KEYINPUT67), .A3(new_n210), .A4(new_n213), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n211), .A2(new_n212), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n218), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n210), .B1(new_n231), .B2(new_n224), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  INV_X1    g049(.A(G143), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT64), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n233), .A2(G143), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(KEYINPUT1), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n242), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT64), .B(G143), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G146), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n232), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n229), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n210), .B1(new_n227), .B2(new_n213), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n229), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n240), .A2(new_n259), .B1(new_n248), .B2(new_n257), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n253), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n254), .B1(new_n223), .B2(new_n228), .ZN(new_n262));
  INV_X1    g076(.A(new_n260), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n262), .A2(KEYINPUT70), .A3(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n209), .B(new_n252), .C1(new_n261), .C2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n252), .B1(new_n262), .B2(new_n263), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n208), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n195), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n195), .B1(new_n266), .B2(new_n208), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n194), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT73), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n243), .B1(new_n238), .B2(new_n239), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n236), .A2(KEYINPUT64), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n234), .A2(G143), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G146), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n277), .A2(new_n242), .A3(new_n249), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n220), .B1(new_n230), .B2(new_n218), .ZN(new_n279));
  OAI22_X1  g093(.A1(new_n274), .A2(new_n278), .B1(new_n210), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n223), .B2(new_n228), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n256), .A2(new_n253), .A3(new_n260), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT70), .B1(new_n262), .B2(new_n263), .ZN(new_n283));
  AOI211_X1 g097(.A(new_n208), .B(new_n281), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n273), .B1(new_n284), .B2(new_n194), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n265), .A2(KEYINPUT72), .A3(new_n193), .ZN(new_n286));
  OAI211_X1 g100(.A(KEYINPUT30), .B(new_n252), .C1(new_n261), .C2(new_n264), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n263), .B1(new_n229), .B2(new_n255), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(new_n281), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n288), .B1(new_n266), .B2(new_n289), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n287), .B(new_n208), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n289), .B1(new_n290), .B2(new_n281), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT68), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n291), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(KEYINPUT71), .A3(new_n208), .A4(new_n287), .ZN(new_n300));
  AOI221_X4 g114(.A(KEYINPUT31), .B1(new_n285), .B2(new_n286), .C1(new_n296), .C2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT31), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n300), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n285), .A2(new_n286), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n272), .A2(new_n301), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n187), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n303), .A2(new_n304), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT31), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n271), .B(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n303), .A2(new_n302), .A3(new_n304), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT32), .A3(new_n307), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n252), .B1(new_n261), .B2(new_n264), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n208), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n265), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT28), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n269), .A2(new_n193), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(G902), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n193), .B1(new_n303), .B2(new_n265), .ZN(new_n325));
  INV_X1    g139(.A(new_n321), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n265), .A2(new_n267), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(KEYINPUT74), .C1(new_n327), .C2(new_n195), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n268), .B2(new_n321), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n322), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n324), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT75), .B1(new_n332), .B2(G472), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n334));
  INV_X1    g148(.A(G472), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n268), .A2(new_n321), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT29), .B1(new_n336), .B2(KEYINPUT74), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n284), .B1(new_n296), .B2(new_n300), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n337), .B(new_n330), .C1(new_n338), .C2(new_n193), .ZN(new_n339));
  AOI211_X1 g153(.A(new_n334), .B(new_n335), .C1(new_n339), .C2(new_n324), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n309), .B(new_n316), .C1(new_n333), .C2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G217), .ZN(new_n342));
  INV_X1    g156(.A(G902), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(G234), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT76), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G137), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G125), .B(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT16), .ZN(new_n350));
  INV_X1    g164(.A(G125), .ZN(new_n351));
  OR3_X1    g165(.A1(new_n351), .A2(KEYINPUT16), .A3(G140), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(G146), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n350), .A2(KEYINPUT80), .A3(G146), .A4(new_n352), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n233), .B2(new_n349), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n241), .A2(KEYINPUT23), .A3(G119), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G110), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n196), .A2(G128), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT78), .B1(new_n363), .B2(KEYINPUT23), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n241), .A2(G119), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n361), .B(new_n362), .C1(new_n364), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT79), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n367), .A2(new_n364), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n362), .A4(new_n361), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n363), .A2(new_n366), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT24), .B(G110), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n369), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n358), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n370), .A2(new_n361), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G110), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n373), .A2(new_n374), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n350), .A2(new_n352), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n233), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n381), .B1(new_n383), .B2(new_n353), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n377), .A2(new_n378), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n378), .B1(new_n377), .B2(new_n385), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n348), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n348), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n377), .A2(new_n385), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(KEYINPUT81), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT25), .ZN(new_n393));
  AOI21_X1  g207(.A(G902), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n392), .A2(new_n393), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n345), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n396), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n388), .A2(new_n398), .A3(new_n391), .A4(new_n394), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n388), .A2(new_n391), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n344), .A2(G902), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G469), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G140), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n189), .A2(G227), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT10), .ZN(new_n411));
  INV_X1    g225(.A(new_n248), .ZN(new_n412));
  AOI21_X1  g226(.A(G146), .B1(new_n275), .B2(new_n276), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT1), .ZN(new_n414));
  OAI21_X1  g228(.A(G128), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n278), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n417));
  INV_X1    g231(.A(G104), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT3), .B1(new_n418), .B2(G107), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT3), .ZN(new_n420));
  INV_X1    g234(.A(G107), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n421), .A3(G104), .ZN(new_n422));
  INV_X1    g236(.A(G101), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n418), .A2(G107), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n419), .A2(new_n422), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n418), .A2(G107), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n421), .A2(G104), .ZN(new_n427));
  OAI21_X1  g241(.A(G101), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n416), .A2(new_n417), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n241), .B1(new_n238), .B2(KEYINPUT1), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n250), .B1(new_n431), .B2(new_n248), .ZN(new_n432));
  INV_X1    g246(.A(new_n429), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT85), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n411), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT86), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n417), .B1(new_n416), .B2(new_n429), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(KEYINPUT85), .A3(new_n433), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n411), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n245), .A2(new_n250), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT10), .A3(new_n433), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT4), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(G101), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(G101), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT4), .A3(new_n425), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n260), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n262), .B1(new_n442), .B2(new_n452), .ZN(new_n453));
  AOI211_X1 g267(.A(new_n256), .B(new_n451), .C1(new_n436), .C2(new_n441), .ZN(new_n454));
  OAI211_X1 g268(.A(KEYINPUT87), .B(new_n410), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n440), .B1(new_n439), .B2(new_n411), .ZN(new_n456));
  AOI211_X1 g270(.A(KEYINPUT86), .B(KEYINPUT10), .C1(new_n437), .C2(new_n438), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n262), .B(new_n452), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n410), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n443), .A2(new_n433), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(new_n437), .B2(new_n438), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT12), .ZN(new_n463));
  OR3_X1    g277(.A1(new_n462), .A2(new_n463), .A3(new_n262), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n463), .B1(new_n462), .B2(new_n262), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n455), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n256), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n458), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT87), .B1(new_n471), .B2(new_n410), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n407), .B(new_n343), .C1(new_n468), .C2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n407), .A2(new_n343), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n459), .B1(new_n466), .B2(new_n458), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n470), .B2(new_n460), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n476), .B2(G469), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT9), .B(G234), .ZN(new_n479));
  OAI21_X1  g293(.A(G221), .B1(new_n479), .B2(G902), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT83), .Z(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT84), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G122), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G116), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n198), .B2(G122), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(KEYINPUT14), .B2(new_n421), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n485), .B(KEYINPUT96), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(G116), .B2(new_n484), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(KEYINPUT14), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(G107), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n236), .A2(G128), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n247), .B2(G128), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(new_n218), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n218), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n489), .B(new_n493), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(KEYINPUT97), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n247), .A2(G128), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n501), .B(G134), .C1(new_n502), .C2(new_n500), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n488), .A2(new_n421), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n491), .A2(G107), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n503), .B(new_n497), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n479), .A2(new_n342), .A3(G953), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n499), .A2(new_n506), .A3(new_n508), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT98), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n515), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n189), .A2(G952), .ZN(new_n518));
  INV_X1    g332(.A(G234), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n518), .B1(new_n519), .B2(new_n188), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n343), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n516), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n418), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n349), .B(KEYINPUT19), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n357), .B1(new_n233), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n531));
  MUX2_X1   g345(.A(G143), .B(new_n247), .S(new_n531), .Z(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G131), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n532), .A2(G131), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT95), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n532), .A2(G131), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n533), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n349), .B(new_n233), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n210), .ZN(new_n543));
  OAI221_X1 g357(.A(new_n541), .B1(new_n532), .B2(new_n543), .C1(new_n533), .C2(new_n542), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n528), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT17), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n383), .B(new_n353), .C1(new_n533), .C2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n528), .B(new_n544), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT20), .ZN(new_n552));
  NOR2_X1   g366(.A1(G475), .A2(G902), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n545), .A2(new_n550), .ZN(new_n555));
  INV_X1    g369(.A(new_n553), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT20), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n544), .B1(new_n546), .B2(new_n548), .ZN(new_n559));
  INV_X1    g373(.A(new_n528), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n343), .B1(new_n561), .B2(new_n550), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G475), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n526), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G214), .B1(G237), .B2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n202), .A2(new_n203), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT5), .ZN(new_n568));
  OAI21_X1  g382(.A(G113), .B1(new_n197), .B2(KEYINPUT5), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n207), .A4(new_n433), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT5), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n202), .B2(new_n203), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n433), .B(new_n207), .C1(new_n575), .C2(new_n569), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT89), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n208), .A2(new_n447), .A3(new_n449), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT88), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n208), .A2(KEYINPUT88), .A3(new_n449), .A4(new_n447), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G122), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n578), .A2(new_n583), .A3(new_n585), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(KEYINPUT6), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT6), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n584), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n263), .A2(G125), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n245), .A2(new_n351), .A3(new_n250), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT90), .B(G224), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n189), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT91), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n594), .B(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n589), .A2(new_n591), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n593), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n260), .A2(new_n351), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT7), .ZN(new_n602));
  OAI22_X1  g416(.A1(new_n600), .A2(new_n601), .B1(new_n602), .B2(new_n597), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n597), .A2(new_n602), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n592), .A2(new_n604), .A3(new_n593), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n206), .B1(new_n568), .B2(new_n570), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n608));
  OR3_X1    g422(.A1(new_n607), .A2(new_n608), .A3(new_n433), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n200), .A2(new_n574), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n207), .B1(new_n610), .B2(new_n569), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n429), .B1(new_n611), .B2(KEYINPUT93), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n612), .B1(KEYINPUT93), .B2(new_n611), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n608), .B1(new_n607), .B2(new_n433), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n609), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT92), .B(KEYINPUT8), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(new_n585), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n606), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n618), .B2(new_n588), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n599), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G210), .B1(G237), .B2(G902), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n599), .A2(new_n621), .A3(new_n619), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n565), .A2(new_n566), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n483), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n341), .A2(new_n406), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  OAI21_X1  g443(.A(G472), .B1(new_n306), .B2(G902), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n315), .A2(new_n307), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n632), .A2(new_n405), .A3(new_n483), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n625), .B2(new_n566), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n599), .A2(new_n621), .A3(new_n619), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n621), .B1(new_n599), .B2(new_n619), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n634), .B(new_n566), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n510), .A2(new_n511), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT33), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n510), .A2(new_n643), .A3(new_n511), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n642), .A2(G478), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n514), .A2(new_n343), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n512), .B2(new_n514), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n645), .A2(new_n647), .A3(KEYINPUT100), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT100), .B1(new_n645), .B2(new_n647), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n564), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n640), .A2(new_n524), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n633), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  INV_X1    g469(.A(new_n564), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n516), .A2(new_n517), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n640), .A2(new_n524), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n633), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n389), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT101), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n390), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n403), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n397), .B2(new_n399), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT102), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n627), .A2(new_n631), .A3(new_n630), .A4(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  NOR2_X1   g487(.A1(new_n483), .A2(new_n669), .ZN(new_n674));
  INV_X1    g488(.A(G900), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n522), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n520), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n566), .B1(new_n636), .B2(new_n637), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT99), .ZN(new_n680));
  AOI211_X1 g494(.A(new_n678), .B(new_n658), .C1(new_n680), .C2(new_n638), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n309), .A2(new_n316), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n340), .A2(new_n333), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n674), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XNOR2_X1  g499(.A(new_n625), .B(KEYINPUT38), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n564), .A2(new_n657), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n686), .A2(new_n566), .A3(new_n668), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n677), .B(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n478), .A2(new_n482), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n689), .B1(new_n692), .B2(KEYINPUT40), .ZN(new_n693));
  INV_X1    g507(.A(new_n310), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n194), .B2(new_n319), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n309), .A2(new_n696), .A3(new_n316), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n693), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n693), .A2(KEYINPUT104), .A3(new_n697), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n247), .ZN(G45));
  OAI211_X1 g518(.A(new_n564), .B(new_n677), .C1(new_n648), .C2(new_n649), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n640), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n674), .B(new_n706), .C1(new_n682), .C2(new_n683), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  OAI21_X1  g522(.A(new_n343), .B1(new_n468), .B2(new_n472), .ZN(new_n709));
  NAND2_X1  g523(.A1(KEYINPUT105), .A2(G469), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n481), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n343), .B(new_n710), .C1(new_n468), .C2(new_n472), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n341), .A2(new_n716), .A3(new_n652), .A4(new_n406), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n341), .A2(new_n716), .A3(new_n659), .A4(new_n406), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NOR2_X1   g535(.A1(new_n715), .A2(new_n640), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n341), .A2(new_n565), .A3(new_n670), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  AOI21_X1  g538(.A(new_n335), .B1(new_n315), .B2(new_n343), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n301), .A2(new_n305), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n320), .A2(new_n269), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n194), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n308), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n725), .A2(new_n729), .A3(new_n405), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n712), .A2(new_n713), .A3(new_n525), .A4(new_n714), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n688), .B1(new_n635), .B2(new_n639), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n730), .A2(new_n733), .A3(KEYINPUT106), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT106), .B1(new_n730), .B2(new_n733), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NOR3_X1   g551(.A1(new_n725), .A2(new_n729), .A3(new_n668), .ZN(new_n738));
  INV_X1    g552(.A(new_n705), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n722), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  AOI21_X1  g555(.A(new_n335), .B1(new_n339), .B2(new_n324), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT75), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n315), .A2(KEYINPUT32), .A3(new_n307), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT110), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n316), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n743), .A2(new_n745), .A3(new_n309), .A4(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT107), .B1(new_n478), .B2(new_n713), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n750));
  AOI211_X1 g564(.A(new_n750), .B(new_n481), .C1(new_n473), .C2(new_n477), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n636), .A2(new_n637), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n566), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n739), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n749), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n748), .A2(KEYINPUT42), .A3(new_n406), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n756), .A2(new_n758), .A3(new_n341), .A4(new_n406), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT32), .B1(new_n315), .B2(new_n307), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n744), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n405), .B1(new_n763), .B2(new_n743), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n758), .B1(new_n764), .B2(new_n756), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n757), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NOR2_X1   g581(.A1(new_n749), .A2(new_n751), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n658), .A2(new_n753), .A3(new_n678), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n341), .A2(new_n768), .A3(new_n406), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  NAND2_X1  g585(.A1(new_n650), .A2(new_n656), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n650), .B(new_n656), .C1(KEYINPUT111), .C2(KEYINPUT43), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n668), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n632), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(new_n632), .A3(KEYINPUT44), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(KEYINPUT112), .A3(new_n754), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n476), .A2(KEYINPUT45), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n453), .A2(new_n454), .A3(new_n410), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n783), .B1(new_n784), .B2(new_n475), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n785), .A3(G469), .ZN(new_n786));
  INV_X1    g600(.A(new_n474), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT46), .ZN(new_n789));
  INV_X1    g603(.A(new_n473), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n786), .A2(new_n787), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n481), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n794), .A2(new_n691), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n781), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n779), .A2(new_n754), .A3(new_n780), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(KEYINPUT113), .B(G137), .Z(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(G39));
  NAND2_X1  g616(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n794), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g618(.A(KEYINPUT114), .B(KEYINPUT47), .Z(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n341), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n755), .A2(new_n406), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  AND2_X1   g625(.A1(new_n684), .A2(new_n740), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  INV_X1    g627(.A(new_n732), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n481), .B1(new_n473), .B2(new_n477), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n668), .A2(new_n677), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n815), .A2(KEYINPUT115), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT115), .B1(new_n815), .B2(new_n816), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n697), .B(new_n814), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n812), .A2(new_n813), .A3(new_n707), .A4(new_n819), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n753), .A2(new_n564), .A3(new_n657), .A4(new_n678), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n341), .A2(new_n674), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n755), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n768), .A2(new_n738), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n770), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n679), .B(new_n524), .C1(new_n651), .C2(new_n658), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n483), .A2(new_n405), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n631), .A4(new_n630), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n628), .A2(new_n671), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n819), .A2(new_n684), .A3(new_n707), .A4(new_n740), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT52), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n820), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n720), .B1(new_n734), .B2(new_n735), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n717), .A2(new_n723), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n766), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT53), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n766), .A2(new_n837), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n684), .A2(new_n740), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n841), .B2(KEYINPUT52), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n833), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n841), .B2(KEYINPUT52), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n820), .A2(new_n830), .A3(new_n832), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n766), .A2(new_n837), .A3(KEYINPUT116), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n847), .B1(new_n833), .B2(new_n840), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n844), .B1(KEYINPUT54), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n855));
  INV_X1    g669(.A(new_n697), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n715), .A2(new_n405), .A3(new_n520), .A4(new_n753), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n858), .A2(new_n564), .A3(new_n650), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n520), .B1(new_n774), .B2(new_n775), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n730), .A2(new_n860), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n715), .A2(new_n686), .A3(new_n566), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT50), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n860), .A2(new_n716), .A3(new_n754), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n738), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT50), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n859), .A2(new_n865), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n712), .A2(new_n714), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n806), .B1(new_n482), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n730), .A2(new_n860), .A3(new_n754), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(KEYINPUT118), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n855), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n748), .A2(new_n406), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n866), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT48), .Z(new_n883));
  NAND3_X1  g697(.A1(new_n730), .A2(new_n860), .A3(new_n722), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n518), .B(new_n884), .C1(new_n858), .C2(new_n651), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n878), .A2(new_n879), .A3(new_n886), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n854), .A2(new_n887), .B1(G952), .B2(G953), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n482), .A2(new_n566), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n772), .A2(new_n405), .A3(new_n889), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n686), .B(new_n890), .C1(KEYINPUT49), .C2(new_n870), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(new_n856), .C1(KEYINPUT49), .C2(new_n870), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n888), .A2(new_n892), .ZN(G75));
  NAND3_X1  g707(.A1(new_n853), .A2(G210), .A3(G902), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n589), .A2(new_n591), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n598), .ZN(new_n897));
  XOR2_X1   g711(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n894), .B2(new_n895), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n189), .A2(G952), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G51));
  XNOR2_X1  g717(.A(new_n474), .B(KEYINPUT57), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n851), .A2(new_n905), .A3(new_n852), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n851), .B2(new_n852), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n468), .A2(new_n472), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n343), .B1(new_n851), .B2(new_n852), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(G469), .A3(new_n782), .A4(new_n785), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n902), .B1(new_n910), .B2(new_n912), .ZN(G54));
  AND2_X1   g727(.A1(KEYINPUT58), .A2(G475), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n902), .B1(new_n915), .B2(new_n555), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n911), .A2(new_n917), .A3(new_n551), .A4(new_n914), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n911), .A2(new_n551), .A3(new_n914), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT120), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n916), .A2(new_n918), .A3(new_n920), .ZN(G60));
  NAND2_X1  g735(.A1(new_n642), .A2(new_n644), .ZN(new_n922));
  XOR2_X1   g736(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n646), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n922), .B(new_n924), .C1(new_n906), .C2(new_n907), .ZN(new_n925));
  INV_X1    g739(.A(new_n902), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n922), .B1(new_n854), .B2(new_n924), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(G63));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n930));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n851), .B2(new_n852), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n665), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n926), .B1(new_n933), .B2(new_n402), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n851), .A2(new_n852), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n401), .B1(new_n938), .B2(new_n932), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(KEYINPUT61), .A3(new_n926), .A4(new_n934), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(G66));
  INV_X1    g755(.A(new_n595), .ZN(new_n942));
  OAI21_X1  g756(.A(G953), .B1(new_n942), .B2(new_n523), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n835), .A2(new_n836), .A3(new_n829), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n896), .B1(G898), .B2(new_n189), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  AOI21_X1  g761(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n299), .A2(new_n287), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(new_n529), .Z(new_n951));
  AOI211_X1 g765(.A(new_n753), .B(new_n692), .C1(new_n651), .C2(new_n658), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n764), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n806), .B2(new_n809), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n796), .B2(new_n799), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n812), .A2(new_n707), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT62), .B1(new_n703), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n956), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n959), .A3(new_n701), .A4(new_n702), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n955), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n951), .B1(new_n961), .B2(new_n189), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n795), .A2(new_n814), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT123), .B1(new_n964), .B2(new_n880), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n881), .A2(new_n966), .A3(new_n814), .A4(new_n795), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(new_n766), .A3(new_n770), .A4(new_n810), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n800), .A2(new_n958), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT122), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n800), .A2(KEYINPUT122), .A3(new_n958), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n189), .ZN(new_n975));
  INV_X1    g789(.A(new_n951), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(G900), .B2(G953), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n949), .B(new_n963), .C1(new_n975), .C2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n974), .B2(new_n189), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n948), .B1(new_n980), .B2(new_n962), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT63), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n325), .A2(KEYINPUT126), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n985), .A2(new_n694), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n325), .A2(KEYINPUT126), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n839), .B2(new_n843), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n955), .A2(new_n960), .A3(new_n944), .A4(new_n957), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n984), .B(KEYINPUT124), .Z(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n338), .A2(new_n194), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n994), .ZN(new_n996));
  AOI211_X1 g810(.A(KEYINPUT125), .B(new_n996), .C1(new_n991), .C2(new_n992), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n926), .B(new_n989), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n338), .A2(new_n194), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n974), .A2(new_n944), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(new_n992), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n998), .A2(new_n1001), .ZN(G57));
endmodule


