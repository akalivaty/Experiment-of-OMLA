//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1045, new_n1046;
  INV_X1    g000(.A(G113gat), .ZN(new_n202));
  NAND3_X1  g001(.A1(new_n202), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G127gat), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n203), .A2(new_n205), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G113gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n202), .A2(G120gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n205), .A2(new_n207), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n210), .A2(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n225), .A3(KEYINPUT23), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n230), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(KEYINPUT23), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n226), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT23), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n241), .A2(G169gat), .A3(G176gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n235), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT67), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245));
  OR2_X1    g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n245), .B(new_n235), .C1(new_n246), .C2(new_n241), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT25), .B1(new_n236), .B2(KEYINPUT23), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n249), .B1(new_n232), .B2(new_n229), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n239), .A2(new_n240), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n252));
  INV_X1    g051(.A(G183gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT27), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT27), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G183gat), .ZN(new_n256));
  INV_X1    g055(.A(G190gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n246), .A2(KEYINPUT26), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT26), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n236), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n235), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT27), .B(G183gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n257), .A3(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n259), .A2(new_n263), .A3(new_n266), .A4(new_n228), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n219), .B1(new_n251), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT1), .B1(new_n212), .B2(new_n213), .ZN(new_n273));
  XNOR2_X1  g072(.A(G127gat), .B(G134gat), .ZN(new_n274));
  OAI22_X1  g073(.A1(new_n272), .A2(new_n209), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n248), .A2(new_n250), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n223), .A2(new_n224), .A3(new_n241), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n237), .B1(new_n278), .B2(new_n222), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT25), .B1(new_n279), .B2(new_n234), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n275), .B(new_n267), .C1(new_n277), .C2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n269), .A2(new_n271), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT32), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT33), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G15gat), .B(G43gat), .Z(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G99gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n288), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n282), .B(KEYINPUT32), .C1(new_n284), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n269), .A2(new_n281), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT34), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n270), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n294), .B1(new_n293), .B2(new_n270), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n293), .A2(KEYINPUT71), .A3(new_n294), .A4(new_n270), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n296), .B2(new_n295), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n303), .A2(new_n289), .A3(new_n291), .A4(new_n300), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT87), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT2), .ZN(new_n310));
  INV_X1    g109(.A(G141gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(G148gat), .ZN(new_n312));
  INV_X1    g111(.A(G148gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G141gat), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n308), .B(new_n310), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G155gat), .B(G162gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(G141gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(G148gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT77), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n316), .B1(new_n321), .B2(new_n310), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT3), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n315), .A2(new_n317), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(new_n316), .A3(new_n310), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n275), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n219), .A2(KEYINPUT4), .A3(new_n324), .A4(new_n326), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n215), .A2(new_n208), .A3(new_n274), .A4(new_n203), .ZN(new_n331));
  XNOR2_X1  g130(.A(G113gat), .B(G120gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n218), .B1(new_n332), .B2(KEYINPUT1), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n324), .A2(new_n331), .A3(new_n326), .A4(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n275), .B1(new_n318), .B2(new_n322), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n334), .ZN(new_n341));
  INV_X1    g140(.A(new_n329), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT79), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344));
  AOI211_X1 g143(.A(new_n344), .B(new_n329), .C1(new_n340), .C2(new_n334), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n337), .B(new_n339), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n334), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n348), .B(new_n338), .C1(new_n334), .C2(new_n335), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n329), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(G1gat), .B(G29gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT0), .ZN(new_n354));
  XNOR2_X1  g153(.A(G57gat), .B(G85gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT6), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n349), .A2(new_n350), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n342), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n344), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n341), .A2(KEYINPUT79), .A3(new_n342), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n324), .A2(new_n326), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n219), .B1(new_n364), .B2(KEYINPUT3), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n342), .B1(new_n365), .B2(new_n327), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n336), .A2(new_n330), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n338), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n359), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n356), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n358), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n356), .B1(new_n346), .B2(new_n351), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n352), .A2(KEYINPUT6), .A3(new_n357), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n371), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G226gat), .ZN(new_n383));
  INV_X1    g182(.A(G233gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n246), .A2(new_n241), .ZN(new_n387));
  OR2_X1    g186(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(KEYINPUT23), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT65), .B(G169gat), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n235), .B(new_n387), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n229), .A2(new_n231), .A3(new_n233), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n240), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n259), .A2(new_n266), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n263), .A2(new_n228), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n394), .A2(new_n276), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n386), .B1(new_n397), .B2(KEYINPUT29), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n385), .B1(new_n251), .B2(new_n268), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT76), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT74), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT22), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT22), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT74), .ZN(new_n404));
  NAND2_X1  g203(.A1(G211gat), .A2(G218gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G211gat), .ZN(new_n407));
  INV_X1    g206(.A(G218gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(KEYINPUT75), .A3(new_n405), .ZN(new_n410));
  XNOR2_X1  g209(.A(G197gat), .B(G204gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n406), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n406), .B2(new_n411), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n400), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n406), .A2(new_n411), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n409), .A2(new_n405), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(KEYINPUT75), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(KEYINPUT76), .A3(new_n412), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n398), .A2(new_n399), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n398), .B2(new_n399), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n382), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n398), .A2(new_n399), .ZN(new_n425));
  INV_X1    g224(.A(new_n421), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n398), .A2(new_n399), .A3(new_n421), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n381), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT30), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n427), .A2(new_n431), .A3(new_n381), .A4(new_n428), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT35), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT31), .B(G50gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n327), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n420), .A3(new_n415), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT29), .B1(new_n419), .B2(new_n412), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n364), .B1(new_n440), .B2(KEYINPUT3), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n439), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n442), .B(KEYINPUT85), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n416), .A2(new_n417), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n418), .A2(new_n406), .A3(new_n411), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n447), .A2(new_n437), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n364), .B1(new_n449), .B2(KEYINPUT3), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n446), .B1(new_n439), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(G22gat), .B1(new_n444), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n439), .A2(new_n450), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n445), .ZN(new_n454));
  INV_X1    g253(.A(G22gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n441), .A3(new_n443), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n458), .B(KEYINPUT84), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n452), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n452), .B2(new_n457), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n436), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n444), .A2(new_n451), .A3(G22gat), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n455), .B1(new_n454), .B2(new_n456), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n452), .A2(new_n457), .A3(new_n460), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n435), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n378), .A2(new_n434), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n307), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n292), .A2(new_n301), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n463), .B2(new_n468), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT70), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n289), .A2(new_n475), .A3(new_n291), .ZN(new_n476));
  AND4_X1   g275(.A1(KEYINPUT72), .A2(new_n474), .A3(new_n301), .A4(new_n476), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n292), .A2(KEYINPUT70), .B1(new_n303), .B2(new_n300), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT72), .B1(new_n478), .B2(new_n476), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n473), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n376), .A2(new_n373), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n369), .B2(new_n356), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n352), .A2(new_n357), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n358), .A2(KEYINPUT81), .A3(new_n370), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n483), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT83), .B1(new_n490), .B2(new_n433), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n372), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT82), .B1(new_n372), .B2(KEYINPUT6), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n358), .A2(KEYINPUT81), .A3(new_n370), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT81), .B1(new_n358), .B2(new_n370), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n498));
  INV_X1    g297(.A(new_n433), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n473), .B(KEYINPUT88), .C1(new_n477), .C2(new_n479), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n482), .A2(new_n491), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n471), .B1(new_n502), .B2(KEYINPUT35), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n427), .A2(KEYINPUT86), .A3(new_n428), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT37), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT38), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n427), .A2(KEYINPUT86), .A3(new_n507), .A4(new_n428), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n505), .A2(new_n506), .A3(new_n382), .A4(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n382), .A3(new_n508), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT38), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n377), .A2(new_n429), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT40), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n328), .B(new_n348), .C1(new_n334), .C2(new_n335), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n342), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n356), .B1(new_n515), .B2(KEYINPUT39), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT39), .B1(new_n341), .B2(new_n342), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n514), .B2(new_n342), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n513), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n356), .B2(new_n369), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n516), .A2(new_n513), .A3(new_n518), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n522), .A2(new_n433), .B1(new_n468), .B2(new_n463), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n305), .A2(KEYINPUT73), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT73), .B1(new_n305), .B2(new_n525), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n472), .A2(new_n525), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n479), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n478), .A2(KEYINPUT72), .A3(new_n476), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n524), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n469), .B1(new_n491), .B2(new_n500), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n503), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n455), .A2(G15gat), .ZN(new_n539));
  INV_X1    g338(.A(G15gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G22gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT90), .ZN(new_n546));
  INV_X1    g345(.A(G1gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT92), .ZN(new_n549));
  INV_X1    g348(.A(G8gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n545), .A2(KEYINPUT90), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n539), .A2(new_n541), .A3(KEYINPUT90), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n554), .A2(KEYINPUT16), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n547), .B1(new_n554), .B2(KEYINPUT91), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n557), .B(G1gat), .C1(new_n552), .C2(new_n553), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n551), .A2(new_n555), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(G8gat), .B1(new_n548), .B2(KEYINPUT92), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(KEYINPUT16), .B2(new_n554), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT91), .B1(new_n544), .B2(new_n546), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(G1gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n560), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT15), .ZN(new_n566));
  INV_X1    g365(.A(G29gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT14), .B(G29gat), .Z(new_n569));
  OAI211_X1 g368(.A(new_n566), .B(new_n568), .C1(new_n569), .C2(G36gat), .ZN(new_n570));
  OR2_X1    g369(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n572));
  AOI21_X1  g371(.A(G36gat), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n568), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT15), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G43gat), .B(G50gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n570), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n578), .B(KEYINPUT15), .C1(new_n573), .C2(new_n574), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT89), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT17), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT89), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n577), .A2(new_n583), .A3(new_n579), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n577), .A2(KEYINPUT17), .A3(new_n579), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n565), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n577), .A2(new_n583), .A3(new_n579), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n583), .B1(new_n577), .B2(new_n579), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(new_n559), .A3(new_n564), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n565), .B1(new_n590), .B2(new_n589), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n592), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n588), .B(KEYINPUT13), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n587), .A2(KEYINPUT18), .A3(new_n588), .A4(new_n592), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n595), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G197gat), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT11), .B(G169gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n595), .A2(new_n606), .A3(new_n600), .A4(new_n599), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n538), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n615));
  XNOR2_X1  g414(.A(G134gat), .B(G162gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT99), .Z(new_n618));
  NAND2_X1  g417(.A1(G85gat), .A2(G92gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT7), .ZN(new_n620));
  OR2_X1    g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(KEYINPUT97), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(KEYINPUT8), .B2(new_n622), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n620), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT97), .B1(new_n621), .B2(new_n622), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n629), .A2(new_n620), .A3(new_n623), .A4(new_n625), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n586), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n591), .B2(new_n582), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n581), .A2(new_n584), .A3(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT98), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n591), .A2(new_n631), .B1(KEYINPUT41), .B2(new_n614), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n585), .A2(new_n586), .A3(new_n632), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n638), .A2(new_n642), .A3(new_n257), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n257), .B1(new_n638), .B2(new_n642), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n643), .A2(new_n644), .A3(G218gat), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n634), .A2(new_n637), .A3(KEYINPUT98), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n641), .B1(new_n639), .B2(new_n640), .ZN(new_n647));
  OAI21_X1  g446(.A(G190gat), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n638), .A2(new_n642), .A3(new_n257), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n408), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n618), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G218gat), .B1(new_n643), .B2(new_n644), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(new_n408), .A3(new_n649), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n617), .A2(KEYINPUT99), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G183gat), .B(G211gat), .ZN(new_n657));
  INV_X1    g456(.A(G71gat), .ZN(new_n658));
  INV_X1    g457(.A(G78gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G71gat), .A2(G78gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT9), .ZN(new_n663));
  XNOR2_X1  g462(.A(G57gat), .B(G64gat), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT93), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(G57gat), .A2(G64gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(G57gat), .A2(G64gat), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(KEYINPUT93), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n662), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT94), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n667), .A2(KEYINPUT94), .A3(new_n668), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT9), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n672), .A2(new_n673), .B1(new_n661), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT95), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n668), .ZN(new_n677));
  NOR2_X1   g476(.A1(G57gat), .A2(G64gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n665), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n669), .A3(KEYINPUT9), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n661), .A3(new_n660), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT95), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n674), .A2(new_n661), .ZN(new_n683));
  INV_X1    g482(.A(new_n673), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT94), .B1(new_n667), .B2(new_n668), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n681), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT21), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n676), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(G231gat), .A2(G233gat), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n206), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n206), .B1(new_n691), .B2(new_n692), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n657), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n695), .ZN(new_n697));
  INV_X1    g496(.A(new_n657), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n698), .A3(new_n693), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n700));
  INV_X1    g499(.A(G155gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT96), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n676), .A2(new_n687), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT21), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n565), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n565), .B2(new_n705), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n702), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n708), .ZN(new_n710));
  INV_X1    g509(.A(new_n702), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n696), .A2(new_n699), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n696), .A2(new_n699), .B1(new_n709), .B2(new_n712), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n656), .A2(KEYINPUT100), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT100), .B1(new_n656), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g517(.A(G120gat), .B(G148gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(G176gat), .B(G204gat), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n719), .B(new_n720), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT102), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n704), .A2(KEYINPUT10), .A3(new_n631), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n628), .A2(new_n630), .B1(new_n681), .B2(new_n686), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n704), .B2(new_n632), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n725), .B2(KEYINPUT10), .ZN(new_n726));
  NAND2_X1  g525(.A1(G230gat), .A2(G233gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n727), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n722), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n721), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n731), .B2(KEYINPUT101), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(KEYINPUT101), .B2(new_n731), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n735), .B2(new_n729), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n717), .A2(new_n718), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n613), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n497), .A2(KEYINPUT103), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n497), .A2(KEYINPUT103), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n547), .ZN(G1324gat));
  NOR2_X1   g543(.A1(new_n738), .A2(new_n499), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT16), .B(G8gat), .Z(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n550), .B2(new_n745), .ZN(new_n748));
  MUX2_X1   g547(.A(new_n747), .B(new_n748), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g548(.A1(new_n529), .A2(new_n534), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G15gat), .B1(new_n738), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n306), .A2(new_n540), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n738), .B2(new_n753), .ZN(G1326gat));
  INV_X1    g553(.A(new_n469), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n613), .A2(new_n755), .A3(new_n737), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT43), .B(G22gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1327gat));
  NOR3_X1   g557(.A1(new_n656), .A2(new_n716), .A3(new_n736), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n613), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n760), .A2(G29gat), .A3(new_n742), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT45), .Z(new_n762));
  AND3_X1   g561(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n763));
  INV_X1    g562(.A(new_n618), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n652), .B2(new_n653), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  OAI211_X1 g565(.A(KEYINPUT44), .B(new_n766), .C1(new_n503), .C2(new_n537), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n736), .B(KEYINPUT104), .Z(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n769), .A2(new_n612), .A3(new_n716), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n771));
  INV_X1    g570(.A(new_n471), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n488), .A2(new_n489), .ZN(new_n774));
  AOI211_X1 g573(.A(KEYINPUT83), .B(new_n433), .C1(new_n774), .C2(new_n494), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n498), .B1(new_n497), .B2(new_n499), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n755), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT105), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n305), .A2(new_n525), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT73), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n526), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n530), .B1(new_n477), .B2(new_n479), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n782), .A2(new_n783), .B1(new_n512), .B2(new_n523), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n785), .B(new_n755), .C1(new_n775), .C2(new_n776), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n778), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n656), .B1(new_n773), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n767), .B(new_n770), .C1(new_n788), .C2(KEYINPUT44), .ZN(new_n789));
  OAI21_X1  g588(.A(G29gat), .B1(new_n789), .B2(new_n742), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n762), .A2(new_n790), .ZN(G1328gat));
  NOR3_X1   g590(.A1(new_n760), .A2(G36gat), .A3(new_n499), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n789), .A2(new_n499), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT107), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G36gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n795), .A2(KEYINPUT107), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(G1329gat));
  OR3_X1    g598(.A1(new_n760), .A2(G43gat), .A3(new_n307), .ZN(new_n800));
  OAI21_X1  g599(.A(G43gat), .B1(new_n789), .B2(new_n751), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT108), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(G1330gat));
  OAI21_X1  g603(.A(G50gat), .B1(new_n789), .B2(new_n469), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n469), .A2(G50gat), .ZN(new_n806));
  OAI221_X1 g605(.A(new_n805), .B1(KEYINPUT109), .B2(KEYINPUT48), .C1(new_n760), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1331gat));
  INV_X1    g608(.A(new_n612), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n773), .B2(new_n787), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n717), .A2(new_n718), .A3(new_n768), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n742), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n499), .ZN(new_n816));
  NOR2_X1   g615(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n817));
  AND2_X1   g616(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n816), .B2(new_n817), .ZN(G1333gat));
  OAI21_X1  g619(.A(G71gat), .B1(new_n813), .B2(new_n751), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n306), .A2(new_n658), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n813), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g623(.A1(new_n813), .A2(new_n469), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(new_n659), .ZN(G1335gat));
  INV_X1    g625(.A(new_n736), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n810), .A2(new_n716), .A3(new_n827), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n767), .B(new_n828), .C1(new_n788), .C2(KEYINPUT44), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n784), .B1(new_n536), .B2(new_n785), .ZN(new_n832));
  INV_X1    g631(.A(new_n786), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n766), .B1(new_n834), .B2(new_n503), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT44), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n837), .A2(KEYINPUT110), .A3(new_n767), .A4(new_n828), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G85gat), .B1(new_n839), .B2(new_n742), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n656), .A2(new_n716), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n612), .B(new_n841), .C1(new_n834), .C2(new_n503), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n811), .A2(KEYINPUT51), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT111), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n742), .A2(G85gat), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n848), .A2(new_n736), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n840), .A2(new_n851), .ZN(G1336gat));
  NOR2_X1   g651(.A1(new_n499), .A2(G92gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n846), .A2(new_n769), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n855));
  OAI21_X1  g654(.A(G92gat), .B1(new_n829), .B2(new_n499), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n831), .A2(new_n838), .A3(new_n433), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G92gat), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT52), .B1(new_n859), .B2(KEYINPUT112), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n854), .A2(KEYINPUT112), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(G92gat), .B2(new_n858), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n857), .B1(new_n860), .B2(new_n862), .ZN(G1337gat));
  OAI21_X1  g662(.A(G99gat), .B1(new_n839), .B2(new_n751), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n307), .A2(G99gat), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n848), .A2(new_n736), .A3(new_n849), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(G1338gat));
  NAND3_X1  g666(.A1(new_n831), .A2(new_n838), .A3(new_n755), .ZN(new_n868));
  XOR2_X1   g667(.A(KEYINPUT113), .B(G106gat), .Z(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n469), .A2(G106gat), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n842), .A2(new_n843), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT51), .B1(new_n811), .B2(new_n841), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n769), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n846), .A2(KEYINPUT114), .A3(new_n769), .A4(new_n871), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT53), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n869), .B1(new_n829), .B2(new_n469), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n874), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(G1339gat));
  OAI21_X1  g682(.A(new_n733), .B1(new_n728), .B2(KEYINPUT54), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n726), .B2(new_n727), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n730), .B(new_n723), .C1(new_n725), .C2(KEYINPUT10), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n887), .A2(KEYINPUT115), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT115), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT55), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n891), .A2(new_n892), .B1(new_n608), .B2(new_n610), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n735), .A2(new_n729), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n728), .A2(KEYINPUT54), .A3(new_n888), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n887), .A2(KEYINPUT115), .A3(new_n888), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n884), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n899), .B2(KEYINPUT55), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n588), .B1(new_n587), .B2(new_n592), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n902));
  OAI22_X1  g701(.A1(new_n901), .A2(new_n902), .B1(new_n597), .B2(new_n598), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT116), .B(new_n588), .C1(new_n587), .C2(new_n592), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n605), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n610), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n893), .A2(new_n900), .B1(new_n906), .B2(new_n736), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n651), .A2(new_n906), .A3(new_n655), .A4(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n900), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n907), .A2(new_n766), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n905), .A2(new_n610), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n892), .B2(new_n891), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n766), .A2(new_n900), .A3(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n916), .B(KEYINPUT117), .C1(new_n766), .C2(new_n907), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n913), .A2(new_n715), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n737), .A2(new_n612), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n741), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n482), .A2(new_n501), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n921), .A2(new_n433), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(G113gat), .B1(new_n924), .B2(new_n810), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n716), .B1(new_n911), .B2(new_n912), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n926), .A2(new_n917), .B1(new_n737), .B2(new_n612), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n755), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n741), .A2(new_n499), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n307), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n202), .A3(new_n612), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n925), .A2(new_n932), .ZN(G1340gat));
  NAND2_X1  g732(.A1(new_n736), .A2(new_n211), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT118), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n924), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G120gat), .B1(new_n931), .B2(new_n768), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT119), .Z(G1341gat));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n206), .A3(new_n716), .ZN(new_n940));
  OAI21_X1  g739(.A(G127gat), .B1(new_n931), .B2(new_n715), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1342gat));
  NOR2_X1   g741(.A1(new_n921), .A2(new_n923), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n656), .A2(G134gat), .A3(new_n433), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT56), .ZN(new_n946));
  OAI21_X1  g745(.A(G134gat), .B1(new_n931), .B2(new_n656), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n943), .A2(new_n948), .A3(new_n944), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT120), .ZN(G1343gat));
  OAI21_X1  g750(.A(KEYINPUT121), .B1(new_n927), .B2(new_n742), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n920), .A2(new_n953), .A3(new_n741), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n750), .A2(new_n469), .ZN(new_n955));
  AND4_X1   g754(.A1(new_n499), .A2(new_n952), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n612), .A2(G141gat), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n929), .A2(new_n750), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT57), .B1(new_n920), .B2(new_n755), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT57), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n469), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n911), .A2(new_n715), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n919), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n810), .B(new_n958), .C1(new_n959), .C2(new_n964), .ZN(new_n965));
  AOI22_X1  g764(.A1(new_n956), .A2(new_n957), .B1(new_n965), .B2(G141gat), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n967), .B1(new_n965), .B2(G141gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n966), .A2(KEYINPUT58), .A3(new_n968), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n954), .A2(new_n955), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n970), .A2(new_n499), .A3(new_n952), .A4(new_n957), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n965), .A2(G141gat), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n971), .B(new_n972), .C1(KEYINPUT122), .C2(KEYINPUT58), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n969), .A2(new_n974), .ZN(G1344gat));
  OR2_X1    g774(.A1(new_n959), .A2(new_n964), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n929), .A2(new_n750), .A3(new_n827), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT59), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n469), .B1(new_n919), .B2(new_n963), .ZN(new_n980));
  OAI22_X1  g779(.A1(new_n980), .A2(KEYINPUT57), .B1(new_n927), .B2(new_n962), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(new_n977), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n978), .A2(new_n313), .ZN(new_n983));
  AOI22_X1  g782(.A1(new_n976), .A2(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n978), .B1(new_n956), .B2(new_n736), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n985), .B2(G148gat), .ZN(G1345gat));
  NAND2_X1  g785(.A1(new_n976), .A2(new_n958), .ZN(new_n987));
  OAI21_X1  g786(.A(G155gat), .B1(new_n987), .B2(new_n715), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n956), .A2(new_n701), .A3(new_n716), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1346gat));
  OAI21_X1  g789(.A(G162gat), .B1(new_n987), .B2(new_n656), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n656), .A2(G162gat), .A3(new_n433), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n970), .A2(new_n952), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1347gat));
  NOR2_X1   g793(.A1(new_n927), .A2(new_n741), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n923), .A2(new_n499), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n997), .A2(new_n391), .A3(new_n612), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n742), .A2(new_n433), .A3(new_n306), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT123), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n928), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(new_n810), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n998), .B1(G169gat), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT124), .ZN(G1348gat));
  INV_X1    g804(.A(new_n997), .ZN(new_n1006));
  AOI21_X1  g805(.A(G176gat), .B1(new_n1006), .B2(new_n736), .ZN(new_n1007));
  NOR3_X1   g806(.A1(new_n1001), .A2(new_n225), .A3(new_n768), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1349gat));
  OAI21_X1  g808(.A(G183gat), .B1(new_n1001), .B2(new_n715), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n716), .A2(new_n264), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1010), .B1(new_n997), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g811(.A(new_n1012), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n928), .A2(new_n1000), .A3(new_n766), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1014), .B1(new_n1015), .B2(G190gat), .ZN(new_n1016));
  INV_X1    g815(.A(KEYINPUT61), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1015), .A2(new_n1014), .A3(G190gat), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1021));
  NOR3_X1   g820(.A1(new_n997), .A2(G190gat), .A3(new_n656), .ZN(new_n1022));
  NOR2_X1   g821(.A1(new_n1022), .A2(KEYINPUT125), .ZN(new_n1023));
  AND2_X1   g822(.A1(new_n1022), .A2(KEYINPUT125), .ZN(new_n1024));
  OAI211_X1 g823(.A(new_n1020), .B(new_n1021), .C1(new_n1023), .C2(new_n1024), .ZN(G1351gat));
  AND3_X1   g824(.A1(new_n995), .A2(new_n433), .A3(new_n955), .ZN(new_n1026));
  AOI21_X1  g825(.A(G197gat), .B1(new_n1026), .B2(new_n810), .ZN(new_n1027));
  NOR3_X1   g826(.A1(new_n741), .A2(new_n750), .A3(new_n499), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n981), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g828(.A(new_n1029), .ZN(new_n1030));
  AND2_X1   g829(.A1(new_n810), .A2(G197gat), .ZN(new_n1031));
  AOI21_X1  g830(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(G1352gat));
  INV_X1    g831(.A(G204gat), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1026), .A2(new_n1033), .A3(new_n736), .ZN(new_n1034));
  XNOR2_X1  g833(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1035));
  OR2_X1    g834(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g835(.A(G204gat), .B1(new_n1029), .B2(new_n768), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1038));
  NAND3_X1  g837(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(G1353gat));
  NAND3_X1  g838(.A1(new_n1026), .A2(new_n407), .A3(new_n716), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1030), .A2(new_n716), .ZN(new_n1041));
  AND3_X1   g840(.A1(new_n1041), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1042));
  AOI21_X1  g841(.A(KEYINPUT63), .B1(new_n1041), .B2(G211gat), .ZN(new_n1043));
  OAI21_X1  g842(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(G1354gat));
  OAI21_X1  g843(.A(G218gat), .B1(new_n1029), .B2(new_n656), .ZN(new_n1045));
  NAND3_X1  g844(.A1(new_n1026), .A2(new_n408), .A3(new_n766), .ZN(new_n1046));
  NAND2_X1  g845(.A1(new_n1045), .A2(new_n1046), .ZN(G1355gat));
endmodule


