//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n462), .A2(G2105), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n466), .A2(G2105), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NOR3_X1   g043(.A1(new_n462), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n460), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT68), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n474), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT69), .Z(new_n483));
  NAND3_X1  g058(.A1(new_n471), .A2(G2105), .A3(new_n473), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n480), .B(new_n483), .C1(G124), .C2(new_n485), .ZN(G162));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  OR2_X1    g062(.A1(KEYINPUT70), .A2(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT70), .A2(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n472), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  OAI22_X1  g066(.A1(new_n484), .A2(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n472), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  AOI211_X1 g070(.A(new_n495), .B(new_n464), .C1(new_n493), .C2(new_n494), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n471), .A2(KEYINPUT71), .A3(new_n473), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(new_n460), .A3(G2104), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n473), .A2(new_n501), .A3(new_n463), .A4(new_n498), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n499), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n496), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n499), .A2(KEYINPUT72), .A3(new_n504), .A4(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n492), .B1(new_n507), .B2(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT74), .Z(new_n519));
  NAND2_X1  g094(.A1(new_n511), .A2(G62), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(new_n515), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(new_n512), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n523), .B(new_n525), .C1(new_n530), .C2(KEYINPUT75), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n530), .A2(KEYINPUT75), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(G52), .A2(new_n524), .B1(new_n512), .B2(G90), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n511), .A2(G64), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n517), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n535), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(G171));
  NAND2_X1  g116(.A1(new_n512), .A2(G81), .ZN(new_n542));
  INV_X1    g117(.A(G43), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(new_n515), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n517), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT77), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT77), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OR3_X1    g132(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n515), .B2(new_n557), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT78), .Z(new_n561));
  NAND2_X1  g136(.A1(new_n512), .A2(G91), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n517), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n512), .A2(G87), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT79), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n511), .A2(G74), .ZN(new_n572));
  AOI22_X1  g147(.A1(G49), .A2(new_n524), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(new_n511), .A2(G61), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(KEYINPUT80), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n575), .A2(KEYINPUT80), .B1(G73), .B2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n517), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(G48), .A2(new_n524), .B1(new_n512), .B2(G86), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n578), .A2(new_n579), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(G47), .A2(new_n524), .B1(new_n512), .B2(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n517), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(new_n512), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  NAND2_X1  g165(.A1(new_n511), .A2(G66), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n517), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(G54), .B2(new_n524), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(G171), .ZN(G284));
  OAI21_X1  g173(.A(new_n597), .B1(new_n596), .B2(G171), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n561), .A2(new_n565), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(new_n595), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT82), .B(G559), .Z(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(G860), .B2(new_n605), .ZN(G148));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g185(.A1(G99), .A2(G2105), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n611), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n612));
  INV_X1    g187(.A(G123), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n484), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(G135), .B2(new_n481), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(G2096), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(G2096), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n636), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n643), .B2(new_n640), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n646), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1971), .B(G1976), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n653), .A2(new_n658), .A3(new_n656), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n653), .A2(new_n658), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n661));
  AOI211_X1 g236(.A(new_n657), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n660), .B2(new_n661), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1981), .B(G1986), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G229));
  INV_X1    g244(.A(G16), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G24), .ZN(new_n671));
  INV_X1    g246(.A(G290), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n672), .B2(new_n670), .ZN(new_n673));
  INV_X1    g248(.A(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(G25), .A2(G29), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n481), .A2(G131), .ZN(new_n677));
  INV_X1    g252(.A(G119), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n472), .A2(G107), .ZN(new_n679));
  OAI21_X1  g254(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n680));
  OAI22_X1  g255(.A1(new_n484), .A2(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n676), .B1(new_n682), .B2(G29), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT35), .B(G1991), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n675), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n683), .B2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G305), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G16), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G6), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT32), .B(G1981), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n692), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n670), .A2(G23), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G288), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n670), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n670), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1971), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n696), .A2(new_n697), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n693), .A2(new_n694), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n687), .B1(new_n705), .B2(KEYINPUT34), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT86), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(KEYINPUT34), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT36), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n670), .A2(G20), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT23), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n601), .B2(new_n670), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(G1956), .Z(new_n714));
  NOR2_X1   g289(.A1(G171), .A2(new_n670), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G5), .B2(new_n670), .ZN(new_n716));
  INV_X1    g291(.A(G1961), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT91), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n551), .A2(new_n670), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n670), .B2(G19), .ZN(new_n722));
  INV_X1    g297(.A(G1341), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n722), .A2(new_n723), .B1(new_n716), .B2(new_n717), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n670), .A2(G21), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G168), .B2(new_n670), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G1966), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT90), .Z(new_n728));
  OAI211_X1 g303(.A(new_n724), .B(new_n728), .C1(new_n723), .C2(new_n722), .ZN(new_n729));
  INV_X1    g304(.A(G2078), .ZN(new_n730));
  NAND2_X1  g305(.A1(G164), .A2(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G27), .B2(G29), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n720), .B(new_n729), .C1(new_n730), .C2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  INV_X1    g310(.A(G139), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n474), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT88), .ZN(new_n738));
  NAND2_X1  g313(.A1(G115), .A2(G2104), .ZN(new_n739));
  INV_X1    g314(.A(G127), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n464), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n738), .B1(G2105), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G29), .B2(G33), .ZN(new_n744));
  INV_X1    g319(.A(G2072), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  INV_X1    g322(.A(G34), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n748), .B2(KEYINPUT24), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(KEYINPUT24), .B2(new_n748), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n476), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT26), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n757), .A2(new_n758), .B1(G105), .B2(new_n467), .ZN(new_n759));
  INV_X1    g334(.A(G129), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n484), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G141), .B2(new_n481), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(new_n751), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n751), .B2(G32), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n754), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n746), .A2(new_n747), .A3(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT89), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n751), .A2(G35), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT92), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n751), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT29), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(G2090), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(G2090), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n764), .A2(new_n765), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n726), .B2(G1966), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G28), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n751), .B1(new_n778), .B2(G28), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n777), .B1(new_n779), .B2(new_n780), .C1(new_n616), .C2(new_n751), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n670), .A2(G4), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n604), .B2(new_n670), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G1348), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n783), .A2(G1348), .B1(new_n753), .B2(new_n752), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n751), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  INV_X1    g364(.A(G128), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n472), .A2(G116), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n792));
  OAI22_X1  g367(.A1(new_n484), .A2(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G140), .B2(new_n481), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(new_n751), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT87), .B(G2067), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n776), .A2(new_n786), .A3(new_n787), .A4(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n773), .A2(new_n774), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n732), .A2(new_n730), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n733), .A2(new_n768), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n710), .A2(new_n801), .ZN(G311));
  OR2_X1    g377(.A1(new_n710), .A2(new_n801), .ZN(G150));
  NAND2_X1  g378(.A1(new_n604), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT96), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT38), .Z(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT93), .B(G93), .ZN(new_n807));
  AOI22_X1  g382(.A1(G55), .A2(new_n524), .B1(new_n512), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n517), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n812), .B(new_n813), .C1(new_n546), .C2(new_n544), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n548), .A2(new_n549), .A3(new_n810), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n814), .A2(new_n815), .A3(KEYINPUT95), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT95), .B1(new_n814), .B2(new_n815), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n806), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n821));
  AOI21_X1  g396(.A(G860), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n812), .A2(new_n813), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(G145));
  XOR2_X1   g402(.A(KEYINPUT98), .B(G37), .Z(new_n828));
  INV_X1    g403(.A(KEYINPUT97), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n742), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n762), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n485), .A2(G130), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n472), .A2(G118), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G142), .B2(new_n481), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(new_n620), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n831), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n504), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT4), .B1(new_n502), .B2(new_n503), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n506), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n496), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n508), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n492), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n794), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n682), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n838), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n615), .B(new_n476), .ZN(new_n849));
  XNOR2_X1  g424(.A(G162), .B(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n848), .A2(new_n850), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n828), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g429(.A1(new_n824), .A2(new_n596), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n819), .B(new_n607), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n601), .A2(new_n604), .ZN(new_n857));
  NAND2_X1  g432(.A1(G299), .A2(new_n595), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(KEYINPUT41), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(new_n862), .A3(new_n858), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n860), .B1(new_n856), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(G305), .B(G166), .ZN(new_n866));
  XNOR2_X1  g441(.A(G288), .B(G290), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT99), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n867), .A2(KEYINPUT99), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n869), .B1(new_n872), .B2(new_n866), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT42), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n865), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n855), .B1(new_n875), .B2(new_n596), .ZN(G295));
  OAI21_X1  g451(.A(new_n855), .B1(new_n875), .B2(new_n596), .ZN(G331));
  OAI21_X1  g452(.A(G168), .B1(new_n817), .B2(new_n818), .ZN(new_n878));
  INV_X1    g453(.A(new_n818), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(G286), .A3(new_n816), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G301), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n880), .A3(G171), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n882), .A2(new_n858), .A3(new_n857), .A4(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n878), .A2(new_n880), .A3(G171), .ZN(new_n885));
  AOI21_X1  g460(.A(G171), .B1(new_n878), .B2(new_n880), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n864), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n873), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n887), .A3(new_n873), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n828), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n859), .A2(KEYINPUT100), .A3(KEYINPUT41), .ZN(new_n895));
  OAI221_X1 g470(.A(new_n895), .B1(KEYINPUT100), .B2(new_n864), .C1(new_n885), .C2(new_n886), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n873), .B1(new_n896), .B2(new_n884), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  MUX2_X1   g474(.A(new_n893), .B(new_n898), .S(new_n899), .Z(new_n900));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n894), .B2(new_n897), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n895), .B1(new_n864), .B2(KEYINPUT100), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(new_n882), .B2(new_n883), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n885), .A2(new_n886), .A3(new_n859), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n889), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n908), .A2(KEYINPUT101), .A3(new_n828), .A4(new_n892), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(KEYINPUT43), .A3(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n890), .A2(new_n899), .A3(new_n891), .A4(new_n892), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n911), .A2(KEYINPUT44), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT102), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT102), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n902), .B1(new_n913), .B2(new_n914), .ZN(G397));
  INV_X1    g490(.A(G1384), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n845), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT45), .ZN(new_n918));
  NAND2_X1  g493(.A1(G160), .A2(G40), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(G1996), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n762), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(KEYINPUT104), .Z(new_n924));
  XNOR2_X1  g499(.A(new_n921), .B(KEYINPUT105), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n794), .B(G2067), .ZN(new_n926));
  INV_X1    g501(.A(G1996), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(new_n927), .B2(new_n762), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n924), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n677), .A2(new_n681), .A3(new_n685), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n682), .A2(new_n684), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n921), .A2(new_n674), .A3(new_n672), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n921), .A2(G1986), .A3(G290), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT103), .Z(new_n937));
  NOR2_X1   g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT106), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT63), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT113), .ZN(new_n941));
  INV_X1    g516(.A(G8), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n845), .A2(KEYINPUT45), .A3(new_n916), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n920), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT107), .B1(G164), .B2(G1384), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n845), .A2(new_n946), .A3(new_n916), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n944), .B1(new_n948), .B2(new_n918), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT112), .B1(new_n949), .B2(G1966), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n946), .B1(new_n845), .B2(new_n916), .ZN(new_n951));
  AOI211_X1 g526(.A(KEYINPUT107), .B(G1384), .C1(new_n843), .C2(new_n844), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n918), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(G164), .A2(G1384), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n919), .B1(new_n954), .B2(KEYINPUT45), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n957));
  INV_X1    g532(.A(G1966), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n950), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n945), .A2(new_n961), .A3(new_n947), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n917), .B2(KEYINPUT50), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n945), .A2(new_n947), .A3(new_n963), .A4(new_n961), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n919), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n753), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n942), .B1(new_n960), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n941), .B1(new_n969), .B2(G168), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n950), .A2(new_n959), .B1(new_n967), .B2(new_n753), .ZN(new_n971));
  NOR4_X1   g546(.A1(new_n971), .A2(KEYINPUT113), .A3(new_n942), .A4(G286), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(G303), .A2(G8), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT55), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n918), .B1(G164), .B2(G1384), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n977), .A2(new_n920), .A3(new_n943), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(G1971), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  AOI211_X1 g555(.A(G2090), .B(new_n919), .C1(new_n965), .C2(new_n966), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(KEYINPUT109), .ZN(new_n982));
  INV_X1    g557(.A(G2090), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n967), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(G8), .B(new_n976), .C1(new_n982), .C2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n920), .B1(new_n917), .B2(KEYINPUT50), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(KEYINPUT50), .B2(new_n948), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n983), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n980), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n976), .B1(new_n991), .B2(G8), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n993));
  INV_X1    g568(.A(G1981), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n583), .A2(new_n994), .A3(new_n580), .A4(new_n581), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n582), .A2(KEYINPUT110), .A3(new_n994), .A4(new_n583), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n688), .A2(new_n994), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n993), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n945), .A2(new_n920), .A3(new_n947), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(new_n942), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n999), .B(KEYINPUT49), .C1(new_n994), .C2(new_n688), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G288), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G1976), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(G288), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1005), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1003), .A2(G8), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT52), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1007), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n992), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n987), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n940), .B1(new_n973), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n960), .A2(new_n968), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(G8), .A3(G168), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT113), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n969), .A2(new_n941), .A3(G168), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1007), .A2(new_n1012), .A3(KEYINPUT63), .A4(new_n1014), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n942), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1027), .B2(new_n976), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n982), .B2(new_n986), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n975), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1023), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1018), .A2(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1007), .A2(new_n1010), .A3(new_n1008), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1005), .B1(new_n1033), .B2(new_n1000), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n987), .B2(new_n1015), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1034), .B(KEYINPUT111), .C1(new_n987), .C2(new_n1015), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n978), .A2(new_n730), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT119), .B(G1961), .Z(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1042), .B1(new_n967), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT123), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n977), .A2(new_n943), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT53), .B1(KEYINPUT122), .B2(G2078), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(KEYINPUT122), .B2(G2078), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1046), .A2(new_n1047), .A3(G301), .A4(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1042), .B(new_n1053), .C1(new_n967), .C2(new_n1044), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT123), .B1(new_n1055), .B2(G171), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n953), .A2(new_n730), .A3(new_n955), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n953), .A2(new_n955), .A3(KEYINPUT118), .A4(new_n730), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1059), .A2(KEYINPUT53), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(G171), .B1(new_n1061), .B2(new_n1045), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1054), .A2(new_n1056), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT124), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(KEYINPUT124), .A3(new_n1064), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n978), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n565), .A2(new_n1072), .A3(new_n560), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1071), .B(new_n1075), .C1(new_n989), .C2(G1956), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n965), .A2(new_n966), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n920), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n785), .ZN(new_n1079));
  INV_X1    g654(.A(G2067), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1004), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n595), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1075), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT50), .B1(new_n951), .B2(new_n952), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n919), .B1(new_n954), .B2(new_n961), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1956), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n977), .A2(new_n920), .A3(new_n943), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1070), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1083), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(KEYINPUT114), .B(new_n1083), .C1(new_n1086), .C2(new_n1089), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1076), .B1(new_n1082), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT60), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1096));
  OAI211_X1 g671(.A(KEYINPUT60), .B(new_n1081), .C1(new_n967), .C2(G1348), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n604), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1079), .A2(KEYINPUT60), .A3(new_n595), .A4(new_n1081), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1090), .A2(new_n1076), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT115), .B(G1996), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(new_n723), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n978), .A2(new_n1103), .B1(new_n1003), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT59), .B1(new_n1106), .B2(new_n550), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1003), .A2(new_n1105), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1103), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1087), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1108), .B(new_n551), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1101), .A2(new_n1102), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1092), .A2(new_n1093), .A3(KEYINPUT61), .A4(new_n1076), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1095), .B1(new_n1100), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1078), .A2(new_n1043), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1059), .A2(KEYINPUT53), .A3(new_n1060), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(G301), .A4(new_n1042), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1064), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1055), .A2(new_n1122), .A3(G171), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1046), .A2(KEYINPUT125), .A3(G301), .A4(new_n1118), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1055), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT126), .B1(new_n1125), .B2(G301), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n987), .A2(new_n1016), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n960), .A2(G168), .A3(new_n968), .ZN(new_n1129));
  AND2_X1   g704(.A1(KEYINPUT117), .A2(G8), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1019), .A2(G8), .A3(G286), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n1134), .A3(new_n1130), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1116), .A2(new_n1127), .A3(new_n1128), .A4(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1032), .B(new_n1039), .C1(new_n1069), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1133), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1134), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT62), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G301), .B1(new_n1046), .B2(new_n1118), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n987), .A2(new_n1016), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1132), .A2(new_n1144), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT127), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n939), .B1(new_n1138), .B2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n922), .B(KEYINPUT46), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n762), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n925), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT47), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n935), .B(KEYINPUT48), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n933), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n929), .A2(new_n930), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n794), .A2(new_n1080), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(new_n925), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1151), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g738(.A(G227), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1165), .A2(G319), .ZN(new_n1166));
  NOR3_X1   g740(.A1(G229), .A2(G401), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g741(.A1(new_n900), .A2(new_n853), .A3(new_n1167), .ZN(G225));
  INV_X1    g742(.A(G225), .ZN(G308));
endmodule


