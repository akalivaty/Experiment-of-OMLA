//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT10), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT65), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n191), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n195), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(new_n198), .A3(new_n191), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n192), .A2(new_n194), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n196), .A2(new_n198), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n201), .A2(new_n202), .B1(new_n205), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT80), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G104), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n215), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G107), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  OR3_X1    g035(.A1(new_n212), .A2(KEYINPUT3), .A3(G107), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n218), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n217), .B1(G104), .B2(new_n216), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G101), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n211), .A2(KEYINPUT81), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n223), .A2(new_n225), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n205), .A2(new_n210), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n207), .A2(new_n209), .A3(new_n202), .A4(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n228), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n189), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n223), .A2(KEYINPUT4), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n218), .A2(new_n220), .A3(new_n222), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G101), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n235), .B(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT0), .A4(G128), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n203), .B1(new_n206), .B2(G143), .ZN(new_n240));
  XOR2_X1   g054(.A(KEYINPUT0), .B(G128), .Z(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n246));
  NOR4_X1   g060(.A1(new_n195), .A2(new_n199), .A3(KEYINPUT1), .A4(new_n200), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT65), .B(G146), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT1), .B1(new_n248), .B2(new_n190), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT68), .B(G128), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n190), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n249), .A2(new_n250), .B1(new_n251), .B2(new_n203), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n246), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n202), .B1(new_n206), .B2(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n200), .A2(KEYINPUT68), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n240), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT69), .A3(new_n231), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n226), .A2(KEYINPUT82), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n223), .A2(new_n225), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n261), .A2(KEYINPUT10), .A3(new_n262), .A4(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT66), .B(G134), .ZN(new_n266));
  INV_X1    g080(.A(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT11), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT67), .B(G131), .Z(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G137), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G134), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n274), .B1(new_n278), .B2(G137), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n270), .B(new_n272), .C1(new_n269), .C2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G131), .ZN(new_n282));
  INV_X1    g096(.A(new_n274), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n266), .B2(new_n267), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT11), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n282), .B1(new_n285), .B2(new_n270), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n234), .A2(new_n245), .A3(new_n265), .A4(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT83), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT81), .B1(new_n211), .B2(new_n226), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n229), .A2(new_n232), .A3(new_n228), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n293), .A2(new_n189), .B1(new_n238), .B2(new_n244), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n294), .A2(KEYINPUT83), .A3(new_n287), .A4(new_n265), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n250), .B1(new_n195), .B2(new_n202), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n201), .A2(new_n202), .B1(new_n297), .B2(new_n240), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n226), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n287), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n300), .A2(KEYINPUT12), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(KEYINPUT12), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(G110), .B(G140), .ZN(new_n304));
  INV_X1    g118(.A(G953), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(G227), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n304), .B(new_n306), .Z(new_n307));
  AND3_X1   g121(.A1(new_n296), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n294), .A2(new_n265), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n281), .B2(new_n286), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n296), .B2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n187), .B(new_n188), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(G469), .A2(G902), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n296), .A2(new_n303), .ZN(new_n314));
  INV_X1    g128(.A(new_n307), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n315), .B1(new_n290), .B2(new_n295), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n310), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(G469), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n312), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G221), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT9), .B(G234), .Z(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(new_n188), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G214), .B1(G237), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G478), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT15), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(G217), .A3(new_n305), .ZN(new_n330));
  INV_X1    g144(.A(G122), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G116), .ZN(new_n332));
  INV_X1    g146(.A(G116), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G122), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n332), .A2(new_n334), .A3(new_n216), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n216), .B1(new_n332), .B2(new_n334), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n200), .B1(new_n196), .B2(new_n198), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n190), .B1(new_n255), .B2(new_n257), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n338), .A2(new_n339), .A3(new_n266), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(KEYINPUT13), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT13), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT64), .B(G143), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(new_n200), .ZN(new_n344));
  INV_X1    g158(.A(new_n339), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n337), .B(new_n340), .C1(G134), .C2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT14), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n332), .A2(new_n334), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n333), .A2(KEYINPUT14), .A3(G122), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(G107), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n345), .B(new_n278), .C1(new_n200), .C2(new_n343), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n266), .B1(new_n338), .B2(new_n339), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n335), .B(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n330), .B1(new_n347), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n335), .B1(new_n353), .B2(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n351), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n337), .B1(new_n346), .B2(G134), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n353), .ZN(new_n361));
  INV_X1    g175(.A(new_n330), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n356), .A2(new_n357), .A3(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT95), .B(new_n330), .C1(new_n347), .C2(new_n355), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n188), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT96), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n329), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n367), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n364), .A2(KEYINPUT96), .A3(new_n188), .A4(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n368), .B1(new_n371), .B2(new_n329), .ZN(new_n372));
  NOR2_X1   g186(.A1(G475), .A2(G902), .ZN(new_n373));
  XNOR2_X1  g187(.A(G125), .B(G140), .ZN(new_n374));
  OR3_X1    g188(.A1(new_n374), .A2(KEYINPUT89), .A3(new_n191), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n206), .A2(new_n374), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n376), .B(KEYINPUT89), .C1(new_n191), .C2(new_n374), .ZN(new_n377));
  INV_X1    g191(.A(G237), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n378), .A2(new_n305), .A3(G214), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n380));
  AOI21_X1  g194(.A(G143), .B1(new_n380), .B2(KEYINPUT64), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(KEYINPUT18), .A2(G131), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n380), .B1(new_n196), .B2(new_n198), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n379), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n378), .A2(new_n305), .A3(G214), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n343), .B2(new_n380), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n383), .B1(new_n388), .B2(new_n382), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n375), .B(new_n377), .C1(new_n386), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT90), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n382), .ZN(new_n392));
  INV_X1    g206(.A(new_n383), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n385), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT90), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n395), .A2(new_n396), .A3(new_n375), .A4(new_n377), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n190), .B1(new_n197), .B2(KEYINPUT88), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(new_n387), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n208), .A2(KEYINPUT88), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(new_n387), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT91), .B1(new_n402), .B2(new_n271), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT17), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n392), .A2(new_n405), .A3(new_n272), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n271), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n403), .A2(new_n404), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n374), .A2(KEYINPUT16), .ZN(new_n409));
  INV_X1    g223(.A(G125), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n410), .A2(KEYINPUT16), .A3(G140), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(G146), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT16), .ZN(new_n414));
  INV_X1    g228(.A(G140), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(G125), .A2(G140), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n191), .B1(new_n418), .B2(new_n411), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n402), .A2(KEYINPUT17), .A3(new_n271), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n408), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G113), .B(G122), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT93), .B(G104), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT94), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n398), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n403), .A2(new_n407), .A3(new_n406), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n374), .B(KEYINPUT19), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(KEYINPUT92), .A3(new_n206), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT92), .ZN(new_n432));
  INV_X1    g246(.A(new_n430), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n248), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n429), .A2(new_n413), .A3(new_n431), .A4(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n426), .B1(new_n398), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n373), .B1(new_n428), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT20), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(new_n373), .C1(new_n428), .C2(new_n436), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n426), .B1(new_n398), .B2(new_n423), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n188), .B1(new_n428), .B2(new_n441), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n438), .A2(new_n440), .B1(G475), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n305), .A2(G952), .ZN(new_n444));
  INV_X1    g258(.A(G234), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(new_n378), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n188), .B(new_n305), .C1(G234), .C2(G237), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT21), .B(G898), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT97), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n372), .A2(new_n443), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n298), .A2(new_n410), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n243), .A2(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G224), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G953), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n333), .A2(KEYINPUT5), .A3(G119), .ZN(new_n461));
  XNOR2_X1  g275(.A(G116), .B(G119), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(KEYINPUT5), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT2), .B(G113), .Z(new_n464));
  AOI22_X1  g278(.A1(new_n463), .A2(G113), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n262), .A2(new_n465), .A3(new_n264), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n235), .A2(G101), .A3(new_n236), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n464), .B(new_n462), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n223), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n262), .A2(KEYINPUT84), .A3(new_n465), .A4(new_n264), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT85), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(KEYINPUT86), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n468), .A2(new_n476), .A3(new_n472), .A4(new_n473), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n460), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT6), .B1(new_n474), .B2(new_n477), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n459), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT7), .ZN(new_n483));
  OR3_X1    g297(.A1(new_n456), .A2(new_n483), .A3(new_n458), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n226), .A2(new_n465), .ZN(new_n485));
  INV_X1    g299(.A(new_n476), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n486), .A2(KEYINPUT8), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n226), .A2(new_n465), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(KEYINPUT8), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n485), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n456), .B1(new_n483), .B2(new_n458), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n479), .A2(new_n484), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n482), .A2(new_n188), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n494));
  OAI21_X1  g308(.A(G210), .B1(G237), .B2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n494), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n482), .A2(new_n188), .A3(new_n498), .A4(new_n492), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n327), .B(new_n453), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n268), .B1(G134), .B2(new_n267), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G131), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n280), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n253), .B2(new_n260), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n278), .A2(G137), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n269), .B1(new_n506), .B2(new_n283), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT11), .B1(new_n266), .B2(new_n267), .ZN(new_n508));
  OAI21_X1  g322(.A(G131), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n243), .B1(new_n509), .B2(new_n280), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n505), .A2(new_n470), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n470), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n508), .B1(KEYINPUT11), .B2(new_n284), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n513), .A2(new_n272), .B1(G131), .B2(new_n502), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n259), .A2(KEYINPUT69), .A3(new_n231), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT69), .B1(new_n259), .B2(new_n231), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n244), .B1(new_n281), .B2(new_n286), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n501), .B(KEYINPUT28), .C1(new_n511), .C2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT28), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n470), .B1(new_n505), .B2(new_n510), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n512), .A3(new_n518), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT71), .B1(new_n523), .B2(new_n521), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n378), .A2(new_n305), .A3(G210), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n221), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n528), .B(new_n529), .Z(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT29), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n188), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(KEYINPUT72), .B(new_n188), .C1(new_n526), .C2(new_n531), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n517), .A2(KEYINPUT30), .A3(new_n518), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n504), .A2(new_n298), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(new_n510), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n470), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT70), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n536), .A2(new_n539), .A3(KEYINPUT70), .A4(new_n470), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n523), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n530), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n523), .A2(new_n521), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n470), .B1(new_n538), .B2(new_n510), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n517), .A2(KEYINPUT28), .A3(new_n512), .A4(new_n518), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n551), .A2(new_n545), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n534), .A2(new_n535), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G472), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT32), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n542), .A2(new_n523), .A3(new_n530), .A4(new_n543), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n557), .A2(KEYINPUT31), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(KEYINPUT31), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n551), .A2(new_n545), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(G472), .A2(G902), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n556), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n557), .A2(KEYINPUT31), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n560), .B1(new_n557), .B2(KEYINPUT31), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n556), .B(new_n562), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n555), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT22), .B(G137), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n321), .A2(new_n445), .A3(G953), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n569), .B(new_n570), .Z(new_n571));
  INV_X1    g385(.A(KEYINPUT76), .ZN(new_n572));
  AOI21_X1  g386(.A(G146), .B1(new_n409), .B2(new_n412), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n418), .A2(new_n191), .A3(new_n411), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT24), .B(G110), .ZN(new_n575));
  OR3_X1    g389(.A1(new_n200), .A2(KEYINPUT73), .A3(G119), .ZN(new_n576));
  INV_X1    g390(.A(G119), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G128), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT73), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n576), .B(new_n579), .C1(new_n250), .C2(new_n577), .ZN(new_n580));
  OAI22_X1  g394(.A1(new_n573), .A2(new_n574), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G110), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n577), .B1(new_n255), .B2(new_n257), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n583), .A2(KEYINPUT23), .B1(new_n577), .B2(G128), .ZN(new_n584));
  OR2_X1    g398(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n585));
  NAND2_X1  g399(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n585), .B(new_n586), .C1(new_n577), .C2(G128), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n582), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT75), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(KEYINPUT23), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n587), .A3(new_n578), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G110), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT75), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n580), .A2(new_n575), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n420), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n413), .A2(new_n376), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n584), .A2(new_n582), .A3(new_n587), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n580), .A2(new_n575), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n572), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  AOI211_X1 g416(.A(KEYINPUT76), .B(new_n600), .C1(new_n589), .C2(new_n595), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n571), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT79), .ZN(new_n605));
  INV_X1    g419(.A(new_n571), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n596), .A2(new_n601), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(KEYINPUT76), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n605), .B1(new_n604), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g424(.A(G217), .B1(new_n445), .B2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n188), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n604), .A2(new_n188), .A3(new_n608), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT78), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT77), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g431(.A(KEYINPUT25), .B(new_n615), .C1(new_n617), .C2(KEYINPUT78), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT78), .B1(new_n614), .B2(new_n616), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT25), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n611), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n613), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n325), .A2(new_n500), .A3(new_n568), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  AND3_X1   g438(.A1(new_n320), .A2(new_n622), .A3(new_n324), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n561), .A2(new_n188), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n626), .A2(G472), .B1(new_n562), .B2(new_n561), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n493), .A2(new_n495), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n482), .A2(new_n188), .A3(new_n496), .A4(new_n492), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n630), .A2(new_n326), .A3(new_n452), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n438), .A2(new_n440), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n442), .A2(G475), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n364), .A2(new_n636), .A3(new_n365), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n356), .A2(KEYINPUT33), .A3(new_n363), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(G478), .A3(new_n188), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n366), .A2(new_n328), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n632), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n629), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NAND2_X1  g460(.A1(new_n440), .A2(KEYINPUT98), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n438), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n437), .A2(KEYINPUT98), .A3(KEYINPUT20), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n648), .A2(new_n649), .B1(G475), .B2(new_n442), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n371), .A2(new_n329), .ZN(new_n651));
  INV_X1    g465(.A(new_n368), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n632), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n629), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  INV_X1    g472(.A(new_n612), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n607), .B(KEYINPUT99), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n606), .A2(KEYINPUT36), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n660), .B(new_n661), .Z(new_n662));
  AOI22_X1  g476(.A1(new_n618), .A2(new_n621), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n325), .A2(new_n500), .A3(new_n627), .A4(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  AND3_X1   g481(.A1(new_n630), .A2(new_n326), .A3(new_n631), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n648), .A2(new_n649), .ZN(new_n669));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n447), .B1(new_n448), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n669), .A2(new_n653), .A3(new_n634), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n650), .A2(new_n675), .A3(new_n653), .A4(new_n672), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n668), .A2(new_n674), .A3(KEYINPUT101), .A4(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n677), .A2(new_n568), .A3(new_n664), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n320), .A2(new_n324), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n668), .A2(new_n674), .A3(new_n676), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  NOR2_X1   g498(.A1(new_n563), .A2(new_n567), .ZN(new_n685));
  INV_X1    g499(.A(G472), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n544), .A2(new_n530), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n511), .A2(new_n519), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n689), .B2(new_n545), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n686), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n671), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n325), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n664), .B(new_n692), .C1(new_n696), .C2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n372), .A2(new_n443), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n497), .A2(new_n499), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT102), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT38), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n699), .A2(new_n326), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n343), .ZN(G45));
  OAI21_X1  g519(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT32), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n707), .A2(new_n566), .B1(G472), .B2(new_n554), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n630), .A2(new_n326), .A3(new_n631), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n443), .B1(new_n640), .B2(new_n639), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n672), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n708), .A2(new_n709), .A3(new_n663), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n325), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT103), .B(G146), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G48));
  NAND2_X1  g529(.A1(KEYINPUT104), .A2(G469), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n296), .A2(new_n310), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n718), .A2(new_n315), .B1(new_n317), .B2(new_n303), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n717), .B1(new_n719), .B2(G902), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n188), .B(new_n716), .C1(new_n308), .C2(new_n311), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n720), .A2(new_n324), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n568), .A2(new_n643), .A3(new_n722), .A4(new_n622), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND4_X1  g539(.A1(new_n568), .A2(new_n655), .A3(new_n722), .A4(new_n622), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NAND4_X1  g541(.A1(new_n568), .A2(new_n722), .A3(new_n668), .A4(new_n664), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n453), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n577), .ZN(G21));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n626), .A2(G472), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n557), .A2(KEYINPUT31), .ZN(new_n734));
  AOI22_X1  g548(.A1(KEYINPUT31), .A2(new_n557), .B1(new_n526), .B2(new_n545), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n526), .A2(new_n545), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n559), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT105), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n733), .B1(new_n741), .B2(new_n562), .ZN(new_n742));
  INV_X1    g556(.A(new_n562), .ZN(new_n743));
  AOI211_X1 g557(.A(KEYINPUT106), .B(new_n743), .C1(new_n737), .C2(new_n740), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n622), .B(new_n732), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n722), .A2(new_n452), .A3(new_n668), .A4(new_n700), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n731), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n732), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n558), .B1(new_n739), .B2(KEYINPUT105), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n735), .A2(new_n736), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n562), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT106), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n741), .A2(new_n733), .A3(new_n562), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n720), .A2(new_n324), .A3(new_n721), .ZN(new_n755));
  NOR4_X1   g569(.A1(new_n755), .A2(new_n632), .A3(new_n372), .A4(new_n443), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n754), .A2(new_n756), .A3(KEYINPUT107), .A4(new_n622), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  OAI211_X1 g573(.A(new_n732), .B(new_n664), .C1(new_n742), .C2(new_n744), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n722), .A2(new_n710), .A3(new_n668), .A4(new_n672), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT108), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n755), .A2(new_n709), .A3(new_n711), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n754), .A2(new_n763), .A3(new_n664), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT109), .B(G125), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G27));
  INV_X1    g582(.A(new_n622), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n708), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n701), .A2(new_n711), .A3(new_n327), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n325), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n770), .A2(KEYINPUT42), .A3(new_n325), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  AOI21_X1  g591(.A(KEYINPUT110), .B1(new_n674), .B2(new_n676), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n778), .A2(new_n708), .A3(new_n679), .A4(new_n769), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n674), .A2(KEYINPUT110), .A3(new_n676), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n701), .A2(new_n327), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  AOI22_X1  g598(.A1(new_n314), .A2(new_n315), .B1(new_n317), .B2(new_n310), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT45), .Z(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(G469), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n313), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n312), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT111), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n791), .A3(new_n312), .ZN(new_n792));
  OAI21_X1  g606(.A(G469), .B1(new_n786), .B2(G902), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n790), .B(new_n792), .C1(KEYINPUT46), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n324), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n627), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT43), .B1(new_n443), .B2(KEYINPUT112), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n443), .A2(new_n641), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n800), .A3(new_n664), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n796), .A2(new_n693), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n781), .B1(new_n801), .B2(new_n802), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n267), .ZN(G39));
  NAND3_X1  g621(.A1(new_n771), .A2(new_n769), .A3(new_n708), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT113), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n794), .A2(KEYINPUT47), .A3(new_n324), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT47), .B1(new_n794), .B2(new_n324), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(KEYINPUT114), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  NOR2_X1   g631(.A1(new_n703), .A2(new_n769), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n799), .A2(new_n327), .A3(new_n323), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n720), .A2(new_n721), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT49), .Z(new_n821));
  NAND4_X1  g635(.A1(new_n818), .A2(new_n692), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n810), .A2(new_n811), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n324), .B2(new_n820), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n447), .A2(new_n754), .A3(new_n622), .A4(new_n800), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n781), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n722), .A2(new_n327), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n703), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n829), .B(new_n825), .C1(new_n827), .C2(new_n828), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT50), .Z(new_n831));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n832));
  INV_X1    g646(.A(new_n781), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n446), .A3(new_n755), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n834), .A2(new_n622), .A3(new_n692), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n635), .A2(new_n641), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n834), .A2(new_n800), .ZN(new_n837));
  INV_X1    g651(.A(new_n760), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n832), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n826), .A2(new_n831), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n826), .A2(new_n839), .A3(new_n831), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(KEYINPUT51), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n678), .A2(new_n682), .B1(new_n712), .B2(new_n325), .ZN(new_n846));
  INV_X1    g660(.A(new_n692), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n664), .A2(new_n671), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n709), .A2(new_n372), .A3(new_n443), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n847), .A2(new_n325), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n766), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n766), .A2(new_n846), .A3(KEYINPUT52), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n642), .B1(new_n372), .B2(new_n635), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n326), .A2(new_n701), .A3(new_n856), .A4(new_n452), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n625), .A3(new_n627), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n623), .A3(new_n665), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT115), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n858), .A2(new_n623), .A3(new_n665), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n723), .B(new_n726), .C1(new_n728), .C2(new_n453), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n747), .B2(new_n757), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n774), .A2(new_n775), .B1(new_n782), .B2(new_n779), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n568), .A2(new_n372), .A3(new_n650), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n732), .B1(new_n742), .B2(new_n744), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n868), .B2(new_n642), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n833), .A2(new_n663), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n325), .A3(new_n672), .A4(new_n870), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n863), .A2(new_n865), .A3(new_n866), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n855), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n855), .A2(new_n872), .A3(KEYINPUT53), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT54), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n837), .A2(new_n770), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT48), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n835), .A2(new_n710), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n825), .A2(new_n668), .A3(new_n722), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n880), .A2(new_n444), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT118), .Z(new_n884));
  NOR3_X1   g698(.A1(new_n845), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(G952), .A2(G953), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n822), .B1(new_n885), .B2(new_n886), .ZN(G75));
  OR2_X1    g701(.A1(new_n480), .A2(new_n481), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(new_n459), .Z(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT119), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT55), .Z(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n188), .B1(new_n875), .B2(new_n876), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n893), .B2(G210), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n305), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(G51));
  INV_X1    g716(.A(new_n878), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n313), .B(KEYINPUT57), .ZN(new_n904));
  OAI22_X1  g718(.A1(new_n903), .A2(new_n904), .B1(new_n311), .B2(new_n308), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n893), .A2(G469), .A3(new_n786), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT121), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n900), .B1(new_n905), .B2(new_n907), .ZN(G54));
  NAND3_X1  g722(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n428), .A2(new_n436), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n900), .ZN(G60));
  XNOR2_X1  g726(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n328), .A2(new_n188), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n878), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n637), .A2(new_n638), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n900), .ZN(G63));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT123), .Z(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT60), .Z(new_n923));
  AND3_X1   g737(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n872), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT53), .B1(new_n855), .B2(new_n872), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n609), .A2(new_n610), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n900), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n662), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n928), .A2(KEYINPUT61), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n931));
  INV_X1    g745(.A(new_n929), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n928), .B2(KEYINPUT124), .ZN(new_n933));
  INV_X1    g747(.A(new_n923), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n875), .B2(new_n876), .ZN(new_n935));
  INV_X1    g749(.A(new_n927), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n901), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n931), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI211_X1 g756(.A(KEYINPUT125), .B(KEYINPUT61), .C1(new_n933), .C2(new_n939), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n930), .B1(new_n942), .B2(new_n943), .ZN(G66));
  OAI21_X1  g758(.A(G953), .B1(new_n450), .B2(new_n457), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n863), .A2(new_n865), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(G953), .ZN(new_n947));
  INV_X1    g761(.A(G898), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n888), .B1(new_n948), .B2(G953), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n947), .B(new_n949), .Z(G69));
  NAND2_X1  g764(.A1(G227), .A2(G900), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n670), .A2(G953), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT127), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n806), .B1(new_n814), .B2(new_n815), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n796), .A2(new_n770), .A3(new_n693), .A4(new_n849), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n766), .A2(new_n846), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n866), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n954), .B1(new_n959), .B2(new_n305), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n536), .A2(new_n539), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n430), .ZN(new_n963));
  OAI211_X1 g777(.A(G953), .B(new_n951), .C1(new_n961), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n704), .A2(new_n957), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n856), .A2(KEYINPUT126), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n695), .A2(new_n770), .A3(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n969), .B(new_n781), .C1(KEYINPUT126), .C2(new_n856), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n955), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n963), .B1(new_n971), .B2(G953), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n951), .A2(G953), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n972), .B(new_n973), .C1(new_n960), .C2(new_n963), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n964), .A2(new_n974), .ZN(G72));
  NAND4_X1  g789(.A1(new_n955), .A2(new_n946), .A3(new_n866), .A4(new_n958), .ZN(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  AOI211_X1 g792(.A(new_n530), .B(new_n544), .C1(new_n976), .C2(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n955), .A2(new_n946), .A3(new_n967), .A4(new_n970), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n688), .B1(new_n980), .B2(new_n978), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n546), .A2(new_n557), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n877), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NOR4_X1   g798(.A1(new_n979), .A2(new_n900), .A3(new_n981), .A4(new_n984), .ZN(G57));
endmodule


