

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  XNOR2_X1 U324 ( .A(n581), .B(n402), .ZN(n464) );
  XNOR2_X1 U325 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U326 ( .A(n299), .B(n292), .ZN(n300) );
  INV_X1 U327 ( .A(n369), .ZN(n310) );
  XNOR2_X1 U328 ( .A(n321), .B(n320), .ZN(n322) );
  AND2_X1 U329 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U330 ( .A(n413), .B(KEYINPUT120), .Z(n293) );
  XOR2_X1 U331 ( .A(G43GAT), .B(G99GAT), .Z(n294) );
  INV_X1 U332 ( .A(KEYINPUT74), .ZN(n382) );
  INV_X1 U333 ( .A(KEYINPUT54), .ZN(n413) );
  XNOR2_X1 U334 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U335 ( .A(n373), .B(n319), .ZN(n320) );
  XNOR2_X1 U336 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U337 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U338 ( .A(n351), .B(n294), .ZN(n324) );
  XNOR2_X1 U339 ( .A(n396), .B(n395), .ZN(n399) );
  XNOR2_X1 U340 ( .A(n312), .B(n311), .ZN(n407) );
  XNOR2_X1 U341 ( .A(n325), .B(n324), .ZN(n326) );
  NOR2_X1 U342 ( .A1(n522), .A2(n514), .ZN(n519) );
  XNOR2_X1 U343 ( .A(KEYINPUT38), .B(n491), .ZN(n511) );
  XNOR2_X1 U344 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n492) );
  XNOR2_X1 U346 ( .A(n468), .B(n467), .ZN(G1349GAT) );
  XNOR2_X1 U347 ( .A(n493), .B(n492), .ZN(G1330GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n296) );
  XOR2_X1 U349 ( .A(G190GAT), .B(G134GAT), .Z(n317) );
  XOR2_X1 U350 ( .A(G218GAT), .B(G162GAT), .Z(n451) );
  XNOR2_X1 U351 ( .A(n317), .B(n451), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n301) );
  XOR2_X1 U353 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n298) );
  XNOR2_X1 U354 ( .A(KEYINPUT66), .B(KEYINPUT79), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U356 ( .A(n302), .B(KEYINPUT9), .Z(n312) );
  XOR2_X1 U357 ( .A(G29GAT), .B(KEYINPUT8), .Z(n304) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(G36GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U360 ( .A(G50GAT), .B(KEYINPUT7), .Z(n305) );
  XOR2_X1 U361 ( .A(n306), .B(n305), .Z(n369) );
  XOR2_X1 U362 ( .A(G92GAT), .B(G85GAT), .Z(n308) );
  XNOR2_X1 U363 ( .A(G99GAT), .B(G106GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n385) );
  XNOR2_X1 U365 ( .A(KEYINPUT82), .B(n385), .ZN(n309) );
  XOR2_X1 U366 ( .A(KEYINPUT83), .B(n407), .Z(n546) );
  XOR2_X1 U367 ( .A(G176GAT), .B(KEYINPUT20), .Z(n314) );
  XNOR2_X1 U368 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n327) );
  XOR2_X1 U370 ( .A(G183GAT), .B(KEYINPUT17), .Z(n316) );
  XNOR2_X1 U371 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n333) );
  XOR2_X1 U373 ( .A(n333), .B(n317), .Z(n323) );
  XNOR2_X1 U374 ( .A(G120GAT), .B(KEYINPUT0), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n318), .B(KEYINPUT91), .ZN(n431) );
  XOR2_X1 U376 ( .A(n431), .B(G71GAT), .Z(n321) );
  XOR2_X1 U377 ( .A(G169GAT), .B(G113GAT), .Z(n373) );
  NAND2_X1 U378 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n325) );
  XOR2_X1 U380 ( .A(G15GAT), .B(G127GAT), .Z(n351) );
  XOR2_X2 U381 ( .A(n327), .B(n326), .Z(n534) );
  INV_X1 U382 ( .A(n534), .ZN(n471) );
  XOR2_X1 U383 ( .A(G204GAT), .B(G36GAT), .Z(n329) );
  NAND2_X1 U384 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n332) );
  XOR2_X1 U386 ( .A(KEYINPUT21), .B(KEYINPUT96), .Z(n331) );
  XNOR2_X1 U387 ( .A(G197GAT), .B(KEYINPUT95), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n440) );
  XOR2_X1 U389 ( .A(n332), .B(n440), .Z(n335) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(n333), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U392 ( .A(KEYINPUT82), .B(G92GAT), .Z(n337) );
  XNOR2_X1 U393 ( .A(G190GAT), .B(G218GAT), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U395 ( .A(n339), .B(n338), .Z(n341) );
  XOR2_X1 U396 ( .A(G8GAT), .B(G211GAT), .Z(n354) );
  XOR2_X1 U397 ( .A(G176GAT), .B(G64GAT), .Z(n388) );
  XNOR2_X1 U398 ( .A(n354), .B(n388), .ZN(n340) );
  XOR2_X1 U399 ( .A(n341), .B(n340), .Z(n526) );
  INV_X1 U400 ( .A(n526), .ZN(n472) );
  XOR2_X1 U401 ( .A(KEYINPUT89), .B(KEYINPUT87), .Z(n343) );
  XNOR2_X1 U402 ( .A(KEYINPUT15), .B(KEYINPUT84), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U404 ( .A(KEYINPUT86), .B(KEYINPUT14), .Z(n345) );
  XNOR2_X1 U405 ( .A(KEYINPUT88), .B(KEYINPUT12), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U407 ( .A(n347), .B(n346), .Z(n353) );
  XOR2_X1 U408 ( .A(KEYINPUT85), .B(KEYINPUT90), .Z(n349) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U413 ( .A(G64GAT), .B(n354), .Z(n356) );
  XOR2_X1 U414 ( .A(G22GAT), .B(G155GAT), .Z(n443) );
  XNOR2_X1 U415 ( .A(G183GAT), .B(n443), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U417 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U418 ( .A(G1GAT), .B(KEYINPUT70), .Z(n372) );
  XOR2_X1 U419 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n360) );
  XNOR2_X1 U420 ( .A(G71GAT), .B(G78GAT), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U422 ( .A(G57GAT), .B(n361), .ZN(n397) );
  XOR2_X1 U423 ( .A(n372), .B(n397), .Z(n362) );
  XOR2_X1 U424 ( .A(n363), .B(n362), .Z(n561) );
  INV_X1 U425 ( .A(n561), .ZN(n584) );
  XNOR2_X1 U426 ( .A(KEYINPUT36), .B(n546), .ZN(n469) );
  NOR2_X1 U427 ( .A1(n584), .A2(n469), .ZN(n365) );
  XNOR2_X1 U428 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n401) );
  XOR2_X1 U430 ( .A(KEYINPUT30), .B(G8GAT), .Z(n367) );
  XNOR2_X1 U431 ( .A(G22GAT), .B(G141GAT), .ZN(n366) );
  XNOR2_X1 U432 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n381) );
  XOR2_X1 U434 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n371) );
  XNOR2_X1 U435 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n377) );
  XOR2_X1 U437 ( .A(G197GAT), .B(G15GAT), .Z(n375) );
  XNOR2_X1 U438 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U440 ( .A(n377), .B(n376), .Z(n379) );
  NAND2_X1 U441 ( .A1(G229GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U443 ( .A(n381), .B(n380), .Z(n576) );
  INV_X1 U444 ( .A(n576), .ZN(n554) );
  XOR2_X1 U445 ( .A(KEYINPUT72), .B(n554), .Z(n490) );
  NAND2_X1 U446 ( .A1(G230GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U447 ( .A(G120GAT), .B(n386), .ZN(n396) );
  XOR2_X1 U448 ( .A(G204GAT), .B(G148GAT), .Z(n444) );
  XOR2_X1 U449 ( .A(KEYINPUT31), .B(KEYINPUT77), .Z(n387) );
  XNOR2_X1 U450 ( .A(n444), .B(n387), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U452 ( .A(n390), .B(KEYINPUT76), .Z(n394) );
  XOR2_X1 U453 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n392) );
  XNOR2_X1 U454 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  INV_X1 U457 ( .A(n397), .ZN(n398) );
  XOR2_X2 U458 ( .A(n399), .B(n398), .Z(n581) );
  NAND2_X1 U459 ( .A1(n490), .A2(n581), .ZN(n400) );
  NOR2_X1 U460 ( .A1(n401), .A2(n400), .ZN(n411) );
  XNOR2_X1 U461 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n402) );
  NAND2_X1 U462 ( .A1(n464), .A2(n554), .ZN(n404) );
  XNOR2_X1 U463 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n561), .B(KEYINPUT111), .ZN(n569) );
  NAND2_X1 U466 ( .A1(n405), .A2(n569), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n406), .B(KEYINPUT113), .ZN(n408) );
  NAND2_X1 U468 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U469 ( .A(KEYINPUT47), .B(n409), .ZN(n410) );
  NOR2_X1 U470 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n412), .B(KEYINPUT48), .ZN(n551) );
  NOR2_X1 U472 ( .A1(n472), .A2(n551), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n414), .B(n293), .ZN(n573) );
  XOR2_X1 U474 ( .A(KEYINPUT4), .B(KEYINPUT100), .Z(n416) );
  XNOR2_X1 U475 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n435) );
  XOR2_X1 U477 ( .A(G134GAT), .B(G127GAT), .Z(n418) );
  XNOR2_X1 U478 ( .A(G29GAT), .B(G113GAT), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U480 ( .A(KEYINPUT101), .B(KEYINPUT5), .Z(n420) );
  XNOR2_X1 U481 ( .A(G148GAT), .B(G155GAT), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U483 ( .A(n422), .B(n421), .Z(n429) );
  XOR2_X1 U484 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n424) );
  XNOR2_X1 U485 ( .A(G141GAT), .B(KEYINPUT97), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n439) );
  XOR2_X1 U487 ( .A(G85GAT), .B(G162GAT), .Z(n426) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n439), .B(n427), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U492 ( .A(n430), .B(G57GAT), .Z(n433) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(n435), .B(n434), .Z(n572) );
  XOR2_X1 U496 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n437) );
  NAND2_X1 U497 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U499 ( .A(n438), .B(G211GAT), .Z(n442) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n448) );
  XOR2_X1 U502 ( .A(G106GAT), .B(n443), .Z(n446) );
  XNOR2_X1 U503 ( .A(G50GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U505 ( .A(n448), .B(n447), .Z(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT22), .B(KEYINPUT99), .Z(n450) );
  XNOR2_X1 U507 ( .A(G78GAT), .B(KEYINPUT98), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n480) );
  AND2_X1 U511 ( .A1(n572), .A2(n480), .ZN(n455) );
  NAND2_X1 U512 ( .A1(n573), .A2(n455), .ZN(n457) );
  XOR2_X1 U513 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n456) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U515 ( .A(n458), .B(KEYINPUT122), .Z(n459) );
  NOR2_X2 U516 ( .A1(n471), .A2(n459), .ZN(n566) );
  INV_X1 U517 ( .A(n566), .ZN(n570) );
  NOR2_X1 U518 ( .A1(n546), .A2(n570), .ZN(n463) );
  XNOR2_X1 U519 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n461) );
  INV_X1 U520 ( .A(G190GAT), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XNOR2_X1 U522 ( .A(KEYINPUT110), .B(n464), .ZN(n537) );
  NAND2_X1 U523 ( .A1(n537), .A2(n566), .ZN(n468) );
  XOR2_X1 U524 ( .A(G176GAT), .B(KEYINPUT57), .Z(n466) );
  XOR2_X1 U525 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n465) );
  XNOR2_X1 U526 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n526), .B(KEYINPUT27), .ZN(n482) );
  NOR2_X1 U528 ( .A1(n534), .A2(n480), .ZN(n470) );
  XNOR2_X1 U529 ( .A(KEYINPUT26), .B(n470), .ZN(n574) );
  NAND2_X1 U530 ( .A1(n482), .A2(n574), .ZN(n478) );
  NOR2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U532 ( .A(KEYINPUT103), .B(n473), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n474), .A2(n480), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT104), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT25), .B(n476), .Z(n477) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n479), .A2(n572), .ZN(n486) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT67), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n481), .B(KEYINPUT28), .ZN(n529) );
  INV_X1 U540 ( .A(n572), .ZN(n524) );
  NAND2_X1 U541 ( .A1(n482), .A2(n524), .ZN(n550) );
  NOR2_X1 U542 ( .A1(n529), .A2(n550), .ZN(n533) );
  XNOR2_X1 U543 ( .A(KEYINPUT102), .B(n533), .ZN(n484) );
  XOR2_X1 U544 ( .A(n534), .B(KEYINPUT94), .Z(n483) );
  NAND2_X1 U545 ( .A1(n484), .A2(n483), .ZN(n485) );
  NAND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n497) );
  NAND2_X1 U547 ( .A1(n584), .A2(n497), .ZN(n487) );
  XOR2_X1 U548 ( .A(KEYINPUT107), .B(n487), .Z(n488) );
  NOR2_X1 U549 ( .A1(n469), .A2(n488), .ZN(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT37), .B(n489), .ZN(n523) );
  INV_X1 U551 ( .A(n490), .ZN(n567) );
  NAND2_X1 U552 ( .A1(n567), .A2(n581), .ZN(n499) );
  NOR2_X1 U553 ( .A1(n523), .A2(n499), .ZN(n491) );
  NAND2_X1 U554 ( .A1(n511), .A2(n534), .ZN(n493) );
  NAND2_X1 U555 ( .A1(n511), .A2(n526), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(KEYINPUT108), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n546), .A2(n561), .ZN(n496) );
  XOR2_X1 U559 ( .A(KEYINPUT16), .B(n496), .Z(n498) );
  NAND2_X1 U560 ( .A1(n498), .A2(n497), .ZN(n514) );
  NOR2_X1 U561 ( .A1(n499), .A2(n514), .ZN(n507) );
  NAND2_X1 U562 ( .A1(n524), .A2(n507), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U565 ( .A1(n526), .A2(n507), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT106), .B(KEYINPUT35), .Z(n504) );
  NAND2_X1 U568 ( .A1(n507), .A2(n534), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n506) );
  XOR2_X1 U570 ( .A(G15GAT), .B(KEYINPUT105), .Z(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1326GAT) );
  NAND2_X1 U572 ( .A1(n507), .A2(n529), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U574 ( .A(G29GAT), .B(KEYINPUT39), .Z(n510) );
  NAND2_X1 U575 ( .A1(n511), .A2(n524), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  XOR2_X1 U577 ( .A(G50GAT), .B(KEYINPUT109), .Z(n513) );
  NAND2_X1 U578 ( .A1(n529), .A2(n511), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1331GAT) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n516) );
  NAND2_X1 U581 ( .A1(n537), .A2(n576), .ZN(n522) );
  NAND2_X1 U582 ( .A1(n519), .A2(n524), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1332GAT) );
  NAND2_X1 U584 ( .A1(n526), .A2(n519), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n517), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n534), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n518), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U589 ( .A1(n519), .A2(n529), .ZN(n520) );
  XNOR2_X1 U590 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NOR2_X1 U591 ( .A1(n523), .A2(n522), .ZN(n530) );
  NAND2_X1 U592 ( .A1(n530), .A2(n524), .ZN(n525) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n526), .A2(n530), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n527), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n530), .A2(n534), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n551), .A2(n535), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n567), .A2(n541), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n539) );
  NAND2_X1 U606 ( .A1(n541), .A2(n537), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  INV_X1 U609 ( .A(n541), .ZN(n545) );
  NOR2_X1 U610 ( .A1(n569), .A2(n545), .ZN(n543) );
  XNOR2_X1 U611 ( .A(KEYINPUT115), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  NOR2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U619 ( .A1(n574), .A2(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT117), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n563), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U626 ( .A(KEYINPUT118), .B(n558), .Z(n560) );
  NAND2_X1 U627 ( .A1(n563), .A2(n464), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n562), .ZN(G1346GAT) );
  INV_X1 U631 ( .A(n407), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(G183GAT), .B(n571), .Z(G1350GAT) );
  AND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n587) );
  NOR2_X1 U640 ( .A1(n587), .A2(n576), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n578) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n587), .ZN(n583) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n587), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n469), .A2(n587), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

