//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT75), .Z(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT81), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(KEYINPUT25), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n195), .B(KEYINPUT80), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT22), .B(G137), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(G128), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G119), .B(G128), .ZN(new_n207));
  INV_X1    g021(.A(G110), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT24), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G110), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n206), .A2(G110), .B1(new_n207), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G125), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n214), .A2(KEYINPUT16), .A3(G140), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G140), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G125), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(G140), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT16), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n216), .A2(new_n220), .A3(G146), .ZN(new_n221));
  AOI21_X1  g035(.A(G146), .B1(new_n216), .B2(new_n220), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n213), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n213), .B(KEYINPUT76), .C1(new_n221), .C2(new_n222), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n204), .A2(G119), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n203), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT24), .B(G110), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n202), .A2(new_n205), .A3(new_n208), .A4(new_n203), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n230), .A2(KEYINPUT77), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT77), .B1(new_n230), .B2(new_n231), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G125), .B(G140), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n215), .B1(new_n235), .B2(KEYINPUT16), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n218), .A2(new_n219), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT78), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT78), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G146), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT79), .B1(new_n234), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n230), .A2(new_n231), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT77), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT79), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n240), .B1(new_n218), .B2(new_n219), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n253), .A2(new_n241), .B1(new_n236), .B2(G146), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  AOI221_X4 g069(.A(new_n199), .B1(new_n225), .B2(new_n226), .C1(new_n245), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n245), .A2(new_n255), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n225), .A2(new_n226), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n198), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G902), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n193), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n234), .A2(KEYINPUT79), .A3(new_n244), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n251), .B1(new_n250), .B2(new_n254), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n199), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n257), .A2(new_n258), .A3(new_n198), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n261), .A3(new_n267), .A4(new_n193), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n190), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n261), .A3(new_n267), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n192), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n268), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT82), .A3(new_n190), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n188), .A2(new_n261), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n260), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n272), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT83), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n282));
  OR2_X1    g096(.A1(KEYINPUT70), .A2(KEYINPUT27), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT70), .A2(KEYINPUT27), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(KEYINPUT71), .A3(new_n284), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(G237), .A2(G953), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G210), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT26), .B(G101), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n287), .A2(new_n291), .A3(new_n288), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n294), .B1(new_n293), .B2(new_n295), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n300));
  XNOR2_X1  g114(.A(G143), .B(G146), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT0), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n204), .A3(KEYINPUT64), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT64), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(KEYINPUT0), .B2(G128), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT0), .A2(G128), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n301), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n301), .A2(new_n307), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n300), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT11), .ZN(new_n312));
  INV_X1    g126(.A(G134), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n312), .B1(new_n313), .B2(G137), .ZN(new_n314));
  INV_X1    g128(.A(G137), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT11), .A3(G134), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(G137), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G131), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT66), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n320), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n322), .A2(new_n314), .A3(new_n316), .A4(new_n317), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n303), .A2(new_n305), .B1(KEYINPUT0), .B2(G128), .ZN(new_n325));
  OAI211_X1 g139(.A(KEYINPUT65), .B(new_n309), .C1(new_n325), .C2(new_n301), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n311), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n301), .ZN(new_n328));
  INV_X1    g142(.A(G143), .ZN(new_n329));
  OAI211_X1 g143(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n329), .C2(G146), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n242), .A2(G143), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT67), .B1(new_n332), .B2(KEYINPUT1), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n328), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(G146), .ZN(new_n336));
  AND4_X1   g150(.A1(new_n335), .A2(new_n332), .A3(new_n336), .A4(G128), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n318), .A2(new_n319), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n315), .A2(G134), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n317), .A3(G131), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n327), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G116), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G119), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT68), .B1(new_n201), .B2(G116), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n346), .A3(G119), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT2), .B(G113), .Z(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n345), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n309), .B1(new_n325), .B2(new_n301), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n339), .A2(new_n343), .B1(new_n324), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n353), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n299), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n324), .A2(new_n355), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT1), .B1(new_n329), .B2(G146), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT67), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(G128), .A3(new_n330), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n337), .B1(new_n364), .B2(new_n328), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n340), .A2(new_n342), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n360), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n353), .B1(new_n367), .B2(KEYINPUT73), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n356), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT28), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n298), .B1(new_n359), .B2(new_n371), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n296), .A2(new_n297), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT69), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n356), .A2(new_n374), .A3(KEYINPUT30), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n374), .B1(new_n356), .B2(KEYINPUT30), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n355), .A2(new_n300), .B1(new_n321), .B2(new_n323), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n378), .A2(new_n326), .B1(new_n339), .B2(new_n343), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n353), .B1(new_n379), .B2(KEYINPUT30), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n358), .B(new_n373), .C1(new_n377), .C2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n372), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n357), .B1(new_n356), .B2(new_n369), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n367), .A2(KEYINPUT73), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n299), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n356), .B(new_n353), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(new_n299), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n298), .A2(KEYINPUT29), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n261), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G472), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n373), .B1(new_n359), .B2(new_n371), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT31), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n298), .A2(new_n358), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n392), .B(new_n394), .C1(new_n377), .C2(new_n380), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n344), .A2(KEYINPUT30), .A3(new_n360), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT69), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n356), .A2(new_n374), .A3(KEYINPUT30), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT30), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n357), .B1(new_n345), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n393), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT72), .B1(new_n403), .B2(new_n392), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n394), .B1(new_n377), .B2(new_n380), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT72), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT31), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n396), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(G472), .A2(G902), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT32), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n390), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n367), .A2(new_n353), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n357), .B1(new_n327), .B2(new_n344), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT28), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n385), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n373), .A2(new_n415), .B1(new_n403), .B2(new_n392), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n406), .B1(new_n405), .B2(KEYINPUT31), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n403), .A2(KEYINPUT72), .A3(new_n392), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT32), .B1(new_n419), .B2(new_n409), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n282), .B1(new_n411), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n422));
  INV_X1    g236(.A(new_n409), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n422), .B1(new_n408), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(KEYINPUT32), .A3(new_n409), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(KEYINPUT74), .A3(new_n425), .A4(new_n390), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n272), .A2(new_n427), .A3(new_n276), .A4(new_n279), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n281), .A2(new_n421), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT9), .B(G234), .ZN(new_n430));
  OAI21_X1  g244(.A(G221), .B1(new_n430), .B2(G902), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n432));
  INV_X1    g246(.A(G237), .ZN(new_n433));
  AND4_X1   g247(.A1(G143), .A2(new_n433), .A3(new_n194), .A4(G214), .ZN(new_n434));
  AOI21_X1  g248(.A(G143), .B1(new_n290), .B2(G214), .ZN(new_n435));
  OAI21_X1  g249(.A(G131), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT17), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n194), .A3(G214), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n329), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n290), .A2(G143), .A3(G214), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n319), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT95), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n221), .A2(new_n222), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT95), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n436), .A2(new_n441), .A3(new_n445), .A4(new_n437), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n436), .A2(new_n437), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n443), .A2(new_n444), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n439), .A2(KEYINPUT92), .A3(new_n440), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT18), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n449), .B1(new_n450), .B2(new_n319), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n319), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n439), .A2(KEYINPUT92), .A3(new_n452), .A4(new_n440), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n238), .A2(G146), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n451), .A2(new_n453), .B1(new_n243), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  XOR2_X1   g270(.A(G113), .B(G122), .Z(new_n457));
  XOR2_X1   g271(.A(KEYINPUT94), .B(G104), .Z(new_n458));
  XOR2_X1   g272(.A(new_n457), .B(new_n458), .Z(new_n459));
  NAND3_X1  g273(.A1(new_n448), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n459), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n436), .A2(new_n441), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n237), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT19), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n464), .B1(new_n252), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT78), .B1(new_n465), .B2(new_n464), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n235), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(G146), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n461), .B1(new_n470), .B2(new_n455), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n460), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(G475), .A2(G902), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n432), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  AOI211_X1 g289(.A(KEYINPUT20), .B(new_n475), .C1(new_n460), .C2(new_n471), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n448), .A2(new_n456), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n461), .ZN(new_n478));
  AOI21_X1  g292(.A(G902), .B1(new_n478), .B2(new_n460), .ZN(new_n479));
  INV_X1    g293(.A(G475), .ZN(new_n480));
  OAI22_X1  g294(.A1(new_n474), .A2(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n329), .A2(G128), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n204), .A2(G143), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n482), .A2(new_n483), .A3(new_n313), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n346), .A2(G122), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n346), .A2(G122), .ZN(new_n486));
  OAI21_X1  g300(.A(G107), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G116), .B(G122), .ZN(new_n488));
  INV_X1    g302(.A(G107), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n484), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT13), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n483), .B1(new_n482), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n492), .B1(new_n204), .B2(G143), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n482), .A2(KEYINPUT96), .A3(new_n492), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n491), .B1(new_n313), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT97), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n313), .B1(new_n482), .B2(new_n483), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n490), .B1(new_n484), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n346), .A2(G122), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT14), .ZN(new_n504));
  OAI21_X1  g318(.A(G107), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(new_n504), .B2(new_n488), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n500), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n501), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n482), .A2(new_n483), .A3(new_n313), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n489), .B1(new_n485), .B2(KEYINPUT14), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n488), .A2(new_n504), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n510), .A2(new_n513), .A3(KEYINPUT97), .A4(new_n490), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n499), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G217), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n430), .A2(new_n516), .A3(G953), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n499), .A2(new_n507), .A3(new_n514), .A4(new_n517), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n261), .ZN(new_n522));
  INV_X1    g336(.A(G478), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G952), .ZN(new_n526));
  AOI211_X1 g340(.A(G953), .B(new_n526), .C1(G234), .C2(G237), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n261), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT21), .B(G898), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(G902), .B1(new_n519), .B2(new_n520), .ZN(new_n532));
  INV_X1    g346(.A(new_n524), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n525), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT98), .B1(new_n481), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n472), .A2(new_n473), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT20), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n472), .A2(new_n432), .A3(new_n473), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n532), .A2(new_n533), .ZN(new_n541));
  AOI211_X1 g355(.A(G902), .B(new_n524), .C1(new_n519), .C2(new_n520), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n541), .A2(new_n542), .A3(new_n530), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n478), .A2(new_n460), .ZN(new_n544));
  OAI21_X1  g358(.A(G475), .B1(new_n544), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT98), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n540), .A2(new_n543), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n536), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT89), .B(G469), .Z(new_n549));
  XNOR2_X1  g363(.A(G110), .B(G140), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n194), .A2(G227), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n489), .A2(G104), .ZN(new_n555));
  OR2_X1    g369(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n556));
  NAND2_X1  g370(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G104), .ZN(new_n559));
  OAI22_X1  g373(.A1(new_n559), .A2(G107), .B1(KEYINPUT86), .B2(KEYINPUT3), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(G107), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(G101), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n559), .A2(G107), .ZN(new_n564));
  AND2_X1   g378(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n565));
  NOR2_X1   g379(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G101), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n561), .A4(new_n560), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n563), .A2(KEYINPUT4), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT4), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n571), .B(G101), .C1(new_n558), .C2(new_n562), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n355), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n361), .A2(KEYINPUT87), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT87), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n332), .A2(new_n576), .A3(KEYINPUT1), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(G128), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n337), .B1(new_n578), .B2(new_n328), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n555), .A2(new_n561), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G101), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n569), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n574), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n339), .A2(KEYINPUT10), .A3(new_n569), .A4(new_n581), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n573), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n585), .A2(new_n324), .ZN(new_n586));
  INV_X1    g400(.A(new_n324), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n573), .A2(new_n583), .A3(new_n584), .A4(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n554), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n554), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n365), .A2(new_n582), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT88), .B1(new_n579), .B2(new_n582), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT88), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n365), .A2(new_n582), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n324), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n593), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n599), .A2(new_n324), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n594), .B(KEYINPUT88), .C1(new_n582), .C2(new_n579), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT12), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n592), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n590), .B1(new_n605), .B2(KEYINPUT90), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT90), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n607), .B(new_n592), .C1(new_n604), .C2(new_n601), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n261), .B(new_n549), .C1(new_n606), .C2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n586), .A2(new_n592), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n597), .A2(new_n593), .A3(new_n600), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT12), .B1(new_n602), .B2(new_n603), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n588), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n610), .B1(new_n613), .B2(new_n554), .ZN(new_n614));
  OAI21_X1  g428(.A(G469), .B1(new_n614), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G214), .B1(G237), .B2(G902), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(G210), .B1(G237), .B2(G902), .ZN(new_n619));
  INV_X1    g433(.A(G113), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT91), .B(KEYINPUT5), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(new_n347), .ZN(new_n622));
  INV_X1    g436(.A(new_n351), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n622), .B1(new_n623), .B2(new_n621), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n351), .A2(new_n352), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n582), .ZN(new_n626));
  XNOR2_X1  g440(.A(G110), .B(G122), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT8), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n351), .A2(KEYINPUT5), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n629), .A2(new_n622), .B1(new_n351), .B2(new_n352), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n626), .B(new_n628), .C1(new_n630), .C2(new_n582), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n353), .A2(new_n570), .A3(new_n572), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n624), .A2(new_n625), .A3(new_n569), .A4(new_n581), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n627), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n355), .A2(G125), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n365), .B2(G125), .ZN(new_n636));
  INV_X1    g450(.A(G224), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(G953), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(KEYINPUT7), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(KEYINPUT7), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n635), .B(new_n641), .C1(G125), .C2(new_n365), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n631), .A2(new_n634), .A3(new_n640), .A4(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n643), .A2(new_n261), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n632), .A2(new_n633), .ZN(new_n645));
  INV_X1    g459(.A(new_n627), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(KEYINPUT6), .A3(new_n634), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n636), .B(new_n639), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT6), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n645), .A2(new_n650), .A3(new_n646), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n619), .B1(new_n644), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n644), .A2(new_n652), .A3(new_n619), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n618), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND4_X1   g470(.A1(new_n431), .A2(new_n548), .A3(new_n616), .A4(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n429), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT99), .B(G101), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G3));
  NAND2_X1  g475(.A1(new_n281), .A2(new_n428), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(G472), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n419), .B(new_n261), .C1(KEYINPUT100), .C2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(KEYINPUT100), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n408), .B2(G902), .ZN(new_n667));
  INV_X1    g481(.A(new_n431), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n609), .B2(new_n615), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n523), .A2(G902), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n521), .A2(KEYINPUT102), .A3(KEYINPUT33), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT33), .B1(new_n521), .B2(KEYINPUT102), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n522), .A2(new_n676), .A3(new_n523), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT103), .B1(new_n532), .B2(G478), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(new_n481), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n644), .A2(new_n652), .A3(new_n619), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n684), .A2(new_n653), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n617), .B1(new_n655), .B2(KEYINPUT101), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n531), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n671), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT34), .B(G104), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G6));
  OR2_X1    g506(.A1(new_n686), .A2(new_n687), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n541), .A2(new_n542), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n540), .A3(new_n545), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n531), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n671), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT105), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT35), .B(G107), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G9));
  NOR2_X1   g516(.A1(new_n199), .A2(KEYINPUT36), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n265), .B(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n277), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n272), .A2(new_n276), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT106), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n667), .A2(new_n665), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n272), .A2(new_n711), .A3(new_n276), .A4(new_n707), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n709), .A2(new_n657), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT37), .B(G110), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G12));
  NAND3_X1  g529(.A1(new_n421), .A2(new_n426), .A3(new_n669), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n709), .A2(new_n712), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n481), .A2(new_n694), .ZN(new_n718));
  INV_X1    g532(.A(G900), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n527), .B1(new_n528), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n688), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n716), .A2(new_n717), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n204), .ZN(G30));
  NOR2_X1   g538(.A1(new_n684), .A2(new_n653), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n725), .B(new_n726), .Z(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n481), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n728), .A2(new_n618), .A3(new_n729), .A4(new_n694), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n720), .B(KEYINPUT39), .Z(new_n731));
  NAND2_X1  g545(.A1(new_n669), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n732), .A2(KEYINPUT40), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(KEYINPUT40), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n412), .B1(new_n400), .B2(new_n402), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n373), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n386), .A2(new_n373), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n261), .ZN(new_n738));
  OAI21_X1  g552(.A(G472), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n424), .A2(new_n425), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT82), .B1(new_n275), .B2(new_n190), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n271), .B(new_n189), .C1(new_n274), .C2(new_n268), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n741), .A2(new_n742), .A3(new_n706), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n730), .A2(new_n733), .A3(new_n734), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G143), .ZN(G45));
  NAND3_X1  g560(.A1(new_n680), .A2(new_n481), .A3(new_n721), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n686), .A2(new_n747), .A3(new_n687), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n709), .A2(new_n712), .A3(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n421), .A2(new_n426), .A3(new_n669), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT108), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n709), .A2(new_n712), .A3(new_n748), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n753), .B2(new_n716), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G146), .ZN(G48));
  OAI21_X1  g570(.A(new_n261), .B1(new_n606), .B2(new_n608), .ZN(new_n757));
  OAI21_X1  g571(.A(G469), .B1(new_n757), .B2(KEYINPUT109), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n611), .A2(new_n612), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n607), .B1(new_n760), .B2(new_n592), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n605), .A2(KEYINPUT90), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n590), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n759), .B1(new_n763), .B2(new_n261), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n431), .B(new_n609), .C1(new_n758), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT110), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n757), .A2(KEYINPUT109), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n759), .A3(new_n261), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(G469), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n431), .A4(new_n609), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n772), .A2(new_n429), .A3(new_n689), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT41), .B(G113), .Z(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G15));
  NOR3_X1   g589(.A1(new_n772), .A2(new_n429), .A3(new_n698), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n346), .ZN(G18));
  AND3_X1   g591(.A1(new_n421), .A2(new_n426), .A3(new_n548), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n765), .A2(new_n693), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n709), .A3(new_n712), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G119), .ZN(G21));
  NOR4_X1   g595(.A1(new_n693), .A2(new_n729), .A3(new_n530), .A4(new_n694), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n403), .B(KEYINPUT31), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n387), .A2(new_n373), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n423), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n419), .A2(new_n261), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n785), .B1(new_n786), .B2(G472), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n280), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n782), .A2(new_n789), .A3(new_n766), .A4(new_n771), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G122), .ZN(G24));
  NAND3_X1  g605(.A1(new_n748), .A2(new_n787), .A3(new_n708), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n765), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n214), .ZN(G27));
  INV_X1    g608(.A(KEYINPUT42), .ZN(new_n795));
  INV_X1    g609(.A(new_n747), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n684), .A2(new_n653), .A3(new_n618), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n669), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n795), .B1(new_n429), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n795), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n272), .A2(new_n276), .A3(new_n279), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n424), .A2(new_n425), .A3(new_n390), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n801), .A2(new_n802), .A3(KEYINPUT111), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT111), .B1(new_n801), .B2(new_n802), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G131), .ZN(G33));
  AND2_X1   g621(.A1(new_n669), .A2(new_n797), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n718), .A3(new_n721), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n429), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(new_n313), .ZN(G36));
  INV_X1    g625(.A(new_n710), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n729), .A2(new_n680), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT43), .Z(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n708), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT44), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n797), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT112), .Z(new_n818));
  OAI21_X1  g632(.A(G469), .B1(new_n614), .B2(KEYINPUT45), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(KEYINPUT45), .B2(new_n614), .ZN(new_n820));
  INV_X1    g634(.A(G469), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n261), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(KEYINPUT46), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n609), .B1(new_n823), .B2(KEYINPUT46), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n431), .B(new_n731), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n816), .B2(new_n815), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n818), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G137), .ZN(G39));
  OAI21_X1  g643(.A(new_n431), .B1(new_n824), .B2(new_n825), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT47), .Z(new_n831));
  NAND2_X1  g645(.A1(new_n796), .A2(new_n797), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n832), .B(new_n663), .C1(new_n421), .C2(new_n426), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n831), .A2(KEYINPUT113), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G140), .ZN(G42));
  OR4_X1    g653(.A1(new_n280), .A2(new_n668), .A3(new_n618), .A4(new_n813), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n842), .A2(new_n843), .A3(new_n740), .A4(new_n727), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n769), .A2(new_n609), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT115), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT49), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(KEYINPUT49), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n743), .A2(new_n711), .ZN(new_n850));
  INV_X1    g664(.A(new_n712), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n850), .A2(new_n851), .A3(new_n722), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n793), .B1(new_n852), .B2(new_n750), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n693), .A2(new_n729), .A3(new_n694), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n744), .A2(new_n854), .A3(new_n669), .A4(new_n721), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT108), .B1(new_n749), .B2(new_n750), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n753), .A2(new_n716), .A3(new_n752), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n853), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT52), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n808), .A2(new_n708), .A3(new_n796), .A4(new_n787), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n429), .B2(new_n809), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n695), .A2(new_n481), .A3(new_n720), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n808), .A2(new_n421), .A3(new_n426), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n717), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n617), .B(new_n531), .C1(new_n684), .C2(new_n653), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n696), .A2(KEYINPUT116), .B1(new_n680), .B2(new_n481), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n718), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n866), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n670), .A2(new_n281), .A3(new_n428), .A4(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n871), .B(new_n713), .C1(new_n429), .C2(new_n658), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n865), .A2(new_n873), .A3(new_n806), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n755), .A2(new_n875), .A3(new_n853), .A4(new_n855), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n780), .A2(new_n790), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n877), .A2(new_n773), .A3(new_n776), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n859), .A2(new_n874), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n853), .A2(new_n875), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(KEYINPUT53), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n885));
  INV_X1    g699(.A(new_n773), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n772), .A2(new_n429), .A3(new_n698), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n780), .A4(new_n790), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n865), .A2(new_n873), .A3(new_n806), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n882), .A2(new_n880), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n876), .A3(new_n859), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n885), .B1(KEYINPUT54), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n797), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n765), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT117), .ZN(new_n897));
  INV_X1    g711(.A(new_n527), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n662), .A2(new_n898), .A3(new_n740), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n729), .A3(new_n679), .A4(new_n675), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT118), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n814), .A2(new_n527), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(new_n789), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n846), .A2(new_n431), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n797), .B(new_n904), .C1(new_n831), .C2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n727), .A2(new_n765), .A3(new_n617), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT50), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n788), .A2(new_n743), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n897), .A2(new_n903), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n902), .A2(new_n906), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n803), .A2(new_n804), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n900), .A2(new_n683), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n526), .B(G953), .C1(new_n904), .C2(new_n779), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n920), .A2(new_n921), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NOR4_X1   g738(.A1(new_n894), .A2(new_n915), .A3(new_n916), .A4(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(G952), .A2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n849), .B1(new_n925), .B2(new_n926), .ZN(G75));
  NOR2_X1   g741(.A1(new_n194), .A2(G952), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n893), .A2(G210), .A3(G902), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n648), .A2(new_n651), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n649), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT55), .Z(new_n935));
  AOI21_X1  g749(.A(KEYINPUT120), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n937));
  INV_X1    g751(.A(new_n935), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n937), .B(new_n938), .C1(new_n930), .C2(new_n931), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n929), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n893), .B2(G902), .ZN(new_n942));
  AOI211_X1 g756(.A(KEYINPUT121), .B(new_n261), .C1(new_n881), .C2(new_n892), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n619), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n935), .A2(KEYINPUT56), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OR3_X1    g760(.A1(new_n944), .A2(KEYINPUT122), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT122), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n940), .B1(new_n947), .B2(new_n948), .ZN(G51));
  XNOR2_X1  g763(.A(new_n893), .B(KEYINPUT54), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n822), .B(KEYINPUT57), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n763), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n942), .A2(new_n943), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n820), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n928), .B1(new_n953), .B2(new_n955), .ZN(G54));
  NAND2_X1  g770(.A1(new_n893), .A2(G902), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(KEYINPUT121), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n893), .A2(new_n941), .A3(G902), .ZN(new_n959));
  AND2_X1   g773(.A1(KEYINPUT58), .A2(G475), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n472), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(KEYINPUT124), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n472), .A2(new_n960), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n964), .B1(new_n954), .B2(new_n965), .ZN(new_n966));
  AND4_X1   g780(.A1(new_n964), .A2(new_n958), .A3(new_n959), .A4(new_n965), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n472), .B1(new_n954), .B2(new_n960), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n929), .B1(new_n969), .B2(KEYINPUT124), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n968), .A2(new_n970), .ZN(G60));
  OR2_X1    g785(.A1(new_n673), .A2(new_n674), .ZN(new_n972));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT59), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n950), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n894), .B2(new_n974), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n975), .A2(new_n976), .A3(new_n928), .ZN(G63));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT60), .Z(new_n979));
  NAND2_X1  g793(.A1(new_n893), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n256), .B2(new_n259), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n929), .C1(new_n705), .C2(new_n980), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n529), .B2(new_n637), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n888), .A2(new_n872), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n933), .B1(G898), .B2(new_n194), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT125), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n986), .B(new_n988), .ZN(G69));
  OAI21_X1  g803(.A(new_n400), .B1(KEYINPUT30), .B2(new_n379), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n466), .A2(new_n468), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n990), .B(new_n991), .Z(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n719), .B2(new_n194), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n755), .A2(new_n853), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n917), .A2(new_n854), .ZN(new_n995));
  INV_X1    g809(.A(new_n826), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n810), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n828), .A2(new_n806), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n836), .B2(new_n837), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n993), .B1(new_n999), .B2(new_n194), .ZN(new_n1000));
  INV_X1    g814(.A(new_n429), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n895), .B1(new_n867), .B2(new_n869), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1001), .A2(new_n669), .A3(new_n731), .A4(new_n1002), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n828), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n994), .A2(new_n745), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1004), .A2(new_n838), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n992), .B1(new_n1008), .B2(new_n194), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1000), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT126), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1010), .B(new_n1012), .Z(G72));
  INV_X1    g827(.A(new_n736), .ZN(new_n1014));
  OR3_X1    g828(.A1(new_n1008), .A2(new_n888), .A3(new_n872), .ZN(new_n1015));
  XNOR2_X1  g829(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n664), .A2(new_n261), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1016), .B(new_n1017), .Z(new_n1018));
  AOI21_X1  g832(.A(new_n1014), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1018), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1020), .B1(new_n999), .B2(new_n985), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n929), .B1(new_n1021), .B2(new_n381), .ZN(new_n1022));
  AND4_X1   g836(.A1(new_n381), .A2(new_n884), .A3(new_n1014), .A4(new_n1018), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .ZN(G57));
endmodule


