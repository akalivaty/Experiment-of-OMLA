//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XOR2_X1   g0007(.A(KEYINPUT64), .B(G238), .Z(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(new_n203), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G87), .A2(G250), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n207), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n207), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n222), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g0028(.A1(new_n218), .A2(new_n219), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT66), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  OR2_X1    g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G222), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G223), .A2(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(new_n223), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n253), .B(new_n255), .C1(G77), .C2(new_n249), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(G274), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n256), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(G179), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n223), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(new_n263), .B2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n224), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n275), .A2(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(G20), .B2(new_n204), .ZN(new_n281));
  INV_X1    g0081(.A(new_n271), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n273), .B1(G50), .B2(new_n274), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n268), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n269), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n268), .A2(G200), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(new_n268), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n283), .B(KEYINPUT69), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT69), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n283), .B(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n291), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(new_n293), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(new_n291), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n287), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  INV_X1    g0106(.A(G238), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n262), .B1(new_n265), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  INV_X1    g0109(.A(new_n249), .ZN(new_n310));
  INV_X1    g0110(.A(G232), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G1698), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G226), .B2(G1698), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n309), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n308), .B1(new_n314), .B2(new_n255), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n306), .B1(new_n315), .B2(KEYINPUT71), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(KEYINPUT71), .B2(new_n315), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n317), .A2(G190), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G13), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G1), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT12), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n203), .A2(G20), .ZN(new_n324));
  INV_X1    g0124(.A(new_n274), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(KEYINPUT12), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n324), .B1(new_n276), .B2(new_n327), .C1(new_n279), .C2(new_n201), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n328), .A2(new_n271), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n326), .B1(new_n329), .B2(KEYINPUT11), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT12), .ZN(new_n331));
  OAI21_X1  g0131(.A(G68), .B1(new_n272), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n330), .B(new_n332), .C1(KEYINPUT11), .C2(new_n329), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n315), .A2(new_n318), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(new_n319), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n320), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n317), .A2(G179), .A3(new_n319), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n284), .B1(new_n335), .B2(new_n319), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT72), .B(KEYINPUT14), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n341), .B1(new_n340), .B2(new_n342), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n338), .B1(new_n339), .B2(new_n340), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n337), .B1(new_n345), .B2(new_n333), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n250), .A2(G232), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n249), .B(new_n347), .C1(new_n208), .C2(new_n250), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n255), .C1(G107), .C2(new_n249), .ZN(new_n349));
  INV_X1    g0149(.A(G244), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n262), .C1(new_n350), .C2(new_n265), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G200), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n289), .B2(new_n351), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n272), .A2(G77), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT68), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n356), .A2(new_n276), .B1(new_n224), .B2(new_n327), .ZN(new_n357));
  INV_X1    g0157(.A(new_n275), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(new_n278), .B2(new_n358), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n355), .B1(G77), .B2(new_n274), .C1(new_n282), .C2(new_n359), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n351), .A2(new_n284), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(new_n362), .C1(G179), .C2(new_n351), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n305), .A2(new_n346), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(G223), .A2(G1698), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n249), .B(new_n365), .C1(G226), .C2(new_n250), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G33), .A2(G87), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n366), .A2(KEYINPUT75), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT75), .B1(new_n366), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n255), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n262), .ZN(new_n371));
  OR3_X1    g0171(.A1(new_n265), .A2(KEYINPUT76), .A3(new_n311), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT76), .B1(new_n265), .B2(new_n311), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(G179), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n370), .A2(new_n374), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n284), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n358), .A2(new_n274), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n272), .B2(new_n358), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n202), .A2(new_n203), .ZN(new_n380));
  NOR2_X1   g0180(.A1(G58), .A2(G68), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G159), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n279), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n247), .A2(new_n224), .A3(new_n248), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n224), .A4(new_n248), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G68), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n384), .B1(new_n390), .B2(KEYINPUT74), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n203), .B1(new_n387), .B2(new_n388), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT74), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT16), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n392), .A2(new_n384), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n271), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n379), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n377), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n379), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n391), .A2(new_n394), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n398), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n334), .B1(new_n370), .B2(new_n374), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(G190), .B2(new_n376), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n370), .A2(G190), .A3(new_n374), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n376), .B2(new_n334), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT17), .B1(new_n414), .B2(new_n399), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n415), .A3(KEYINPUT77), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT77), .B1(new_n412), .B2(new_n415), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n402), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n364), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n263), .A2(G33), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n274), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n271), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n325), .A2(KEYINPUT25), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT25), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n274), .B2(G107), .ZN(new_n427));
  AOI22_X1  g0227(.A1(G107), .A2(new_n423), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT86), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT23), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n224), .B2(G107), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n424), .A2(KEYINPUT23), .A3(G20), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G116), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n257), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n224), .ZN(new_n436));
  AND2_X1   g0236(.A1(KEYINPUT3), .A2(G33), .ZN(new_n437));
  NOR2_X1   g0237(.A1(KEYINPUT3), .A2(G33), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n224), .B(G87), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n433), .B(new_n436), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n440), .ZN(new_n443));
  AOI21_X1  g0243(.A(G20), .B1(new_n247), .B2(new_n248), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(G87), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT24), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n447));
  INV_X1    g0247(.A(new_n440), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(G87), .A3(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n431), .A2(new_n432), .B1(new_n435), .B2(new_n224), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT24), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n447), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n429), .B1(new_n453), .B2(new_n271), .ZN(new_n454));
  AOI211_X1 g0254(.A(KEYINPUT86), .B(new_n282), .C1(new_n446), .C2(new_n452), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n428), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(KEYINPUT87), .B(new_n428), .C1(new_n454), .C2(new_n455), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n249), .A2(G257), .A3(G1698), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G294), .ZN(new_n461));
  OAI21_X1  g0261(.A(G250), .B1(new_n437), .B2(new_n438), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n460), .B(new_n461), .C1(G1698), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n255), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n260), .A2(G1), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G41), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n255), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G264), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n464), .A2(G179), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(G274), .B1(new_n254), .B2(new_n223), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n464), .A2(new_n472), .A3(new_n476), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n478), .A2(KEYINPUT88), .A3(G169), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT88), .B1(new_n478), .B2(G169), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n458), .A2(new_n459), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT89), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT89), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n458), .A2(new_n481), .A3(new_n484), .A4(new_n459), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n478), .A2(G200), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n478), .A2(new_n289), .ZN(new_n487));
  OR3_X1    g0287(.A1(new_n456), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  OR2_X1    g0290(.A1(KEYINPUT81), .A2(G303), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT81), .A2(G303), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n247), .A2(new_n491), .A3(new_n248), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n250), .A2(G257), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G264), .A2(G1698), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n494), .B(new_n495), .C1(new_n437), .C2(new_n438), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(new_n496), .A3(new_n255), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n493), .A2(new_n496), .A3(new_n499), .A4(new_n255), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n469), .A2(G270), .A3(new_n259), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT80), .B1(new_n503), .B2(new_n475), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT80), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n476), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  INV_X1    g0308(.A(G97), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n224), .C1(G33), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n434), .A2(G20), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n271), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n510), .A2(KEYINPUT20), .A3(new_n271), .A4(new_n511), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n274), .A2(G116), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n423), .B2(G116), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n284), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n507), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT83), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n507), .A2(new_n523), .A3(new_n519), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT84), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT84), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n521), .A2(new_n527), .A3(new_n522), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n507), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n516), .A2(new_n518), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(G179), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n507), .A2(KEYINPUT21), .A3(new_n519), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n507), .B2(G200), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n289), .B2(new_n507), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n423), .A2(G97), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(G97), .B2(new_n274), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n279), .A2(new_n327), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  AND2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n424), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n540), .B1(new_n546), .B2(G20), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT78), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT78), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n224), .B1(new_n544), .B2(new_n545), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n540), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n389), .A2(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n539), .B1(new_n553), .B2(new_n271), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(G1698), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(G244), .C1(new_n438), .C2(new_n437), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n350), .B1(new_n247), .B2(new_n248), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n508), .C1(new_n558), .C2(KEYINPUT4), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n250), .B1(new_n462), .B2(KEYINPUT4), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n255), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n475), .B1(new_n471), .B2(G257), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n554), .B(new_n564), .C1(new_n289), .C2(new_n563), .ZN(new_n565));
  INV_X1    g0365(.A(new_n465), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT79), .B1(new_n474), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT79), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n259), .A2(new_n568), .A3(G274), .A4(new_n465), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n307), .A2(new_n250), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n350), .A2(G1698), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n437), .C2(new_n438), .ZN(new_n573));
  INV_X1    g0373(.A(new_n435), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n255), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n259), .A2(new_n566), .A3(G250), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n570), .A2(new_n576), .A3(new_n578), .A4(G190), .ZN(new_n579));
  INV_X1    g0379(.A(G87), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n509), .A3(new_n424), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n309), .A2(new_n224), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT19), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n224), .B(G68), .C1(new_n437), .C2(new_n438), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n276), .B2(new_n509), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(new_n271), .B1(new_n325), .B2(new_n356), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n423), .A2(G87), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n579), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n577), .B1(new_n569), .B2(new_n567), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n334), .B1(new_n591), .B2(new_n576), .ZN(new_n592));
  INV_X1    g0392(.A(G179), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n570), .A2(new_n576), .A3(new_n578), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n587), .A2(new_n271), .ZN(new_n595));
  OR3_X1    g0395(.A1(new_n422), .A2(new_n356), .A3(new_n271), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n356), .A2(new_n325), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(G169), .B1(new_n591), .B2(new_n576), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n590), .A2(new_n592), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n563), .A2(new_n284), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n561), .A2(new_n562), .A3(new_n593), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n547), .A2(KEYINPUT78), .B1(new_n389), .B2(G107), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n282), .B1(new_n605), .B2(new_n551), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n603), .B(new_n604), .C1(new_n606), .C2(new_n539), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n565), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n529), .A2(new_n535), .A3(new_n537), .A4(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n420), .A2(new_n490), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g0410(.A(new_n610), .B(KEYINPUT90), .Z(G372));
  NAND2_X1  g0411(.A1(new_n345), .A2(new_n333), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n337), .B2(new_n363), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n412), .A2(new_n415), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT77), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n416), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n402), .ZN(new_n619));
  INV_X1    g0419(.A(new_n304), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n303), .B1(new_n302), .B2(new_n291), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n287), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n420), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n534), .B1(new_n526), .B2(new_n528), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n481), .A2(new_n456), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n565), .A2(new_n607), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n576), .A2(KEYINPUT91), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT91), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n575), .A2(new_n631), .A3(new_n255), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n591), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G200), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT92), .ZN(new_n635));
  INV_X1    g0435(.A(new_n590), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT92), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(new_n637), .A3(G200), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n488), .A2(new_n629), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n628), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n603), .A2(new_n604), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n554), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n633), .A2(new_n284), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n645), .A2(new_n594), .A3(new_n598), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n639), .A2(new_n643), .A3(new_n644), .A4(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT26), .B1(new_n607), .B2(new_n601), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n647), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n624), .B1(new_n625), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n651), .B(KEYINPUT93), .Z(G369));
  NAND2_X1  g0452(.A1(new_n322), .A2(new_n224), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n531), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n626), .A2(new_n537), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n626), .B2(new_n659), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n458), .A2(new_n459), .A3(new_n658), .ZN(new_n664));
  INV_X1    g0464(.A(new_n658), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n489), .A2(new_n664), .B1(new_n482), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n481), .A2(new_n456), .A3(new_n665), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n626), .A2(new_n658), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n490), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n220), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G1), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n581), .A2(G116), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n675), .A2(new_n676), .B1(new_n226), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n658), .B1(new_n641), .B2(new_n649), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(KEYINPUT29), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n483), .A2(new_n626), .A3(new_n485), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n640), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n644), .B1(new_n607), .B2(new_n601), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT94), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(KEYINPUT94), .B(new_n644), .C1(new_n607), .C2(new_n601), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n639), .A2(new_n643), .A3(KEYINPUT26), .A4(new_n646), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n646), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(KEYINPUT95), .A3(new_n665), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT95), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n689), .B1(new_n640), .B2(new_n681), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n658), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n680), .B1(new_n696), .B2(KEYINPUT29), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n483), .A2(new_n485), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n609), .A3(new_n488), .A4(new_n665), .ZN(new_n700));
  INV_X1    g0500(.A(new_n563), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n591), .A2(new_n576), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n473), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  OR3_X1    g0504(.A1(new_n703), .A2(new_n704), .A3(new_n507), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n530), .A2(new_n701), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n593), .A3(new_n478), .A4(new_n633), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n704), .B1(new_n703), .B2(new_n507), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n658), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n698), .B1(new_n700), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n697), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n678), .B1(new_n716), .B2(G1), .ZN(G364));
  NAND3_X1  g0517(.A1(new_n224), .A2(G13), .A3(G45), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n674), .A2(G1), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n663), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G330), .B2(new_n661), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n223), .B1(G20), .B2(new_n284), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G179), .A2(G200), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n224), .B1(new_n725), .B2(G190), .ZN(new_n726));
  INV_X1    g0526(.A(G294), .ZN(new_n727));
  INV_X1    g0527(.A(G303), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n224), .A2(new_n289), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n334), .A2(G179), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI221_X1 g0531(.A(new_n310), .B1(new_n726), .B2(new_n727), .C1(new_n728), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n224), .A2(G190), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n593), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G311), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n729), .A2(new_n734), .ZN(new_n738));
  INV_X1    g0538(.A(G322), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n733), .A2(new_n730), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n733), .A2(new_n725), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n744), .A2(G329), .ZN(new_n745));
  NOR4_X1   g0545(.A1(new_n732), .A2(new_n737), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G326), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n224), .A2(new_n593), .A3(new_n334), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT98), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n289), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n749), .A2(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT33), .B(G317), .Z(new_n754));
  OAI221_X1 g0554(.A(new_n746), .B1(new_n747), .B2(new_n751), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G50), .A2(new_n750), .B1(new_n752), .B2(G68), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n743), .A2(new_n383), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT32), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n740), .A2(new_n424), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n731), .A2(new_n580), .ZN(new_n760));
  INV_X1    g0560(.A(new_n738), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n759), .B(new_n760), .C1(G58), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n726), .A2(new_n509), .ZN(new_n763));
  INV_X1    g0563(.A(new_n735), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n310), .B(new_n763), .C1(G77), .C2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n756), .A2(new_n758), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n724), .B1(new_n755), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT97), .Z(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n723), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n310), .A2(new_n220), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n260), .B2(new_n227), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(new_n242), .B2(new_n260), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT96), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n672), .B(new_n310), .C1(new_n775), .C2(G355), .ZN(new_n776));
  OR2_X1    g0576(.A1(G355), .A2(new_n775), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n776), .A2(new_n777), .B1(new_n434), .B2(new_n672), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n719), .B(new_n767), .C1(new_n771), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n770), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n661), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n722), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(G396));
  OR2_X1    g0584(.A1(new_n363), .A2(new_n658), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n360), .A2(new_n658), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n361), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n363), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n679), .B(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(new_n715), .Z(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n719), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n723), .A2(new_n768), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n789), .A2(new_n769), .B1(G77), .B2(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n424), .A2(new_n731), .B1(new_n738), .B2(new_n727), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n310), .B1(new_n735), .B2(new_n434), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n740), .A2(new_n580), .B1(new_n743), .B2(new_n736), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n763), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n799), .B1(new_n751), .B2(new_n728), .C1(new_n741), .C2(new_n753), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT99), .B(G143), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n761), .A2(new_n801), .B1(new_n764), .B2(G159), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(new_n751), .B2(new_n803), .C1(new_n277), .C2(new_n753), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT100), .Z(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  INV_X1    g0606(.A(G132), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n249), .B1(new_n743), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT101), .ZN(new_n809));
  INV_X1    g0609(.A(new_n740), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G68), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n201), .B2(new_n731), .ZN(new_n812));
  INV_X1    g0612(.A(new_n726), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G58), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n806), .A2(new_n809), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n800), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n795), .B1(new_n817), .B2(new_n723), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n792), .B1(new_n719), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT102), .Z(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G384));
  OR2_X1    g0621(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n822), .A2(G116), .A3(new_n225), .A4(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT36), .Z(new_n825));
  OAI211_X1 g0625(.A(new_n227), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n201), .A2(G68), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n263), .B(G13), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n408), .A2(new_n410), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n379), .B1(new_n398), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n377), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT103), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n408), .A2(new_n410), .B1(new_n377), .B2(new_n833), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT103), .ZN(new_n839));
  INV_X1    g0639(.A(new_n656), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n837), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n656), .B(KEYINPUT104), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n399), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n831), .A2(new_n843), .A3(new_n400), .A4(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT105), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  AOI22_X1  g0649(.A1(KEYINPUT37), .A2(new_n842), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n841), .B1(new_n617), .B2(new_n402), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n830), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n848), .A2(new_n849), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n835), .A2(new_n836), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n841), .B1(new_n838), .B2(KEYINPUT103), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n419), .A2(new_n840), .A3(new_n833), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n700), .A2(new_n714), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n333), .A2(new_n658), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n346), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n333), .B(new_n658), .C1(new_n345), .C2(new_n337), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n861), .A2(new_n865), .A3(new_n789), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT40), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n831), .A2(new_n400), .A3(new_n845), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n848), .A2(new_n849), .B1(KEYINPUT37), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n845), .B1(new_n402), .B2(new_n614), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n830), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n868), .B1(new_n859), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n866), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n869), .A2(G330), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n420), .A2(new_n715), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT106), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n867), .A2(new_n868), .B1(new_n866), .B2(new_n874), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n420), .A3(new_n861), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n786), .B1(new_n679), .B2(new_n789), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n860), .A2(new_n865), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n402), .B2(new_n844), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n345), .A2(new_n333), .A3(new_n665), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n850), .A2(new_n851), .A3(new_n830), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n857), .B2(new_n858), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT39), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n859), .A2(new_n873), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n887), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n624), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n697), .B2(new_n420), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n894), .B(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n882), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(KEYINPUT107), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n263), .B1(G13), .B2(new_n224), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n882), .B2(new_n897), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT107), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n902), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n829), .B1(new_n900), .B2(new_n904), .ZN(G367));
  OAI21_X1  g0705(.A(new_n771), .B1(new_n220), .B2(new_n356), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n236), .A2(new_n220), .A3(new_n310), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n720), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n750), .A2(new_n801), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n752), .A2(G159), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n738), .A2(new_n277), .B1(new_n735), .B2(new_n201), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n731), .A2(new_n202), .B1(new_n743), .B2(new_n803), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n249), .B1(new_n740), .B2(new_n327), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(G68), .B2(new_n813), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n909), .A2(new_n910), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n727), .A2(new_n753), .B1(new_n751), .B2(new_n736), .ZN(new_n917));
  INV_X1    g0717(.A(new_n731), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G116), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT46), .ZN(new_n920));
  INV_X1    g0720(.A(G317), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n743), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n740), .A2(new_n509), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(G283), .C2(new_n764), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n491), .A2(new_n492), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n310), .B1(new_n926), .B2(new_n738), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(G107), .B2(new_n813), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n920), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n916), .B1(new_n917), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT111), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT47), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n908), .B1(new_n932), .B2(new_n723), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n588), .A2(new_n589), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n658), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n639), .A2(new_n646), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n646), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n933), .B1(new_n781), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n629), .B1(new_n554), .B2(new_n665), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n643), .A2(new_n658), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n670), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n607), .B1(new_n699), .B2(new_n939), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n944), .A2(new_n945), .B1(new_n665), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT108), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT108), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT109), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n947), .A2(new_n955), .A3(new_n948), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n954), .B1(new_n953), .B2(new_n956), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n958), .A2(new_n959), .B1(new_n667), .B2(new_n942), .ZN(new_n960));
  INV_X1    g0760(.A(new_n959), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n667), .A2(new_n942), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n962), .A3(new_n957), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n673), .B(KEYINPUT41), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n670), .A2(new_n668), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n942), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT110), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT44), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n967), .A2(KEYINPUT110), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n970), .B1(new_n969), .B2(new_n971), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n670), .A2(new_n668), .A3(new_n941), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT45), .Z(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n667), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n670), .B1(new_n666), .B2(new_n669), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n662), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n716), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n972), .A2(new_n667), .A3(new_n973), .A4(new_n975), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n978), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n965), .B1(new_n985), .B2(new_n716), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n718), .A2(G1), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n938), .B1(new_n964), .B2(new_n988), .ZN(G387));
  AOI211_X1 g0789(.A(G45), .B(new_n676), .C1(G68), .C2(G77), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n275), .A2(G50), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT50), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n772), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n233), .B2(new_n260), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n310), .A2(new_n672), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n995), .A2(new_n676), .B1(new_n424), .B2(new_n672), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(KEYINPUT112), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n771), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT112), .B1(new_n994), .B2(new_n996), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n720), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G159), .A2(new_n750), .B1(new_n752), .B2(new_n358), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n738), .A2(new_n201), .B1(new_n735), .B2(new_n203), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n726), .A2(new_n356), .ZN(new_n1003));
  NOR4_X1   g0803(.A1(new_n1002), .A2(new_n923), .A3(new_n1003), .A4(new_n310), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n731), .A2(new_n327), .B1(new_n743), .B2(new_n277), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT113), .Z(new_n1006));
  NAND3_X1  g0806(.A1(new_n1001), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n918), .A2(G294), .B1(new_n813), .B2(G283), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G317), .A2(new_n761), .B1(new_n764), .B2(new_n925), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n751), .B2(new_n739), .C1(new_n736), .C2(new_n753), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT114), .Z(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT49), .Z(new_n1016));
  OAI221_X1 g0816(.A(new_n310), .B1(new_n743), .B2(new_n747), .C1(new_n434), .C2(new_n740), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1007), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1000), .B1(new_n1018), .B2(new_n723), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n666), .A2(new_n781), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1019), .A2(new_n1020), .B1(new_n981), .B2(new_n987), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n716), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(KEYINPUT115), .A3(new_n980), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(new_n673), .A3(new_n982), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT115), .B1(new_n1022), .B2(new_n980), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(G393));
  NAND3_X1  g0826(.A1(new_n978), .A2(new_n987), .A3(new_n984), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n771), .B1(new_n509), .B2(new_n220), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n245), .A2(new_n772), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n720), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n750), .A2(G317), .B1(G311), .B2(new_n761), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT52), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n753), .A2(new_n926), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n764), .A2(G294), .B1(new_n744), .B2(G322), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n741), .B2(new_n731), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n310), .B1(new_n726), .B2(new_n434), .C1(new_n424), .C2(new_n740), .ZN(new_n1036));
  NOR4_X1   g0836(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT116), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(KEYINPUT116), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n750), .A2(G150), .B1(G159), .B2(new_n761), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT51), .Z(new_n1041));
  OAI221_X1 g0841(.A(new_n249), .B1(new_n726), .B2(new_n327), .C1(new_n580), .C2(new_n740), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n358), .A2(new_n764), .B1(new_n744), .B2(new_n801), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n203), .B2(new_n731), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(G50), .C2(new_n752), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1038), .A2(new_n1039), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1030), .B1(new_n1047), .B2(new_n723), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n941), .B2(new_n781), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1027), .A2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n985), .A2(new_n673), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n978), .A2(new_n984), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n982), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1050), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(G390));
  OAI21_X1  g0855(.A(new_n720), .B1(new_n358), .B2(new_n794), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G128), .A2(new_n750), .B1(new_n752), .B2(G137), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n731), .A2(new_n277), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT53), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(KEYINPUT54), .B(G143), .ZN(new_n1060));
  INV_X1    g0860(.A(G125), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n735), .A2(new_n1060), .B1(new_n743), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G50), .B2(new_n810), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n249), .B1(new_n738), .B2(new_n807), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G159), .B2(new_n813), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1057), .A2(new_n1059), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n752), .A2(G107), .B1(G97), .B2(new_n764), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n741), .B2(new_n751), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT117), .Z(new_n1069));
  OAI221_X1 g0869(.A(new_n811), .B1(new_n434), .B2(new_n738), .C1(new_n727), .C2(new_n743), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n726), .A2(new_n327), .ZN(new_n1071));
  OR4_X1    g0871(.A1(new_n249), .A2(new_n1070), .A3(new_n760), .A4(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1066), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1056), .B1(new_n1073), .B2(new_n723), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n890), .A2(new_n892), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n769), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT118), .Z(new_n1077));
  NAND3_X1  g0877(.A1(new_n692), .A2(new_n695), .A3(new_n785), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n788), .A2(new_n363), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n865), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n887), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n859), .B2(new_n873), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n863), .A2(new_n864), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n887), .B1(new_n883), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n890), .A2(new_n1085), .A3(new_n892), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n715), .A2(new_n789), .A3(new_n865), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1083), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1077), .B1(new_n987), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n529), .A2(new_n535), .A3(new_n608), .A4(new_n537), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n489), .A2(new_n1092), .A3(new_n658), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n712), .A2(new_n713), .ZN(new_n1094));
  OAI211_X1 g0894(.A(G330), .B(new_n789), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1084), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n883), .B1(new_n1087), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1087), .A2(new_n1096), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT95), .B1(new_n691), .B2(new_n665), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n694), .A2(new_n693), .A3(new_n658), .ZN(new_n1103));
  OAI21_X1  g0903(.A(KEYINPUT29), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n680), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n420), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n624), .A3(new_n877), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1101), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1095), .A2(new_n1084), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1083), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n865), .B1(new_n715), .B2(new_n789), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n884), .B1(new_n1114), .B2(new_n1110), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n1098), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n896), .A3(new_n877), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1113), .A2(new_n1119), .A3(new_n673), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1091), .A2(new_n1120), .ZN(G378));
  INV_X1    g0921(.A(KEYINPUT122), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n286), .B1(new_n620), .B2(new_n621), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1124), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n305), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n292), .A2(new_n656), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1128), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1122), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1131), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(KEYINPUT122), .A3(new_n1129), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n880), .A2(new_n1135), .A3(G330), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1129), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n880), .B2(G330), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n886), .A2(new_n893), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n876), .A2(new_n1129), .A3(new_n1133), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n880), .A2(new_n1135), .A3(G330), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n894), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n987), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n720), .B1(G50), .B2(new_n794), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT121), .ZN(new_n1147));
  AOI21_X1  g0947(.A(G50), .B1(new_n248), .B2(new_n258), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G97), .A2(new_n752), .B1(new_n750), .B2(G116), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n738), .A2(new_n424), .B1(new_n743), .B2(new_n741), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n356), .A2(new_n735), .B1(new_n740), .B2(new_n202), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G68), .C2(new_n813), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n310), .B(new_n258), .C1(new_n327), .C2(new_n731), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT119), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1149), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT58), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1148), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G125), .A2(new_n750), .B1(new_n752), .B2(G132), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1159), .A2(new_n738), .B1(new_n731), .B2(new_n1060), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT120), .Z(new_n1161));
  AOI22_X1  g0961(.A1(G137), .A2(new_n764), .B1(new_n813), .B2(G150), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1158), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n257), .B(new_n258), .C1(new_n740), .C2(new_n383), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G124), .B2(new_n744), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1157), .B1(new_n1156), .B2(new_n1155), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1147), .B1(new_n1169), .B2(new_n723), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1135), .B2(new_n769), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1145), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1107), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1113), .A2(KEYINPUT123), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT123), .B1(new_n1113), .B2(new_n1174), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1144), .B(KEYINPUT57), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n673), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1144), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1173), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(G375));
  NAND2_X1  g0984(.A1(new_n1084), .A2(new_n768), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n720), .B1(G68), .B2(new_n794), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n509), .A2(new_n731), .B1(new_n738), .B2(new_n741), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n310), .B1(new_n740), .B2(new_n327), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n735), .A2(new_n424), .B1(new_n743), .B2(new_n728), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1003), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n751), .B2(new_n727), .C1(new_n434), .C2(new_n753), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n249), .B1(new_n726), .B2(new_n201), .C1(new_n202), .C2(new_n740), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n735), .A2(new_n277), .B1(new_n743), .B2(new_n1159), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n803), .A2(new_n738), .B1(new_n731), .B2(new_n383), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n751), .B2(new_n807), .C1(new_n753), .C2(new_n1060), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT125), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n724), .B1(new_n1197), .B2(KEYINPUT125), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1186), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1117), .A2(new_n987), .B1(new_n1185), .B2(new_n1200), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n965), .B(KEYINPUT124), .Z(new_n1202));
  NAND2_X1  g1002(.A1(new_n1118), .A2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1174), .A2(new_n1117), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(G381));
  OR2_X1    g1005(.A1(G393), .A2(G396), .ZN(new_n1206));
  OR4_X1    g1006(.A1(G384), .A2(G378), .A3(new_n1206), .A4(G381), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1054), .B(new_n938), .C1(new_n964), .C2(new_n988), .ZN(new_n1208));
  OR3_X1    g1008(.A1(G375), .A2(new_n1207), .A3(new_n1208), .ZN(G407));
  INV_X1    g1009(.A(G378), .ZN(new_n1210));
  INV_X1    g1010(.A(G213), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(G343), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1183), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT126), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(G407), .A3(G213), .ZN(G409));
  NAND2_X1  g1015(.A1(G387), .A2(G390), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(G393), .B(G396), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1216), .A2(new_n1208), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1216), .B2(new_n1208), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT61), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n674), .B(new_n1108), .C1(new_n1204), .C2(KEYINPUT60), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(KEYINPUT60), .B2(new_n1204), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n820), .B1(new_n1223), .B2(new_n1201), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n820), .A3(new_n1201), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1212), .A2(G2897), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1227), .B(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT123), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1118), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n1107), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1113), .A2(KEYINPUT123), .A3(new_n1174), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n1144), .A3(new_n1202), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G378), .B1(new_n1172), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1144), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G378), .B(new_n1172), .C1(new_n1178), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT127), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1182), .A2(new_n673), .A3(new_n1177), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT127), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1240), .A2(new_n1241), .A3(G378), .A4(new_n1172), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1236), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1229), .B1(new_n1243), .B2(new_n1212), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1227), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1243), .A2(new_n1212), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT62), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1221), .B(new_n1244), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1236), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1212), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1253), .A2(KEYINPUT62), .A3(new_n1245), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1220), .B1(new_n1248), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT63), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1253), .B2(new_n1245), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1229), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1246), .A2(KEYINPUT63), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1261), .ZN(G405));
  NAND2_X1  g1062(.A1(G375), .A2(new_n1210), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1220), .A2(new_n1249), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1249), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1259), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(new_n1245), .ZN(G402));
endmodule


