//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n568, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT64), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(G137), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT65), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n462), .A2(G125), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR3_X1    g053(.A1(KEYINPUT66), .A2(G100), .A3(G2105), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n463), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT66), .B1(G100), .B2(G2105), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n479), .A2(new_n480), .A3(G2104), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n476), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(G2104), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT67), .B(G114), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n487), .A2(new_n488), .B1(G126), .B2(new_n477), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n463), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n492), .A2(KEYINPUT68), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(KEYINPUT68), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n462), .A2(new_n496), .A3(G138), .A4(new_n463), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(G651), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n504), .A2(KEYINPUT69), .A3(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT6), .B1(new_n506), .B2(G651), .ZN(new_n507));
  OAI211_X1 g082(.A(G543), .B(new_n503), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n504), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n506), .A2(new_n501), .A3(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n502), .B1(KEYINPUT69), .B2(new_n504), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n515), .A2(KEYINPUT71), .A3(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XOR2_X1   g096(.A(KEYINPUT72), .B(G88), .Z(new_n522));
  NAND3_X1  g097(.A1(new_n514), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n504), .A2(KEYINPUT69), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n506), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n510), .B(new_n523), .C1(new_n524), .C2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND3_X1  g105(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n514), .A2(new_n521), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n509), .A2(G51), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n533), .A2(new_n535), .A3(new_n537), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n513), .A2(new_n512), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT74), .B(G90), .Z(new_n543));
  NAND4_X1  g118(.A1(new_n521), .A2(new_n542), .A3(new_n503), .A4(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n542), .A2(G52), .A3(G543), .A4(new_n503), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n515), .A2(KEYINPUT71), .A3(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT71), .B1(new_n515), .B2(G543), .ZN(new_n549));
  OAI211_X1 g124(.A(G64), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(new_n527), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n541), .B1(new_n546), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n544), .A2(new_n545), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n528), .B1(new_n550), .B2(new_n551), .ZN(new_n556));
  NOR3_X1   g131(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT75), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  NAND4_X1  g134(.A1(new_n542), .A2(G43), .A3(G543), .A4(new_n503), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n521), .A2(new_n542), .A3(G81), .A4(new_n503), .ZN(new_n561));
  INV_X1    g136(.A(G68), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(new_n518), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n521), .B2(G56), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n560), .B(new_n561), .C1(new_n564), .C2(new_n528), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(G188));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT9), .B1(new_n508), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n514), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n514), .A2(G91), .A3(new_n521), .ZN(new_n578));
  OAI211_X1 g153(.A(G65), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n579));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(G299));
  NAND3_X1  g158(.A1(new_n514), .A2(G49), .A3(G543), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n514), .A2(G87), .A3(new_n521), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT76), .Z(new_n589));
  OAI21_X1  g164(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(new_n527), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT77), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n514), .A2(new_n521), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  INV_X1    g171(.A(G48), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n595), .A2(new_n596), .B1(new_n597), .B2(new_n508), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n594), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n509), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OAI221_X1 g178(.A(new_n601), .B1(new_n595), .B2(new_n602), .C1(new_n528), .C2(new_n603), .ZN(G290));
  NAND4_X1  g179(.A1(new_n521), .A2(new_n542), .A3(G92), .A4(new_n503), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n514), .A2(KEYINPUT10), .A3(G92), .A4(new_n521), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n509), .A2(G54), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n590), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G651), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n609), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G171), .B2(new_n616), .ZN(G284));
  OAI21_X1  g193(.A(new_n617), .B1(G171), .B2(new_n616), .ZN(G321));
  NAND2_X1  g194(.A1(G299), .A2(new_n616), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G168), .B2(new_n616), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(G168), .B2(new_n616), .ZN(G280));
  INV_X1    g197(.A(new_n615), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n566), .ZN(G323));
  XOR2_X1   g203(.A(G323), .B(KEYINPUT78), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n475), .A2(G2104), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2100), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n477), .A2(G123), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT79), .Z(new_n636));
  OR2_X1    g211(.A1(G99), .A2(G2105), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n637), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n475), .A2(G135), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2096), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  INV_X1    g219(.A(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  OAI21_X1  g222(.A(KEYINPUT14), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT80), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2443), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT81), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n652), .A2(new_n656), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n657), .B2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n643), .B1(new_n664), .B2(G14), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n657), .A2(new_n660), .ZN(new_n666));
  INV_X1    g241(.A(new_n659), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND4_X1   g243(.A1(new_n643), .A2(new_n668), .A3(G14), .A4(new_n661), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  AOI21_X1  g251(.A(KEYINPUT18), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2072), .B(G2078), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT83), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(KEYINPUT18), .B2(new_n674), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n677), .B(new_n680), .Z(new_n681));
  XNOR2_X1  g256(.A(G2096), .B(G2100), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n684), .A2(new_n685), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n693));
  AOI21_X1  g268(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n694), .B(new_n695), .C1(new_n692), .C2(new_n693), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1996), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1981), .B(G1986), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT86), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT85), .B(G1991), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n699), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G26), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT94), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n477), .A2(G128), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT93), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(G104), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n475), .A2(G140), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n708), .B1(new_n715), .B2(new_n705), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2067), .ZN(new_n717));
  OR2_X1    g292(.A1(G29), .A2(G33), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n475), .A2(G139), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT25), .Z(new_n721));
  AOI22_X1  g296(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT95), .Z(new_n723));
  OAI211_X1 g298(.A(new_n719), .B(new_n721), .C1(new_n723), .C2(new_n463), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n718), .B1(new_n724), .B2(new_n705), .ZN(new_n725));
  INV_X1    g300(.A(G2072), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n717), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G1341), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n566), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(G19), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n705), .A2(G35), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G162), .B2(new_n705), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT29), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n728), .B1(new_n729), .B2(new_n732), .C1(G2090), .C2(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  NOR2_X1   g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n737), .A2(new_n738), .A3(G29), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n471), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT96), .Z(new_n743));
  AND2_X1   g318(.A1(new_n740), .A2(new_n741), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n640), .A2(G29), .ZN(new_n745));
  OR2_X1    g320(.A1(G29), .A2(G32), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n477), .A2(G129), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n475), .A2(G141), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n746), .B1(new_n752), .B2(new_n705), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(G28), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n758), .A2(new_n759), .A3(new_n705), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n745), .A2(new_n755), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n736), .A2(new_n743), .A3(new_n744), .A4(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(KEYINPUT97), .B1(G16), .B2(G21), .ZN(new_n763));
  NAND2_X1  g338(.A1(G168), .A2(G16), .ZN(new_n764));
  MUX2_X1   g339(.A(KEYINPUT97), .B(new_n763), .S(new_n764), .Z(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT98), .B(G1966), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n730), .A2(G4), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n623), .B2(new_n730), .ZN(new_n771));
  INV_X1    g346(.A(G1348), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n729), .A2(new_n732), .B1(new_n735), .B2(G2090), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n762), .A2(new_n768), .A3(new_n769), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n765), .A2(new_n767), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT99), .Z(new_n778));
  AND2_X1   g353(.A1(new_n725), .A2(new_n726), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n730), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n730), .ZN(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n730), .A2(G20), .ZN(new_n784));
  AND3_X1   g359(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(new_n785));
  OAI211_X1 g360(.A(KEYINPUT23), .B(new_n784), .C1(new_n785), .C2(new_n730), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT23), .B2(new_n784), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n776), .A2(new_n778), .A3(new_n779), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n705), .A2(G27), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G164), .B2(new_n705), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT100), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2078), .ZN(new_n794));
  INV_X1    g369(.A(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(KEYINPUT91), .B1(new_n795), .B2(G16), .ZN(new_n796));
  OR3_X1    g371(.A1(new_n795), .A2(KEYINPUT91), .A3(G16), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n796), .B(new_n797), .C1(G166), .C2(new_n730), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G1971), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n798), .A2(G1971), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n730), .A2(G6), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G305), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT32), .B(G1981), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT88), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n799), .B(new_n800), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n802), .A2(new_n804), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G23), .ZN(new_n807));
  INV_X1    g382(.A(G288), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G16), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT89), .B(KEYINPUT90), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT33), .B(G1976), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n805), .A2(new_n806), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT34), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n805), .A2(new_n816), .A3(new_n806), .A4(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n730), .A2(G24), .ZN(new_n818));
  INV_X1    g393(.A(G290), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n730), .ZN(new_n820));
  INV_X1    g395(.A(G1986), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n705), .A2(G25), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n475), .A2(G131), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n477), .A2(G119), .ZN(new_n825));
  OR2_X1    g400(.A1(G95), .A2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n823), .B1(new_n829), .B2(new_n705), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT87), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G1991), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n817), .A2(new_n822), .A3(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT92), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(KEYINPUT92), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n815), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI211_X1 g414(.A(KEYINPUT36), .B(new_n815), .C1(new_n835), .C2(new_n836), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n790), .B(new_n794), .C1(new_n839), .C2(new_n840), .ZN(G150));
  INV_X1    g416(.A(G150), .ZN(G311));
  XNOR2_X1  g417(.A(KEYINPUT102), .B(G860), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n521), .A2(new_n542), .A3(G93), .A4(new_n503), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n542), .A2(G55), .A3(G543), .A4(new_n503), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G67), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n590), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G80), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n518), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n527), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n843), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n850), .B1(new_n521), .B2(G67), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n845), .B(new_n844), .C1(new_n854), .C2(new_n528), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n565), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n623), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(KEYINPUT101), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(KEYINPUT101), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n843), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n859), .A2(new_n860), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n853), .B1(new_n864), .B2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(new_n715), .B(new_n499), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n752), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n632), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n868), .A2(new_n632), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n828), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n829), .A3(new_n869), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n471), .B(G162), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI22_X1  g452(.A1(G130), .A2(new_n477), .B1(new_n475), .B2(G142), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n881), .B(new_n882), .C1(G118), .C2(new_n463), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n724), .B(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n877), .A2(new_n885), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(new_n640), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n640), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n875), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n874), .A3(new_n872), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(new_n855), .A2(new_n616), .ZN(new_n898));
  NAND2_X1  g473(.A1(G303), .A2(new_n808), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n536), .A2(new_n522), .B1(G50), .B2(new_n509), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n524), .A2(new_n528), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(G288), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n899), .A2(new_n902), .A3(G290), .ZN(new_n903));
  AOI21_X1  g478(.A(G290), .B1(new_n899), .B2(new_n902), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n903), .A2(new_n904), .A3(G305), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n593), .A2(KEYINPUT77), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n593), .A2(KEYINPUT77), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n598), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(G303), .A2(new_n808), .ZN(new_n909));
  AOI21_X1  g484(.A(G288), .B1(new_n900), .B2(new_n901), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n819), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n899), .A2(new_n902), .A3(G290), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n905), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT42), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n626), .B(new_n856), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n785), .A2(new_n615), .ZN(new_n917));
  NAND4_X1  g492(.A1(G299), .A2(new_n610), .A3(new_n609), .A4(new_n614), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT41), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n918), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n922), .B1(new_n923), .B2(new_n916), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n915), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n898), .B1(new_n925), .B2(new_n616), .ZN(G295));
  OAI21_X1  g501(.A(new_n898), .B1(new_n925), .B2(new_n616), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  INV_X1    g503(.A(new_n923), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n554), .B2(new_n557), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n856), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n553), .A2(new_n541), .A3(new_n545), .A4(new_n544), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT75), .B1(new_n555), .B2(new_n556), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT105), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n935), .A2(G286), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n521), .A2(G56), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n527), .B1(new_n937), .B2(new_n563), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n561), .A2(new_n560), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n855), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n565), .A2(new_n846), .A3(new_n851), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT105), .B1(new_n933), .B2(new_n934), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n932), .A2(new_n936), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n936), .B1(new_n932), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n929), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n935), .A2(G286), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n942), .A2(new_n943), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n942), .A2(new_n943), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n932), .A2(new_n936), .A3(new_n944), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n921), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n914), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n947), .A2(new_n953), .ZN(new_n956));
  INV_X1    g531(.A(new_n914), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI211_X1 g533(.A(KEYINPUT106), .B(new_n914), .C1(new_n947), .C2(new_n953), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n895), .B(new_n954), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n928), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT44), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT107), .B1(new_n960), .B2(KEYINPUT43), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n969));
  NOR4_X1   g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n964), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n966), .A2(KEYINPUT44), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n968), .A2(new_n964), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT108), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n965), .B1(new_n970), .B2(new_n973), .ZN(G397));
  INV_X1    g549(.A(G2067), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n715), .B(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n499), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n465), .A2(G40), .A3(new_n470), .A4(new_n466), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n978), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT110), .Z(new_n982));
  XNOR2_X1  g557(.A(new_n752), .B(G1996), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n980), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n828), .B(new_n832), .Z(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(new_n821), .A3(new_n819), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n980), .A2(G1986), .A3(G290), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n990), .B(KEYINPUT109), .Z(new_n991));
  NOR2_X1   g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n908), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n598), .B(KEYINPUT113), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n995), .A2(new_n593), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n996), .B2(new_n993), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT49), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n499), .A2(new_n977), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(new_n979), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1976), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(G288), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n808), .A2(G1976), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1006), .A2(KEYINPUT112), .A3(new_n1002), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(KEYINPUT112), .A3(new_n1007), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(new_n1009), .A3(new_n1005), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n998), .A2(new_n1002), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n979), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n499), .A2(KEYINPUT50), .A3(new_n977), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT50), .B1(new_n499), .B2(new_n977), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(G2090), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n979), .B1(new_n1017), .B2(new_n999), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT111), .B1(new_n999), .B2(new_n1017), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n499), .A2(new_n1020), .A3(KEYINPUT45), .A4(new_n977), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1971), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1001), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT55), .Z(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1011), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n741), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n978), .A2(KEYINPUT45), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n766), .B1(new_n1018), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(G8), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G286), .A2(G8), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT123), .B(KEYINPUT51), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n1037), .B(KEYINPUT124), .Z(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(new_n1035), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1042));
  OAI22_X1  g617(.A1(new_n1038), .A2(new_n1041), .B1(new_n1042), .B2(new_n1037), .ZN(new_n1043));
  INV_X1    g618(.A(G2078), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1018), .A2(new_n1019), .A3(new_n1044), .A4(new_n1021), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1045), .A2(new_n1046), .B1(new_n782), .B2(new_n1015), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G171), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1018), .A2(new_n1033), .A3(KEYINPUT53), .A4(new_n1044), .ZN(new_n1051));
  AOI21_X1  g626(.A(G301), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1043), .B1(new_n1053), .B2(KEYINPUT54), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT125), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1049), .B2(G171), .ZN(new_n1056));
  AOI211_X1 g631(.A(KEYINPUT125), .B(G301), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1048), .A2(G301), .A3(new_n1051), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT54), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1956), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1015), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT56), .B(G2072), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .A4(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n578), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n504), .B1(new_n579), .B2(new_n580), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT115), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n578), .B(new_n1071), .C1(new_n1072), .C2(new_n504), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n577), .A3(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n577), .A2(KEYINPUT57), .A3(new_n578), .A4(new_n582), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT116), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT57), .A4(new_n577), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT117), .B1(new_n1076), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1083), .A2(KEYINPUT119), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1067), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1066), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1066), .A2(new_n1090), .A3(KEYINPUT122), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1089), .A2(new_n1093), .A3(KEYINPUT61), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1015), .A2(new_n772), .B1(new_n975), .B2(new_n1000), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(KEYINPUT60), .B2(new_n623), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n615), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(KEYINPUT60), .A3(new_n623), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT58), .B(G1341), .ZN(new_n1101));
  OAI22_X1  g676(.A1(new_n1022), .A2(G1996), .B1(new_n1000), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n566), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT59), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1105), .A3(new_n566), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1099), .A2(new_n1100), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1095), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1109));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1066), .A2(new_n1090), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n1066), .B2(new_n1090), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1066), .A2(new_n1090), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1109), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1096), .A2(new_n615), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1085), .B1(new_n1120), .B2(new_n1084), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1086), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1083), .A2(KEYINPUT119), .A3(new_n1086), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1118), .B1(new_n1125), .B2(new_n1067), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1091), .A2(KEYINPUT118), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1066), .A2(new_n1090), .A3(new_n1110), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1117), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1118), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1089), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n1113), .A3(KEYINPUT120), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1061), .B1(new_n1116), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1043), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT126), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1043), .A2(new_n1140), .A3(KEYINPUT62), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1138), .A2(new_n1052), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1030), .B1(new_n1135), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1035), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1011), .A2(new_n1028), .A3(new_n1029), .A4(new_n1144), .ZN(new_n1145));
  OR3_X1    g720(.A1(new_n1145), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1011), .A2(new_n1027), .A3(new_n1025), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT63), .B1(new_n1145), .B2(G286), .ZN(new_n1148));
  AOI211_X1 g723(.A(G1976), .B(G288), .C1(new_n998), .C2(new_n1002), .ZN(new_n1149));
  INV_X1    g724(.A(new_n994), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1002), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n992), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT46), .ZN(new_n1154));
  OR3_X1    g729(.A1(new_n985), .A2(new_n1154), .A3(G1996), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n980), .B1(new_n976), .B2(new_n752), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n985), .B2(G1996), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n988), .B(KEYINPUT48), .Z(new_n1161));
  NOR2_X1   g736(.A1(new_n828), .A2(new_n832), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n984), .A2(new_n1162), .B1(new_n975), .B2(new_n715), .ZN(new_n1163));
  OAI221_X1 g738(.A(new_n1160), .B1(new_n987), .B2(new_n1161), .C1(new_n1163), .C2(new_n985), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1153), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g741(.A(G227), .ZN(new_n1168));
  OAI21_X1  g742(.A(new_n1168), .B1(new_n665), .B2(new_n669), .ZN(new_n1169));
  NOR2_X1   g743(.A1(G229), .A2(new_n460), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n896), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g745(.A(new_n964), .ZN(new_n1172));
  AOI211_X1 g746(.A(new_n1169), .B(new_n1171), .C1(new_n962), .C2(new_n1172), .ZN(G308));
  AOI21_X1  g747(.A(new_n1169), .B1(new_n962), .B2(new_n1172), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n1174), .A2(new_n896), .A3(new_n1170), .ZN(G225));
endmodule


