//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT68), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AND2_X1   g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n458), .A2(G567), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n471), .B1(new_n473), .B2(G101), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n470), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n467), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n477), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n468), .A2(new_n469), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(KEYINPUT71), .ZN(new_n483));
  OR2_X1    g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n484), .A2(KEYINPUT71), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n483), .B2(new_n486), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n484), .B2(new_n485), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(KEYINPUT72), .B2(G114), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT72), .A2(G114), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2105), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G102), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(new_n472), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT3), .B(G2104), .ZN(new_n509));
  AND3_X1   g084(.A1(new_n504), .A2(KEYINPUT4), .A3(G138), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n502), .B(new_n506), .C1(G2105), .C2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(new_n520), .A3(G88), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G50), .A3(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT74), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n519), .B1(new_n525), .B2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(new_n520), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n531), .A2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n518), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT75), .B(G90), .Z(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n534), .A2(new_n540), .B1(new_n529), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n518), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT76), .B(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n534), .A2(new_n546), .B1(new_n529), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n529), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n520), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n516), .A2(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT79), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n518), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n516), .A2(new_n520), .A3(G91), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n558), .A2(KEYINPUT78), .A3(new_n559), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  XNOR2_X1  g146(.A(G168), .B(KEYINPUT80), .ZN(G286));
  INV_X1    g147(.A(new_n526), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT74), .B1(new_n521), .B2(new_n522), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n573), .A2(new_n574), .B1(new_n518), .B2(new_n517), .ZN(G303));
  OR2_X1    g150(.A1(new_n516), .A2(G74), .ZN(new_n576));
  INV_X1    g151(.A(new_n529), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n576), .A2(G651), .B1(new_n577), .B2(G49), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT81), .B1(new_n534), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n516), .A2(new_n520), .A3(new_n581), .A4(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n583), .ZN(G288));
  AND2_X1   g159(.A1(G73), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n516), .B2(G61), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n518), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n516), .A2(new_n520), .A3(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n577), .A2(G48), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n518), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n534), .A2(new_n593), .B1(new_n529), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n516), .A2(new_n520), .A3(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT10), .Z(new_n600));
  NAND2_X1  g175(.A1(new_n516), .A2(G66), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT82), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n518), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(G54), .B2(new_n577), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G321));
  NOR2_X1   g184(.A1(G299), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G286), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  AOI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  INV_X1    g190(.A(new_n549), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n606), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n509), .A2(new_n473), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n488), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n491), .A2(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n628), .A2(new_n629), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n629), .B2(new_n628), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n626), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  INV_X1    g209(.A(new_n633), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n625), .A2(new_n634), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT14), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n644), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT84), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XNOR2_X1  g231(.A(G2084), .B(G2090), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(KEYINPUT17), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n660), .B(new_n657), .C1(new_n655), .C2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n657), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n655), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n636), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT85), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n670), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1986), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  INV_X1    g258(.A(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n680), .A2(new_n681), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(new_n681), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G35), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G162), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT29), .Z(new_n695));
  INV_X1    g270(.A(G2090), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n488), .A2(G141), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n491), .A2(G129), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT26), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n703), .A2(new_n704), .B1(G105), .B2(new_n473), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n699), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(KEYINPUT94), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n699), .A2(new_n700), .A3(new_n708), .A4(new_n705), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n692), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n692), .B2(G32), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n697), .A2(new_n698), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G5), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G171), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G1961), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n549), .A2(new_n716), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n716), .B2(G19), .ZN(new_n721));
  INV_X1    g296(.A(G1341), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G168), .A2(new_n716), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n716), .B2(G21), .ZN(new_n725));
  INV_X1    g300(.A(G1966), .ZN(new_n726));
  OAI22_X1  g301(.A1(new_n725), .A2(new_n726), .B1(G1961), .B2(new_n718), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n692), .A2(G27), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G164), .B2(new_n692), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G2078), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n723), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n692), .B1(KEYINPUT24), .B2(G34), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(KEYINPUT24), .B2(G34), .ZN(new_n734));
  INV_X1    g309(.A(G160), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G29), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n721), .A2(new_n722), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT31), .B(G11), .Z(new_n738));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n692), .B1(new_n739), .B2(G28), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n740), .A2(KEYINPUT95), .B1(new_n739), .B2(G28), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n737), .B(new_n743), .C1(new_n692), .C2(new_n633), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n716), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n607), .B2(new_n716), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1348), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n692), .A2(G26), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n750));
  INV_X1    g325(.A(G104), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n467), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n491), .B2(G128), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n488), .A2(G140), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n749), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n731), .A2(new_n744), .A3(new_n747), .A4(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n725), .A2(new_n726), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT97), .B(KEYINPUT23), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n716), .A2(G20), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G299), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1956), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n692), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n509), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n467), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n488), .B2(G139), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(new_n692), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(new_n442), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n736), .A2(new_n732), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n762), .A2(new_n767), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n715), .A2(new_n760), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n716), .A2(G22), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G166), .B2(new_n716), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT90), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G1971), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n587), .A2(G16), .A3(new_n588), .A4(new_n589), .ZN(new_n786));
  OR2_X1    g361(.A1(G6), .A2(G16), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(KEYINPUT32), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT32), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n786), .A2(new_n790), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G1981), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n789), .A2(new_n684), .A3(new_n791), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n783), .A2(KEYINPUT90), .ZN(new_n796));
  INV_X1    g371(.A(G1971), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n783), .A2(KEYINPUT90), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G16), .A2(G23), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT89), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G288), .B2(new_n716), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT33), .B(G1976), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  AND4_X1   g379(.A1(new_n785), .A2(new_n795), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT88), .B(KEYINPUT34), .Z(new_n806));
  OAI21_X1  g381(.A(KEYINPUT91), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n785), .A2(new_n795), .A3(new_n799), .A4(new_n804), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n809));
  INV_X1    g384(.A(new_n806), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  INV_X1    g389(.A(KEYINPUT86), .ZN(new_n815));
  INV_X1    g390(.A(G119), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n490), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n815), .B1(new_n490), .B2(new_n816), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(new_n467), .B2(G107), .ZN(new_n821));
  INV_X1    g396(.A(G95), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n467), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n488), .B2(G131), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n692), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n692), .A2(G25), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n814), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n819), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n824), .B1(new_n828), .B2(new_n817), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n826), .B1(new_n829), .B2(G29), .ZN(new_n830));
  INV_X1    g405(.A(new_n814), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT87), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n827), .A2(new_n832), .A3(KEYINPUT87), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n716), .A2(G24), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n596), .B2(new_n716), .ZN(new_n838));
  INV_X1    g413(.A(G1986), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n835), .A2(new_n836), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n805), .B2(new_n806), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n812), .A2(new_n813), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n813), .B1(new_n812), .B2(new_n842), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n781), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n812), .A2(new_n842), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT92), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n848), .A2(KEYINPUT36), .A3(new_n843), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n780), .B1(new_n846), .B2(new_n849), .ZN(G311));
  NOR3_X1   g425(.A1(new_n844), .A2(new_n781), .A3(new_n845), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT36), .B1(new_n848), .B2(new_n843), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n779), .B1(new_n851), .B2(new_n852), .ZN(G150));
  XOR2_X1   g428(.A(KEYINPUT98), .B(G93), .Z(new_n854));
  INV_X1    g429(.A(G55), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n534), .A2(new_n854), .B1(new_n529), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT99), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(new_n518), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(KEYINPUT100), .A3(new_n859), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n616), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n857), .A2(KEYINPUT100), .A3(new_n549), .A4(new_n859), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n607), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g445(.A(G860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n860), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(G145));
  XNOR2_X1  g451(.A(new_n633), .B(KEYINPUT102), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G162), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n877), .A2(G162), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n735), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n878), .A3(G160), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n706), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n885), .A2(new_n773), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n707), .A2(new_n709), .A3(new_n773), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n829), .B(new_n623), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n623), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n829), .B(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n886), .A3(new_n887), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n755), .A2(G164), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n753), .A2(new_n512), .A3(new_n754), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n488), .A2(G142), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n491), .A2(G130), .ZN(new_n897));
  OR2_X1    g472(.A1(G106), .A2(G2105), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n898), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n894), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(new_n894), .B2(new_n895), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n890), .A2(new_n893), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n890), .B2(new_n893), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n884), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT103), .A3(new_n884), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT104), .B1(new_n911), .B2(new_n884), .ZN(new_n914));
  INV_X1    g489(.A(new_n884), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n915), .A2(new_n910), .A3(new_n916), .A4(new_n904), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n913), .A2(KEYINPUT40), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT40), .B1(new_n913), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(G395));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n922));
  XNOR2_X1  g497(.A(G305), .B(KEYINPUT105), .ZN(new_n923));
  INV_X1    g498(.A(G288), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(G166), .B(new_n596), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n923), .B(G288), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n926), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n930), .A3(KEYINPUT42), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n864), .A2(new_n619), .A3(new_n865), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n619), .B1(new_n864), .B2(new_n865), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(G299), .B(new_n606), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT41), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n607), .A2(G299), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(new_n606), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n939), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n936), .B2(new_n937), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n935), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n933), .A2(new_n947), .A3(new_n934), .A4(new_n949), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n617), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n860), .A2(new_n617), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n922), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n955), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n953), .A2(KEYINPUT106), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n956), .A2(new_n958), .ZN(G295));
  NAND2_X1  g534(.A1(new_n954), .A2(new_n955), .ZN(G331));
  NOR2_X1   g535(.A1(G171), .A2(G168), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(G286), .B2(G301), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n864), .A2(new_n865), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n864), .B2(new_n865), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n948), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n966), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n946), .A3(new_n964), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n969), .A3(new_n931), .ZN(new_n970));
  INV_X1    g545(.A(G37), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n931), .B1(new_n967), .B2(new_n969), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n940), .A2(new_n945), .A3(KEYINPUT107), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n939), .A2(new_n976), .A3(KEYINPUT41), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n968), .A2(new_n975), .A3(new_n964), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n967), .ZN(new_n979));
  INV_X1    g554(.A(new_n931), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n971), .A4(new_n970), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n974), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n972), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n967), .A2(new_n969), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n980), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n986), .A2(new_n987), .A3(new_n982), .A4(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n989), .A2(new_n982), .A3(new_n971), .A4(new_n970), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT108), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n931), .B1(new_n978), .B2(new_n967), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT43), .B1(new_n972), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n990), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n985), .B1(new_n995), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g571(.A(new_n755), .B(new_n757), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n707), .A2(new_n709), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(G1996), .ZN(new_n999));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n506), .B1(new_n511), .B2(G2105), .ZN(new_n1001));
  INV_X1    g576(.A(new_n501), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n509), .A2(G126), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n467), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n477), .ZN(new_n1008));
  INV_X1    g583(.A(new_n480), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(G40), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n999), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(G1996), .A3(new_n706), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT110), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1011), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n829), .A2(new_n831), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n820), .A2(new_n814), .A3(new_n824), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1012), .B(new_n1014), .C1(new_n1015), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n596), .A2(new_n839), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT109), .Z(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n839), .B2(new_n596), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1019), .B1(new_n1011), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1010), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1027), .B2(G2078), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT124), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1005), .A2(KEYINPUT50), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n512), .A2(new_n1035), .A3(new_n1000), .ZN(new_n1036));
  INV_X1    g611(.A(G40), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n477), .A2(new_n480), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT121), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1010), .B1(new_n1005), .B2(KEYINPUT50), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(new_n1036), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1961), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1027), .A2(KEYINPUT124), .A3(new_n1028), .ZN(new_n1045));
  OR3_X1    g620(.A1(new_n1033), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1024), .B1(new_n1046), .B2(G171), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1031), .ZN(new_n1048));
  INV_X1    g623(.A(G1961), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1043), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1042), .B1(new_n1041), .B2(new_n1036), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n504), .A2(KEYINPUT4), .A3(G138), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n482), .A2(new_n1053), .B1(new_n507), .B2(new_n472), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1054), .A2(new_n467), .B1(new_n505), .B2(new_n503), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1384), .B1(new_n1055), .B2(new_n502), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT45), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1026), .A2(KEYINPUT116), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n1059), .A3(new_n1025), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(new_n1028), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1052), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1048), .B1(new_n1063), .B2(KEYINPUT123), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1052), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1064), .A2(KEYINPUT125), .A3(G301), .A4(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT123), .B1(new_n1044), .B2(new_n1061), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1066), .A2(new_n1068), .A3(G301), .A4(new_n1031), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT125), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1047), .A2(new_n1067), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1056), .B2(new_n1038), .ZN(new_n1075));
  AND4_X1   g650(.A1(new_n1074), .A2(new_n1038), .A3(new_n512), .A4(new_n1000), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n757), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT120), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n757), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1348), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1073), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1348), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1085), .A2(KEYINPUT60), .A3(new_n1080), .A4(new_n1078), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n607), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1038), .A2(new_n512), .A3(new_n1074), .A4(new_n1000), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1996), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1007), .A2(new_n1092), .A3(new_n1038), .A4(new_n1026), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n549), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT122), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1098), .A3(new_n549), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1094), .B2(new_n549), .ZN(new_n1101));
  AOI211_X1 g676(.A(KEYINPUT122), .B(new_n616), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT59), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1081), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1105), .A2(KEYINPUT60), .A3(new_n606), .A4(new_n1085), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n568), .A2(new_n1107), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n943), .A2(new_n1107), .B1(new_n560), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  AND4_X1   g685(.A1(new_n1038), .A2(new_n1007), .A3(new_n1026), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(G1956), .B1(new_n1041), .B2(new_n1036), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NOR4_X1   g688(.A1(new_n560), .A2(KEYINPUT57), .A3(new_n566), .A4(new_n567), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1025), .A2(new_n1026), .A3(new_n1110), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1115), .B(new_n1116), .C1(new_n1117), .C2(G1956), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1113), .A2(new_n1118), .A3(KEYINPUT61), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT61), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1087), .A2(new_n1104), .A3(new_n1106), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1113), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1105), .A2(new_n1085), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1118), .A2(new_n607), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(G301), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1128));
  NOR4_X1   g703(.A1(new_n1033), .A2(new_n1044), .A3(G171), .A4(new_n1045), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1024), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT111), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1041), .A2(new_n696), .A3(new_n1036), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1971), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT113), .ZN(new_n1136));
  INV_X1    g711(.A(G8), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1138));
  NOR3_X1   g713(.A1(G166), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT55), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(KEYINPUT112), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(G303), .B2(G8), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1136), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1138), .ZN(new_n1144));
  NAND3_X1  g719(.A1(G303), .A2(G8), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G166), .A2(new_n1137), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1145), .B(KEYINPUT113), .C1(new_n1146), .C2(new_n1141), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1027), .A2(new_n797), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT111), .A3(new_n1132), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1135), .A2(new_n1148), .A3(new_n1150), .A4(G8), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1153), .B2(new_n1137), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1137), .B1(new_n1056), .B2(new_n1038), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n587), .A2(new_n684), .A3(new_n588), .A4(new_n589), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n586), .A2(new_n518), .ZN(new_n1158));
  INV_X1    g733(.A(G48), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n588), .B1(new_n1159), .B2(new_n529), .ZN(new_n1160));
  OAI21_X1  g735(.A(G1981), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1157), .A2(KEYINPUT49), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT49), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1156), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n924), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1165));
  INV_X1    g740(.A(G1976), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT114), .B1(G288), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT114), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n578), .A2(new_n583), .A3(new_n1168), .A4(G1976), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1155), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT52), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1171), .A2(KEYINPUT115), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1165), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1155), .A2(new_n1167), .A3(new_n1172), .A4(new_n1169), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1164), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1151), .A2(new_n1154), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1060), .A2(new_n726), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1117), .A2(new_n732), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(G168), .ZN(new_n1181));
  OAI21_X1  g756(.A(G8), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n726), .A2(new_n1060), .B1(new_n1117), .B2(new_n732), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1183), .A2(G168), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT51), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1137), .B1(new_n1183), .B2(G168), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT51), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1177), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  AND4_X1   g764(.A1(new_n1072), .A2(new_n1127), .A3(new_n1130), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n611), .A2(G8), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1183), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1151), .A2(new_n1154), .A3(new_n1176), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT117), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT118), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1149), .A2(new_n1132), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1137), .B1(new_n1199), .B2(new_n1131), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1198), .B1(new_n1200), .B2(new_n1150), .ZN(new_n1201));
  AND4_X1   g776(.A1(new_n1198), .A2(new_n1135), .A3(G8), .A4(new_n1150), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1152), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AND4_X1   g778(.A1(KEYINPUT63), .A2(new_n1151), .A3(new_n1176), .A4(new_n1192), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1193), .A2(KEYINPUT117), .A3(new_n1194), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1197), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  OR3_X1    g782(.A1(new_n1164), .A2(G1976), .A3(G288), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1156), .B1(new_n1208), .B2(new_n1157), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1151), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1209), .B1(new_n1210), .B2(new_n1176), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1187), .B1(new_n1186), .B2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1182), .A2(KEYINPUT51), .ZN(new_n1214));
  OAI21_X1  g789(.A(KEYINPUT62), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1185), .A2(new_n1216), .A3(new_n1188), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1177), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1215), .A2(new_n1217), .A3(new_n1128), .A4(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1207), .A2(new_n1211), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1023), .B1(new_n1190), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1011), .A2(new_n1092), .ZN(new_n1222));
  XOR2_X1   g797(.A(new_n1222), .B(KEYINPUT46), .Z(new_n1223));
  AOI21_X1  g798(.A(new_n1015), .B1(new_n997), .B2(new_n885), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  XOR2_X1   g800(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1226));
  XNOR2_X1  g801(.A(new_n1225), .B(new_n1226), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1021), .A2(new_n1015), .ZN(new_n1228));
  XNOR2_X1  g803(.A(new_n1228), .B(KEYINPUT48), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1227), .B1(new_n1019), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1231));
  OAI22_X1  g806(.A1(new_n1231), .A2(new_n1017), .B1(G2067), .B2(new_n755), .ZN(new_n1232));
  AOI21_X1  g807(.A(KEYINPUT126), .B1(new_n1232), .B2(new_n1011), .ZN(new_n1233));
  AND3_X1   g808(.A1(new_n1232), .A2(KEYINPUT126), .A3(new_n1011), .ZN(new_n1234));
  NOR3_X1   g809(.A1(new_n1230), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1221), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g811(.A1(G227), .A2(new_n465), .A3(G401), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1238), .B1(new_n687), .B2(new_n690), .ZN(new_n1239));
  NAND2_X1  g813(.A1(new_n913), .A2(new_n918), .ZN(new_n1240));
  NAND2_X1  g814(.A1(new_n974), .A2(new_n983), .ZN(new_n1241));
  AND3_X1   g815(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(G308));
  NAND3_X1  g816(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(G225));
endmodule


