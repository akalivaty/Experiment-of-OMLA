//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G224), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT0), .B(G128), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT64), .B1(new_n194), .B2(G143), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(G143), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n193), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(G146), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT0), .A4(G128), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT82), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT82), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n208), .B(G125), .C1(new_n201), .C2(new_n204), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n200), .A3(new_n202), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n197), .A2(G146), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n214), .B1(new_n195), .B2(new_n198), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n200), .B2(KEYINPUT1), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n206), .B(new_n213), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT83), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n192), .B1(new_n210), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n217), .B(KEYINPUT83), .ZN(new_n221));
  INV_X1    g035(.A(new_n192), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n207), .A4(new_n209), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n225));
  INV_X1    g039(.A(G107), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G104), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n227), .A2(KEYINPUT3), .B1(new_n228), .B2(G107), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n225), .A2(new_n230), .A3(new_n226), .A4(G104), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(G101), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G116), .ZN(new_n236));
  INV_X1    g050(.A(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n241), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n227), .A2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g060(.A(G101), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n228), .A2(G107), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n231), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT4), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n229), .B2(new_n231), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n234), .B(new_n245), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n226), .A2(G104), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n248), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT80), .A3(G101), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT80), .ZN(new_n256));
  XNOR2_X1  g070(.A(G104), .B(G107), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n247), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n249), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n240), .A2(KEYINPUT5), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n236), .A2(KEYINPUT5), .ZN(new_n261));
  INV_X1    g075(.A(G113), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n260), .A2(new_n263), .B1(new_n240), .B2(new_n242), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n252), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G122), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n252), .A2(new_n265), .A3(new_n267), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(KEYINPUT6), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n272), .A3(new_n268), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n224), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT7), .ZN(new_n275));
  OAI22_X1  g089(.A1(new_n210), .A2(new_n219), .B1(new_n275), .B2(new_n192), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n192), .A2(new_n275), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n221), .A2(new_n207), .A3(new_n209), .A4(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n267), .B(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n265), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n259), .A2(new_n264), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n276), .A2(new_n270), .A3(new_n278), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n190), .B1(new_n274), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n224), .A2(new_n271), .A3(new_n273), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n288), .A2(new_n285), .A3(new_n189), .A4(new_n284), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n188), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(new_n285), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n249), .A2(new_n255), .A3(new_n258), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n200), .A2(new_n202), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n213), .B1(new_n298), .B2(new_n216), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(new_n249), .A3(new_n255), .A4(new_n258), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G134), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G137), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT11), .ZN(new_n304));
  INV_X1    g118(.A(G137), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(G134), .B2(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n302), .A2(KEYINPUT11), .A3(G137), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G131), .ZN(new_n309));
  INV_X1    g123(.A(G131), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n310), .B(new_n303), .C1(new_n306), .C2(new_n307), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(KEYINPUT66), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT81), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n308), .A2(new_n314), .A3(G131), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT12), .B1(new_n301), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n316), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT12), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n297), .A2(new_n300), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n234), .B(new_n205), .C1(new_n251), .C2(new_n250), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT10), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n300), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n312), .A2(new_n315), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n258), .A2(new_n255), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n326), .A2(KEYINPUT10), .A3(new_n294), .A4(new_n249), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n322), .A2(new_n324), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n317), .A2(new_n321), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G140), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n331), .A2(G227), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n324), .A2(new_n327), .ZN(new_n336));
  INV_X1    g150(.A(new_n322), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n315), .B(new_n312), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n329), .A2(new_n333), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n293), .B1(new_n339), .B2(G469), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n317), .A3(new_n321), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n324), .A2(new_n327), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n325), .B1(new_n342), .B2(new_n322), .ZN(new_n343));
  INV_X1    g157(.A(new_n328), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n333), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n292), .A3(new_n285), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT9), .B(G234), .ZN(new_n349));
  OAI21_X1  g163(.A(G221), .B1(new_n349), .B2(G902), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n291), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n353));
  INV_X1    g167(.A(new_n245), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT67), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n305), .B2(G134), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n305), .A2(G134), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n302), .A2(KEYINPUT67), .A3(G137), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G131), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n311), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT68), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n311), .A3(KEYINPUT68), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(new_n294), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n312), .A2(new_n205), .A3(new_n315), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT30), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT65), .B1(new_n201), .B2(new_n204), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT65), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n203), .B(new_n370), .C1(new_n215), .C2(new_n193), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n312), .A2(new_n369), .A3(new_n315), .A4(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT30), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n294), .A2(new_n311), .A3(new_n360), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n354), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n377));
  NOR2_X1   g191(.A1(G237), .A2(G953), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G210), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n377), .B(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT26), .B(G101), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n365), .A2(new_n366), .A3(new_n354), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n376), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n382), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n354), .B1(new_n372), .B2(new_n374), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT28), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n386), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n353), .B1(new_n385), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n391), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n367), .A2(new_n245), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n383), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n394), .B1(KEYINPUT28), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n386), .A2(new_n353), .ZN(new_n398));
  AOI21_X1  g212(.A(G902), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G472), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT32), .ZN(new_n402));
  INV_X1    g216(.A(new_n387), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n372), .A2(new_n374), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n245), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n405), .B2(new_n383), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n386), .B1(new_n406), .B2(new_n394), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n383), .A2(new_n382), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT31), .B1(new_n376), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n373), .B1(new_n365), .B2(new_n366), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n245), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT31), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n382), .A4(new_n383), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G472), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n285), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT71), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n402), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n415), .A2(new_n402), .A3(new_n419), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n401), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G217), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(G234), .B2(new_n285), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT25), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT77), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT76), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT22), .B(G137), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n206), .A2(G140), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT16), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G140), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT73), .B1(new_n436), .B2(G125), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT73), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n206), .A3(G140), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n432), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n435), .B1(new_n440), .B2(new_n434), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G146), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT23), .B1(new_n211), .B2(G119), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n211), .A2(G119), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT74), .ZN(new_n446));
  INV_X1    g260(.A(G110), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n211), .A2(KEYINPUT23), .A3(G119), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n445), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n235), .B2(G128), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n235), .A2(G128), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n451), .A2(new_n448), .A3(new_n447), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT74), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT72), .B1(new_n235), .B2(G128), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT72), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n211), .A3(G119), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n457), .A3(new_n452), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT24), .B(G110), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n449), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n206), .A2(G140), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n433), .A2(new_n462), .A3(new_n194), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n442), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n451), .A2(new_n452), .A3(new_n448), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G110), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n459), .B2(new_n458), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n194), .B(new_n435), .C1(new_n440), .C2(new_n434), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n442), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT75), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n464), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n442), .A2(new_n468), .ZN(new_n472));
  INV_X1    g286(.A(new_n467), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n442), .A2(new_n461), .A3(new_n463), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT75), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n431), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n431), .B1(new_n474), .B2(new_n475), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n426), .B1(new_n480), .B2(new_n285), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n470), .B1(new_n464), .B2(new_n469), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n474), .A2(KEYINPUT75), .A3(new_n475), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n430), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n285), .B(new_n426), .C1(new_n484), .C2(new_n478), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n424), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n424), .A2(G902), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT78), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n480), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n352), .A2(new_n422), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n197), .A2(KEYINPUT85), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(G214), .A3(new_n378), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT85), .B(G143), .ZN(new_n497));
  INV_X1    g311(.A(G237), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n498), .A2(new_n331), .A3(G214), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n496), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT17), .A3(G131), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n442), .A2(new_n468), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G143), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n506), .A2(new_n495), .B1(new_n378), .B2(G214), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n498), .A2(new_n331), .A3(G214), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n505), .A2(G143), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G131), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n496), .B(new_n310), .C1(new_n497), .C2(new_n499), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(KEYINPUT88), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n507), .A2(new_n510), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT88), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n310), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n442), .A2(KEYINPUT89), .A3(new_n468), .A4(new_n501), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n504), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(G113), .B(G122), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(new_n228), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n437), .A2(new_n439), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n433), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT87), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n440), .A2(KEYINPUT86), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n527), .A2(new_n528), .A3(G146), .A4(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n500), .B1(new_n531), .B2(new_n310), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n310), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n496), .B(new_n533), .C1(new_n497), .C2(new_n499), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n526), .B(new_n432), .C1(new_n437), .C2(new_n439), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT86), .B1(new_n524), .B2(new_n433), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n536), .A2(new_n537), .A3(new_n194), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n463), .A2(KEYINPUT87), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n530), .B(new_n535), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n521), .A2(new_n523), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT19), .B1(new_n536), .B2(new_n537), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT19), .B1(new_n433), .B2(new_n462), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(G146), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n513), .A2(new_n442), .A3(new_n516), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n523), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n541), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(G475), .A2(G902), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n494), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n551), .ZN(new_n553));
  AOI211_X1 g367(.A(KEYINPUT20), .B(new_n553), .C1(new_n541), .C2(new_n549), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n521), .A2(new_n540), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n548), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n556), .B2(new_n541), .ZN(new_n557));
  INV_X1    g371(.A(G475), .ZN(new_n558));
  OAI22_X1  g372(.A1(new_n552), .A2(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT90), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI221_X1 g375(.A(KEYINPUT90), .B1(new_n557), .B2(new_n558), .C1(new_n552), .C2(new_n554), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n331), .A2(G952), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(G902), .A3(G953), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT96), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n211), .A2(G143), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n197), .A2(G128), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT92), .B1(new_n574), .B2(new_n576), .ZN(new_n579));
  INV_X1    g393(.A(new_n577), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n573), .B1(new_n580), .B2(KEYINPUT13), .ZN(new_n581));
  OAI211_X1 g395(.A(G134), .B(new_n578), .C1(new_n579), .C2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n574), .A2(new_n580), .A3(new_n302), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  INV_X1    g398(.A(G122), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n584), .B1(new_n585), .B2(G116), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n237), .A2(KEYINPUT91), .A3(G122), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n586), .A2(new_n587), .B1(G116), .B2(new_n585), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(new_n226), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n226), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n582), .B(new_n583), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G134), .B1(new_n573), .B2(new_n577), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n583), .A2(new_n592), .B1(new_n588), .B2(new_n226), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n587), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n594), .A2(KEYINPUT14), .B1(G116), .B2(new_n585), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT14), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n586), .A2(new_n596), .A3(new_n587), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n226), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n593), .B1(new_n598), .B2(KEYINPUT93), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT93), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n600), .B(new_n226), .C1(new_n595), .C2(new_n597), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n591), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n349), .A2(new_n423), .A3(G953), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n591), .B(new_n603), .C1(new_n599), .C2(new_n601), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n602), .A2(KEYINPUT94), .A3(new_n604), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n285), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G478), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(KEYINPUT15), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n612), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n608), .A2(new_n285), .A3(new_n609), .A4(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n613), .A2(KEYINPUT95), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT95), .B1(new_n613), .B2(new_n615), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n563), .A2(new_n572), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n563), .A2(KEYINPUT97), .A3(new_n572), .A4(new_n618), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n493), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT98), .B(G101), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G3));
  NAND2_X1  g439(.A1(new_n415), .A2(new_n285), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G472), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n415), .A2(new_n419), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n629), .A2(new_n491), .A3(new_n351), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n608), .A2(new_n631), .A3(new_n609), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n605), .A2(KEYINPUT33), .A3(new_n607), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(G478), .A3(new_n285), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT99), .B(G478), .Z(new_n635));
  NAND2_X1  g449(.A1(new_n610), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n561), .A2(new_n562), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n290), .A2(new_n572), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n630), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n228), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NOR3_X1   g459(.A1(new_n618), .A2(new_n640), .A3(new_n559), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n630), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  INV_X1    g463(.A(new_n350), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n340), .B2(new_n347), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n431), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT101), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n471), .A2(new_n476), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n489), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n424), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n484), .A2(new_n478), .ZN(new_n661));
  OAI211_X1 g475(.A(KEYINPUT77), .B(new_n425), .C1(new_n661), .C2(G902), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n660), .B1(new_n662), .B2(new_n485), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n651), .B(new_n290), .C1(new_n659), .C2(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(new_n629), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n621), .B2(new_n622), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NAND2_X1  g482(.A1(new_n628), .A2(KEYINPUT32), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n415), .A2(new_n402), .A3(new_n419), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n669), .A2(new_n670), .B1(G472), .B2(new_n400), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n664), .ZN(new_n672));
  INV_X1    g486(.A(new_n559), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n569), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT102), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n566), .B(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n673), .B(new_n678), .C1(new_n616), .C2(new_n617), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  NAND2_X1  g496(.A1(new_n287), .A2(new_n289), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT38), .Z(new_n684));
  NAND3_X1  g498(.A1(new_n487), .A2(new_n187), .A3(new_n658), .ZN(new_n685));
  NOR4_X1   g499(.A1(new_n684), .A2(new_n563), .A3(new_n618), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n678), .B(KEYINPUT39), .Z(new_n687));
  NOR2_X1   g501(.A1(new_n351), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT40), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n386), .B1(new_n412), .B2(new_n383), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n285), .B1(new_n396), .B2(new_n382), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g508(.A(KEYINPUT104), .B(G472), .C1(new_n690), .C2(new_n691), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n421), .B2(new_n420), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT105), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n696), .B(new_n699), .C1(new_n421), .C2(new_n420), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n686), .A2(new_n689), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  INV_X1    g517(.A(new_n678), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n638), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n672), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  NOR2_X1   g521(.A1(new_n671), .A2(new_n491), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n292), .B1(new_n346), .B2(new_n285), .ZN(new_n709));
  AOI211_X1 g523(.A(G469), .B(G902), .C1(new_n341), .C2(new_n345), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n350), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n708), .A2(new_n639), .A3(new_n641), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT106), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n714), .B(new_n716), .ZN(G15));
  NAND3_X1  g531(.A1(new_n708), .A2(new_n646), .A3(new_n713), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NAND3_X1  g533(.A1(new_n711), .A2(new_n290), .A3(new_n350), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n487), .A2(new_n658), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n422), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n621), .B2(new_n622), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n235), .ZN(G21));
  OAI211_X1 g539(.A(new_n409), .B(new_n414), .C1(new_n397), .C2(new_n382), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n626), .A2(G472), .B1(new_n419), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n492), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n290), .B1(new_n616), .B2(new_n617), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n563), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n730), .A3(new_n572), .A4(new_n713), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND2_X1  g546(.A1(new_n726), .A2(new_n419), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n722), .A2(new_n627), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n720), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n705), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n351), .B(KEYINPUT107), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n683), .B2(new_n188), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n287), .A2(KEYINPUT108), .A3(new_n187), .A4(new_n289), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n739), .A2(new_n708), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n705), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n738), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n422), .A2(new_n492), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n743), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(KEYINPUT42), .A3(new_n705), .A4(new_n739), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  NOR2_X1   g566(.A1(new_n745), .A2(new_n679), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n302), .ZN(G36));
  NAND2_X1  g568(.A1(new_n563), .A2(new_n637), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n629), .A2(new_n722), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT44), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(new_n761), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n743), .B(KEYINPUT109), .Z(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(G469), .B1(new_n339), .B2(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(KEYINPUT45), .B2(new_n339), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  OR3_X1    g583(.A1(new_n768), .A2(new_n769), .A3(new_n293), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n768), .B2(new_n293), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n347), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n350), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n687), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n766), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  NOR3_X1   g592(.A1(new_n422), .A2(new_n743), .A3(new_n492), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(KEYINPUT111), .A3(new_n705), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n772), .A2(KEYINPUT47), .A3(new_n350), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT47), .B1(new_n772), .B2(new_n350), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT111), .B1(new_n779), .B2(new_n705), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  INV_X1    g601(.A(new_n677), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n743), .A2(new_n712), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n757), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n701), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n567), .A3(new_n492), .A4(new_n789), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n563), .A2(new_n636), .A3(new_n634), .ZN(new_n793));
  OAI22_X1  g607(.A1(new_n790), .A2(new_n734), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n757), .A2(new_n788), .A3(new_n728), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n684), .A2(new_n188), .A3(new_n713), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT119), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n796), .A2(KEYINPUT50), .A3(new_n798), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n794), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n782), .A2(new_n783), .ZN(new_n804));
  INV_X1    g618(.A(new_n711), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n350), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n765), .A3(new_n796), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n803), .A2(KEYINPUT51), .A3(new_n807), .ZN(new_n808));
  OAI221_X1 g622(.A(new_n564), .B1(new_n792), .B2(new_n638), .C1(new_n795), .C2(new_n720), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n790), .A2(new_n748), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT48), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT48), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n796), .A2(new_n765), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n804), .A2(KEYINPUT118), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n804), .A2(KEYINPUT118), .B1(new_n650), .B2(new_n711), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT51), .B1(new_n819), .B2(new_n803), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT120), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  INV_X1    g636(.A(new_n803), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n822), .B1(new_n823), .B2(new_n818), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n808), .A4(new_n813), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n651), .A2(new_n487), .A3(new_n658), .A4(new_n678), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n563), .A3(new_n729), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n701), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n706), .A3(new_n681), .A4(new_n736), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n701), .A2(new_n829), .B1(new_n672), .B2(new_n705), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n680), .A2(new_n672), .B1(new_n735), .B2(new_n705), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT113), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n831), .A2(KEYINPUT52), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT114), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n834), .A2(KEYINPUT113), .A3(new_n835), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT113), .B1(new_n834), .B2(new_n835), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n845), .A3(new_n838), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n753), .B1(new_n747), .B2(new_n750), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n621), .A2(new_n622), .B1(new_n665), .B2(new_n493), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n613), .A2(new_n615), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n561), .B2(new_n562), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT112), .B1(new_n639), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(KEYINPUT112), .B2(new_n639), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n630), .A2(new_n641), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n848), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n714), .A2(new_n731), .A3(new_n718), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n724), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n739), .A2(new_n705), .A3(new_n727), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n673), .A2(new_n651), .A3(new_n849), .A4(new_n678), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n671), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n722), .A3(new_n744), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n847), .A2(new_n854), .A3(new_n856), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n840), .A2(new_n846), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n842), .A2(new_n843), .A3(new_n841), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT115), .B1(new_n865), .B2(new_n837), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n833), .A2(KEYINPUT52), .A3(new_n836), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n844), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n869), .A3(new_n862), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(KEYINPUT54), .B(new_n864), .C1(new_n871), .C2(new_n863), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n863), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n714), .A2(new_n731), .ZN(new_n874));
  INV_X1    g688(.A(new_n724), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT116), .A4(new_n718), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n855), .B2(new_n724), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n854), .A3(new_n878), .A4(KEYINPUT53), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n847), .A2(new_n860), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n840), .A3(new_n846), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n883));
  NAND3_X1  g697(.A1(new_n873), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n872), .A2(new_n884), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n827), .A2(new_n885), .B1(G952), .B2(G953), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n805), .A2(KEYINPUT49), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n805), .A2(KEYINPUT49), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n637), .A3(new_n888), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n889), .A2(new_n491), .A3(new_n188), .A4(new_n650), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n563), .A3(new_n684), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n886), .B1(new_n701), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n331), .A2(G952), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n844), .A2(new_n867), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n861), .B1(new_n894), .B2(KEYINPUT115), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n895), .B2(new_n869), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n881), .A2(new_n840), .A3(new_n846), .ZN(new_n897));
  OAI211_X1 g711(.A(G210), .B(G902), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n271), .A2(new_n273), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(new_n224), .Z(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n893), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n873), .A2(new_n882), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(KEYINPUT121), .A3(G210), .A4(G902), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n903), .A2(KEYINPUT56), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n904), .A2(new_n910), .ZN(G51));
  XNOR2_X1  g725(.A(new_n293), .B(KEYINPUT57), .ZN(new_n912));
  INV_X1    g726(.A(new_n883), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n896), .A2(new_n897), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n883), .B1(new_n873), .B2(new_n882), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n346), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n285), .B1(new_n873), .B2(new_n882), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n768), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n893), .B1(new_n917), .B2(new_n919), .ZN(G54));
  AND2_X1   g734(.A1(KEYINPUT58), .A2(G475), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n907), .A2(G902), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n550), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT122), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n893), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n918), .A2(new_n926), .A3(new_n550), .A4(new_n921), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(G60));
  AND2_X1   g742(.A1(new_n632), .A2(new_n633), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT59), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n929), .B(new_n931), .C1(new_n914), .C2(new_n915), .ZN(new_n932));
  INV_X1    g746(.A(new_n893), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n885), .B2(new_n931), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n873), .B2(new_n882), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(new_n480), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n656), .A2(new_n657), .ZN(new_n941));
  INV_X1    g755(.A(new_n938), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n941), .B(new_n942), .C1(new_n896), .C2(new_n897), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n940), .A2(KEYINPUT61), .A3(new_n933), .A4(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n943), .B(new_n933), .C1(new_n939), .C2(new_n480), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n947), .ZN(G66));
  OAI21_X1  g762(.A(G953), .B1(new_n570), .B2(new_n191), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n854), .A2(new_n856), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n951), .B2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n901), .B1(G898), .B2(new_n331), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT123), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n952), .B(new_n954), .ZN(G69));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n835), .A2(new_n706), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n774), .A2(new_n708), .A3(new_n730), .ZN(new_n958));
  AND4_X1   g772(.A1(new_n786), .A2(new_n847), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n777), .A2(new_n331), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n368), .A2(new_n375), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n542), .A2(new_n544), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n961), .B(new_n962), .Z(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(G900), .B2(G953), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n956), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n852), .A2(new_n688), .A3(new_n749), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n784), .B2(new_n785), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n957), .B2(new_n702), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n957), .A2(new_n969), .A3(new_n702), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n957), .A2(new_n702), .A3(KEYINPUT124), .A4(new_n969), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n971), .B(new_n976), .C1(new_n775), .C2(new_n776), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n331), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT125), .B1(new_n978), .B2(new_n964), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n980), .B(new_n963), .C1(new_n977), .C2(new_n331), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n966), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n331), .B1(G227), .B2(G900), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n966), .B(new_n985), .C1(new_n979), .C2(new_n981), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n977), .B2(new_n950), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n893), .B1(new_n990), .B2(new_n690), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n959), .B(new_n951), .C1(new_n776), .C2(new_n775), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n989), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n385), .ZN(new_n994));
  INV_X1    g808(.A(new_n385), .ZN(new_n995));
  INV_X1    g809(.A(new_n690), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n996), .A3(new_n989), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n864), .B(new_n998), .C1(new_n871), .C2(new_n863), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n991), .A2(new_n994), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(KEYINPUT127), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n991), .A2(new_n994), .A3(new_n1002), .A4(new_n999), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G57));
endmodule


