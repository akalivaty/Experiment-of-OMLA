//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XOR2_X1   g044(.A(KEYINPUT66), .B(G2105), .Z(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(G137), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT67), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n460), .A3(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(KEYINPUT68), .B1(new_n477), .B2(G101), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  INV_X1    g054(.A(G101), .ZN(new_n480));
  AOI211_X1 g055(.A(new_n479), .B(new_n480), .C1(new_n474), .C2(new_n476), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n469), .B(new_n472), .C1(new_n478), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n460), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n463), .B1(new_n485), .B2(new_n486), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n489), .B1(new_n492), .B2(G124), .ZN(G162));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n496), .B2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT71), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n471), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n461), .B(new_n462), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n470), .A2(new_n510), .A3(G138), .A4(new_n471), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n504), .B1(new_n509), .B2(new_n511), .ZN(G164));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT72), .B1(new_n513), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT6), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(new_n517), .B1(new_n513), .B2(G651), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n518), .A2(G50), .A3(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(new_n517), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n513), .A2(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n518), .A2(KEYINPUT74), .A3(new_n525), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G88), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n516), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n520), .A2(new_n532), .A3(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  NAND3_X1  g111(.A1(new_n518), .A2(G51), .A3(G543), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n541), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n525), .A2(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G89), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n530), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n516), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n528), .A2(G90), .A3(new_n529), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n518), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G52), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n550), .A2(KEYINPUT75), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(KEYINPUT75), .B1(new_n550), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND2_X1  g131(.A1(new_n531), .A2(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n523), .A2(new_n524), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n551), .A2(G43), .B1(new_n561), .B2(G651), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  AOI22_X1  g143(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n516), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n528), .A2(G91), .A3(new_n529), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n521), .A2(G53), .A3(G543), .A4(new_n522), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n518), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n574), .B1(new_n573), .B2(new_n576), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n570), .B(new_n571), .C1(new_n578), .C2(new_n579), .ZN(G299));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n546), .B(new_n581), .ZN(G286));
  OR2_X1    g157(.A1(new_n525), .A2(G74), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n551), .A2(G49), .B1(G651), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n528), .A2(G87), .A3(new_n529), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G288));
  NAND3_X1  g161(.A1(new_n528), .A2(G86), .A3(new_n529), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n521), .A2(G48), .A3(G543), .A4(new_n522), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n518), .A2(KEYINPUT79), .A3(G48), .A4(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n523), .B2(new_n524), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n594), .B2(new_n595), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n587), .A2(new_n592), .A3(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n551), .A2(G47), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI221_X1 g179(.A(new_n602), .B1(new_n516), .B2(new_n603), .C1(new_n530), .C2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n516), .B1(new_n607), .B2(KEYINPUT80), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(KEYINPUT80), .B2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n551), .A2(G54), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n530), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n611), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(G868), .B2(new_n616), .ZN(G284));
  OAI21_X1  g192(.A(new_n606), .B1(G868), .B2(new_n616), .ZN(G321));
  NOR2_X1   g193(.A1(G299), .A2(G868), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n546), .B(KEYINPUT77), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  XOR2_X1   g196(.A(G280), .B(KEYINPUT81), .Z(G297));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n557), .A2(new_n562), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n616), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n629), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n492), .A2(G123), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n470), .A2(G111), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n633), .B2(KEYINPUT83), .ZN(new_n636));
  INV_X1    g211(.A(new_n487), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n634), .A2(new_n636), .B1(new_n637), .B2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT84), .Z(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2096), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n477), .A2(new_n471), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2100), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(new_n642), .A3(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT86), .B(KEYINPUT14), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1341), .B(G1348), .Z(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  OR2_X1    g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(G401));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT87), .Z(new_n667));
  XOR2_X1   g242(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n667), .B2(new_n670), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(new_n670), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n667), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n672), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n686), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT20), .Z(new_n690));
  AOI211_X1 g265(.A(new_n688), .B(new_n690), .C1(new_n683), .C2(new_n687), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1981), .B(G1986), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT89), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n693), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G22), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1971), .ZN(new_n703));
  MUX2_X1   g278(.A(G23), .B(G288), .S(G16), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT92), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G6), .B(G305), .S(G16), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT91), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT32), .B(G1981), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT34), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  OAI221_X1 g293(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n719));
  INV_X1    g294(.A(G131), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n487), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n492), .B2(G119), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n718), .B1(new_n722), .B2(new_n717), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XOR2_X1   g299(.A(new_n723), .B(new_n724), .Z(new_n725));
  OR2_X1    g300(.A1(G290), .A2(KEYINPUT90), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n700), .B1(G290), .B2(KEYINPUT90), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n726), .A2(new_n727), .B1(new_n700), .B2(G24), .ZN(new_n728));
  INV_X1    g303(.A(G1986), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT93), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(KEYINPUT36), .ZN(new_n733));
  NOR4_X1   g308(.A1(new_n725), .A2(new_n730), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n715), .A2(new_n716), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(KEYINPUT36), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n736), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n715), .A2(new_n738), .A3(new_n716), .A4(new_n734), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n717), .A2(G35), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G162), .B2(new_n717), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT29), .Z(new_n742));
  INV_X1    g317(.A(G2090), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n700), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G299), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n700), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT102), .B(G1956), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n744), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT103), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n717), .A2(G32), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n492), .A2(G129), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT26), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n477), .A2(G105), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n758), .B(new_n759), .C1(new_n637), .C2(G141), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n755), .B1(new_n762), .B2(new_n717), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT27), .B(G1996), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G164), .A2(new_n717), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G27), .B2(new_n717), .ZN(new_n767));
  INV_X1    g342(.A(G2078), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G28), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT30), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n770), .B2(KEYINPUT30), .ZN(new_n772));
  OR2_X1    g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  NAND2_X1  g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT24), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n717), .B1(new_n778), .B2(G34), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(G34), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n779), .B2(KEYINPUT99), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n482), .A2(new_n717), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n776), .B1(new_n768), .B2(new_n767), .C1(new_n777), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n765), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G168), .A2(new_n700), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n700), .B2(G21), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI22_X1  g363(.A1(new_n640), .A2(new_n717), .B1(G1966), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n783), .A2(new_n777), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT100), .Z(new_n791));
  NOR2_X1   g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n742), .A2(new_n743), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n700), .A2(G19), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n563), .B2(new_n700), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1341), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G1966), .B2(new_n788), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n785), .A2(new_n792), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n700), .A2(G5), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G171), .B2(new_n700), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1961), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n717), .A2(G26), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT28), .ZN(new_n803));
  INV_X1    g378(.A(G140), .ZN(new_n804));
  NOR2_X1   g379(.A1(G104), .A2(G2105), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT95), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(new_n470), .B2(G116), .ZN(new_n807));
  OAI22_X1  g382(.A1(new_n487), .A2(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n492), .B2(G128), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n803), .B1(new_n809), .B2(new_n717), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2067), .ZN(new_n811));
  NOR2_X1   g386(.A1(G29), .A2(G33), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT96), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G139), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n487), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n470), .B1(new_n820), .B2(KEYINPUT98), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(KEYINPUT98), .B2(new_n820), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n813), .B1(new_n823), .B2(G29), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n811), .B1(new_n824), .B2(G2072), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n700), .A2(G4), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n616), .B2(new_n700), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT94), .B(G1348), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n825), .B(new_n829), .C1(G2072), .C2(new_n824), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n798), .A2(new_n801), .A3(new_n830), .ZN(new_n831));
  AND4_X1   g406(.A1(new_n737), .A2(new_n739), .A3(new_n754), .A4(new_n831), .ZN(G311));
  NAND4_X1  g407(.A1(new_n737), .A2(new_n739), .A3(new_n754), .A4(new_n831), .ZN(G150));
  NAND2_X1  g408(.A1(new_n551), .A2(G55), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI221_X1 g411(.A(new_n834), .B1(new_n516), .B2(new_n835), .C1(new_n530), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n616), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT104), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n625), .B(new_n837), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n844), .A2(new_n845), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n839), .B1(new_n848), .B2(new_n849), .ZN(G145));
  XNOR2_X1  g425(.A(new_n722), .B(new_n645), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n823), .A2(new_n762), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n819), .A2(new_n822), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n761), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n852), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n492), .A2(G130), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT106), .ZN(new_n859));
  OAI221_X1 g434(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n470), .C2(G118), .ZN(new_n860));
  INV_X1    g435(.A(G142), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n487), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n509), .A2(new_n511), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n460), .B1(KEYINPUT71), .B2(new_n498), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n496), .A2(G114), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n494), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n501), .B1(new_n465), .B2(new_n466), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT105), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n864), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n809), .B(new_n872), .Z(new_n873));
  OR2_X1    g448(.A1(new_n863), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n863), .A2(new_n873), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n853), .A2(new_n855), .A3(new_n852), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n857), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  INV_X1    g453(.A(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n856), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n640), .A2(G160), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n639), .B(KEYINPUT84), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n482), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G162), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(G162), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n881), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n877), .A2(new_n880), .A3(new_n888), .A4(new_n887), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(G395));
  XNOR2_X1  g470(.A(G303), .B(G305), .ZN(new_n896));
  XNOR2_X1  g471(.A(G290), .B(G288), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT109), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n629), .B(new_n843), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n748), .A2(new_n616), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n748), .A2(new_n616), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n628), .A2(G299), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n906), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n909), .A2(new_n910), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n906), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n905), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n902), .B(new_n904), .C1(new_n915), .C2(new_n917), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n837), .A2(new_n626), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(G295));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n925), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  NAND2_X1  g503(.A1(G171), .A2(new_n620), .ZN(new_n929));
  NAND2_X1  g504(.A1(G301), .A2(new_n546), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n843), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n843), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n916), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n563), .B(new_n837), .ZN(new_n934));
  INV_X1    g509(.A(new_n930), .ZN(new_n935));
  NOR2_X1   g510(.A1(G286), .A2(G301), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n843), .A2(new_n929), .A3(new_n930), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n937), .A2(new_n911), .A3(new_n938), .A4(new_n913), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n898), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n891), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n933), .A2(new_n939), .A3(new_n898), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n898), .B1(new_n933), .B2(new_n939), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT110), .B1(new_n948), .B2(G37), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n942), .A2(new_n891), .A3(new_n945), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n928), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n944), .A2(new_n945), .A3(new_n949), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n948), .A2(G37), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n954), .A2(KEYINPUT43), .B1(new_n955), .B2(new_n947), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n953), .B1(new_n956), .B2(new_n928), .ZN(G397));
  INV_X1    g532(.A(G1996), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n761), .B(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n809), .B(G2067), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n722), .B(new_n724), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(G290), .B(new_n729), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n872), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n477), .A2(G101), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n479), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n477), .A2(KEYINPUT68), .A3(G101), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n973), .A2(G40), .A3(new_n469), .A4(new_n472), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n965), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n872), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n482), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n968), .B1(G164), .B2(G1384), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1971), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n872), .A2(new_n984), .A3(new_n966), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(KEYINPUT111), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n498), .A2(KEYINPUT71), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n867), .A2(new_n988), .A3(G2105), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n989), .A2(new_n495), .B1(new_n471), .B2(new_n502), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n509), .A2(new_n511), .B1(new_n990), .B2(KEYINPUT105), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n991), .B2(new_n870), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n993), .A3(new_n984), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n979), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n983), .B1(new_n996), .B2(G2090), .ZN(new_n997));
  NAND2_X1  g572(.A1(G303), .A2(G8), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n1000), .A3(G8), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT78), .B1(new_n559), .B2(new_n593), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n596), .A3(new_n598), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1005), .A2(G651), .B1(new_n590), .B2(new_n591), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1006), .B2(new_n587), .ZN(new_n1007));
  AND4_X1   g582(.A1(new_n1003), .A2(new_n587), .A3(new_n592), .A4(new_n600), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n967), .A2(new_n974), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G305), .A2(G1981), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1006), .A2(new_n1003), .A3(new_n587), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(KEYINPUT49), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n584), .A2(G1976), .A3(new_n585), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1017), .B(G8), .C1(new_n967), .C2(new_n974), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT52), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n992), .A2(new_n979), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(G8), .A4(new_n1017), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1016), .A2(new_n1019), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1012), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G288), .A2(G1976), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1008), .B1(new_n1016), .B2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1001), .A2(new_n1024), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n995), .A2(new_n777), .A3(new_n979), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT45), .B1(new_n872), .B2(new_n966), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n974), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT113), .B(new_n979), .C1(new_n992), .C2(KEYINPUT45), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n864), .A2(new_n990), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n995), .A2(KEYINPUT114), .A3(new_n777), .A4(new_n979), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1031), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(G8), .A3(new_n620), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT63), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1024), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1001), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n997), .A2(G8), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1044), .B(new_n1047), .C1(new_n1000), .C2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n998), .B(KEYINPUT55), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1036), .A2(new_n984), .A3(new_n966), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n979), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n984), .B1(new_n872), .B2(new_n966), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1052), .A2(G2090), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n982), .B2(new_n981), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1050), .B1(new_n1055), .B2(new_n1011), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1023), .A2(new_n1019), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1057), .A2(KEYINPUT112), .A3(new_n1016), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT112), .B1(new_n1057), .B2(new_n1016), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1001), .B(new_n1056), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1045), .B1(new_n1060), .B2(new_n1043), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1028), .B1(new_n1049), .B2(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n469), .A2(G40), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n472), .B1(new_n478), .B2(new_n481), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(KEYINPUT122), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n973), .B2(new_n472), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT123), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n973), .A2(new_n1066), .A3(new_n472), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(KEYINPUT122), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1063), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n969), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT124), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1068), .A2(new_n969), .A3(new_n1075), .A4(new_n1072), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G2078), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n977), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1961), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n996), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1077), .B1(new_n981), .B2(G2078), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(new_n1082), .A3(G301), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n974), .B1(new_n987), .B2(new_n994), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1085), .B2(G1961), .ZN(new_n1086));
  AND4_X1   g661(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .A4(new_n1078), .ZN(new_n1087));
  OAI21_X1  g662(.A(G171), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT125), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1093), .A3(new_n1090), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n573), .B2(new_n576), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1096), .A2(new_n570), .A3(new_n571), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n1101));
  INV_X1    g676(.A(new_n579), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n577), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n571), .A2(new_n570), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1101), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT115), .B1(new_n1106), .B2(new_n1097), .ZN(new_n1107));
  INV_X1    g682(.A(G1956), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n977), .A2(new_n979), .A3(new_n980), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1100), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n828), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n995), .B2(new_n979), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1022), .A2(G2067), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1098), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n616), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1113), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT116), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1122), .B(new_n1113), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT117), .B(new_n1125), .C1(new_n967), .C2(new_n974), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n977), .A2(new_n958), .A3(new_n979), .A4(new_n980), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT117), .B1(new_n1022), .B2(new_n1125), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n563), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT118), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1132), .B(new_n563), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(KEYINPUT59), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1135), .B(new_n563), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1131), .A2(KEYINPUT119), .A3(KEYINPUT59), .A4(new_n1133), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1143));
  OAI221_X1 g718(.A(KEYINPUT60), .B1(G2067), .B2(new_n1022), .C1(new_n1085), .C2(new_n1114), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n616), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1117), .A2(KEYINPUT60), .A3(new_n628), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1113), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1148));
  INV_X1    g723(.A(new_n1118), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1098), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1124), .B1(new_n1141), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1095), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT114), .B1(new_n1085), .B2(new_n777), .ZN(new_n1156));
  OAI21_X1  g731(.A(G8), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n546), .A2(G8), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT51), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1158), .B2(KEYINPUT121), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(G8), .B(new_n1160), .C1(new_n1042), .C2(new_n546), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1158), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1042), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1080), .A2(new_n1082), .A3(KEYINPUT126), .A4(new_n1083), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1170), .A2(G171), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1090), .B1(new_n1173), .B2(G301), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1060), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1167), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1062), .B1(new_n1154), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1167), .A2(KEYINPUT62), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1060), .A2(new_n1088), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1166), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1180), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1179), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n976), .B1(new_n1177), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n975), .A2(new_n958), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT46), .Z(new_n1187));
  INV_X1    g762(.A(new_n975), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1188), .B1(new_n960), .B2(new_n762), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT47), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1188), .A2(G290), .A3(G1986), .ZN(new_n1192));
  XNOR2_X1  g767(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1194), .B1(new_n963), .B2(new_n1188), .ZN(new_n1195));
  AND4_X1   g770(.A1(new_n724), .A2(new_n959), .A3(new_n722), .A4(new_n960), .ZN(new_n1196));
  INV_X1    g771(.A(G2067), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1196), .B1(new_n1197), .B2(new_n809), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1195), .B1(new_n1198), .B2(new_n1188), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1191), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1185), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g776(.A(G319), .ZN(new_n1203));
  NOR3_X1   g777(.A1(G401), .A2(G227), .A3(new_n1203), .ZN(new_n1204));
  AND2_X1   g778(.A1(new_n698), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n893), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n1206), .A2(new_n956), .ZN(G308));
  OR2_X1    g781(.A1(new_n1206), .A2(new_n956), .ZN(G225));
endmodule


