//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  INV_X1    g0012(.A(G13), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n212), .B1(new_n205), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g0014(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n215));
  AND2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n206), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT65), .Z(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n211), .B1(new_n218), .B2(new_n219), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n246), .A2(G50), .B1(G20), .B2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n248), .B1(new_n251), .B2(new_n202), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n214), .A2(new_n215), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT11), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n213), .A2(new_n206), .A3(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n247), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n257), .B(KEYINPUT12), .Z(new_n258));
  NOR2_X1   g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n252), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n214), .A2(new_n215), .A3(new_n253), .ZN(new_n261));
  INV_X1    g0061(.A(new_n256), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n205), .A2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G68), .A3(new_n265), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n259), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT13), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n249), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n205), .A2(new_n213), .ZN(new_n273));
  NAND3_X1  g0073(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G274), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n277), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(G238), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT69), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n249), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(G1698), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n292), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n286), .A2(new_n291), .ZN(new_n294));
  AND4_X1   g0094(.A1(KEYINPUT74), .A2(new_n294), .A3(G232), .A4(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n286), .B2(new_n291), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT74), .B1(new_n297), .B2(G232), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT75), .B(new_n293), .C1(new_n295), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n214), .A2(new_n215), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n249), .B2(new_n271), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n294), .A2(G232), .A3(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT74), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n297), .A2(KEYINPUT74), .A3(G232), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT75), .B1(new_n308), .B2(new_n293), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n269), .B(new_n283), .C1(new_n303), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT77), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n293), .B1(new_n295), .B2(new_n298), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(new_n302), .A3(new_n299), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT77), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n269), .A4(new_n283), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n283), .B1(new_n303), .B2(new_n309), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G179), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT78), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n319), .B2(KEYINPUT13), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT78), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n311), .A3(new_n325), .A4(new_n317), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n320), .B2(new_n310), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n268), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n286), .A2(new_n291), .ZN(new_n333));
  AOI22_X1  g0133(.A1(G238), .A2(new_n297), .B1(new_n333), .B2(G107), .ZN(new_n334));
  INV_X1    g0134(.A(G232), .ZN(new_n335));
  INV_X1    g0135(.A(new_n292), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n302), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n279), .B1(G244), .B2(new_n282), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n323), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n265), .A2(G77), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n264), .A2(new_n342), .B1(new_n202), .B2(new_n256), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT8), .B(G58), .Z(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n246), .B1(G20), .B2(G77), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT71), .A3(new_n250), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT71), .B1(new_n347), .B2(new_n250), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n254), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n339), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n337), .B2(new_n302), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n340), .B(new_n352), .C1(G169), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n338), .A2(G190), .A3(new_n339), .ZN(new_n356));
  INV_X1    g0156(.A(new_n352), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n354), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n355), .A2(new_n359), .A3(KEYINPUT72), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT72), .B1(new_n355), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT7), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n286), .A2(new_n291), .A3(new_n363), .A4(new_n206), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n290), .A2(new_n206), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT79), .B(G33), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n287), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n364), .B(G68), .C1(new_n363), .C2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(G58), .B(G68), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(G20), .B1(G159), .B2(new_n246), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n206), .B(new_n288), .C1(new_n366), .C2(new_n287), .ZN(new_n374));
  OAI21_X1  g0174(.A(G68), .B1(new_n374), .B2(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n249), .A2(KEYINPUT79), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G33), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n285), .B1(new_n379), .B2(KEYINPUT3), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n363), .B1(new_n380), .B2(new_n206), .ZN(new_n381));
  OAI211_X1 g0181(.A(KEYINPUT16), .B(new_n370), .C1(new_n375), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n373), .A2(new_n254), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT70), .A2(G58), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT8), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n384), .B(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n205), .B2(G20), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n264), .A2(new_n387), .B1(new_n256), .B2(new_n386), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n288), .B1(new_n366), .B2(new_n287), .ZN(new_n389));
  NOR2_X1   g0189(.A1(G223), .A2(G1698), .ZN(new_n390));
  INV_X1    g0190(.A(G226), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(G1698), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G87), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n301), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n275), .A2(G232), .A3(new_n280), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n278), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(G169), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n392), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n380), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n394), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n302), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n397), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(G179), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n383), .A2(new_n388), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT18), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n403), .A3(G190), .ZN(new_n407));
  OAI21_X1  g0207(.A(G200), .B1(new_n395), .B2(new_n397), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n383), .A2(new_n388), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT17), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n278), .B1(new_n281), .B2(new_n391), .ZN(new_n411));
  AOI22_X1  g0211(.A1(G223), .A2(new_n297), .B1(new_n333), .B2(G77), .ZN(new_n412));
  INV_X1    g0212(.A(G222), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n336), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n414), .B2(new_n302), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n415), .A2(new_n323), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n246), .A2(G150), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n417), .B1(new_n206), .B2(new_n201), .C1(new_n386), .C2(new_n251), .ZN(new_n418));
  INV_X1    g0218(.A(G50), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n418), .A2(new_n254), .B1(new_n419), .B2(new_n256), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n264), .A2(G50), .A3(new_n265), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n415), .B2(G169), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT73), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n425), .A3(KEYINPUT9), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n425), .A2(KEYINPUT9), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(KEYINPUT9), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n420), .A2(new_n421), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n415), .A2(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n415), .A2(new_n358), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT10), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n433), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT10), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n431), .A4(new_n430), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n424), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n362), .A2(new_n406), .A3(new_n410), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n320), .A2(G190), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n267), .B1(new_n318), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n320), .A2(new_n310), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G200), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n358), .B1(new_n320), .B2(new_n310), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT76), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n442), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n332), .A2(new_n440), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT82), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n294), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n453));
  INV_X1    g0253(.A(G283), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n249), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n294), .A2(G250), .A3(G1698), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n287), .B1(new_n376), .B2(new_n378), .ZN(new_n459));
  OAI211_X1 g0259(.A(G244), .B(new_n296), .C1(new_n459), .C2(new_n285), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT4), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n302), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n205), .A2(G45), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT5), .B(G41), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n275), .A2(G274), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n465), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n275), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n470), .A2(G257), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n463), .A2(G190), .A3(new_n467), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n262), .A2(G97), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n249), .A2(G1), .ZN(new_n476));
  OR3_X1    g0276(.A1(new_n254), .A2(new_n256), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT6), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT6), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G97), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(KEYINPUT80), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT80), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G107), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n481), .A2(new_n483), .A3(new_n485), .A4(new_n487), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n206), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n202), .A2(G20), .A3(G33), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT81), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND4_X1   g0293(.A1(new_n481), .A2(new_n483), .A3(new_n485), .A4(new_n487), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n481), .A2(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n495));
  OAI21_X1  g0295(.A(G20), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT81), .ZN(new_n497));
  INV_X1    g0297(.A(new_n492), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n364), .B(G107), .C1(new_n363), .C2(new_n367), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n493), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n479), .B1(new_n501), .B2(new_n254), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n473), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n455), .B1(new_n297), .B2(G250), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n460), .A2(new_n461), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(new_n453), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n471), .B1(new_n506), .B2(new_n302), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n358), .B1(new_n507), .B2(new_n467), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n452), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n463), .A2(new_n467), .A3(new_n472), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G200), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n511), .A2(KEYINPUT82), .A3(new_n502), .A4(new_n473), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n502), .A2(KEYINPUT83), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n502), .A2(KEYINPUT83), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n510), .A2(new_n323), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n328), .B1(new_n507), .B2(new_n467), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n389), .A2(new_n206), .A3(G68), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT19), .B1(new_n250), .B2(G97), .ZN(new_n520));
  NAND3_X1  g0320(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n206), .ZN(new_n522));
  INV_X1    g0322(.A(G87), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(new_n478), .A3(new_n480), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n261), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n263), .A2(new_n476), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n347), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n347), .A2(new_n262), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G250), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n464), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n464), .A2(G274), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n275), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n296), .A2(G238), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT84), .B1(new_n380), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n389), .A2(G244), .A3(G1698), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT84), .ZN(new_n541));
  INV_X1    g0341(.A(new_n538), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n389), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n379), .A2(G116), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n539), .A2(new_n540), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n537), .B1(new_n545), .B2(new_n302), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n532), .B1(new_n546), .B2(G169), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI211_X1 g0348(.A(G179), .B(new_n537), .C1(new_n545), .C2(new_n302), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n528), .A2(G87), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n527), .A2(new_n551), .A3(new_n531), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(G190), .B2(new_n546), .ZN(new_n553));
  OR2_X1    g0353(.A1(new_n546), .A2(new_n358), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n548), .A2(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n513), .A2(new_n518), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G270), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n467), .B1(new_n469), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G257), .B(new_n296), .C1(new_n459), .C2(new_n285), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT85), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n389), .A2(KEYINPUT85), .A3(G257), .A4(new_n296), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n286), .A2(new_n291), .A3(G303), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G264), .A2(G1698), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n380), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n558), .B1(new_n568), .B2(new_n302), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n256), .A2(G116), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n477), .B2(G116), .ZN(new_n571));
  AOI21_X1  g0371(.A(G20), .B1(G33), .B2(G283), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n249), .A2(G97), .ZN(new_n573));
  INV_X1    g0373(.A(G116), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n572), .A2(new_n573), .B1(G20), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n254), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n254), .A2(new_n575), .A3(new_n577), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n579), .A2(new_n580), .B1(KEYINPUT86), .B2(KEYINPUT20), .ZN(new_n581));
  OAI21_X1  g0381(.A(G169), .B1(new_n571), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT87), .B1(new_n569), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT21), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT21), .ZN(new_n585));
  OAI211_X1 g0385(.A(KEYINPUT87), .B(new_n585), .C1(new_n569), .C2(new_n582), .ZN(new_n586));
  INV_X1    g0386(.A(new_n558), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n566), .B1(new_n561), .B2(new_n562), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n587), .B(G179), .C1(new_n588), .C2(new_n301), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n571), .A2(new_n581), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n584), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G264), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n467), .B1(new_n469), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT90), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n533), .A2(G1698), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n380), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n389), .A2(G257), .A3(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n389), .A2(KEYINPUT90), .A3(new_n596), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n379), .A2(G294), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n594), .B1(new_n602), .B2(new_n302), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n323), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(G169), .B2(new_n603), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT24), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n206), .B(G87), .C1(new_n459), .C2(new_n285), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT88), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT88), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n389), .A2(new_n609), .A3(new_n206), .A4(G87), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(KEYINPUT22), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT89), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT22), .ZN(new_n613));
  AOI211_X1 g0413(.A(G20), .B(new_n523), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n294), .B(new_n614), .C1(new_n612), .C2(new_n613), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n480), .A2(G20), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT23), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n617), .B(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n544), .B2(G20), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n606), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  AOI211_X1 g0422(.A(KEYINPUT24), .B(new_n620), .C1(new_n611), .C2(new_n615), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n254), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT25), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n262), .B2(G107), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n480), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n528), .A2(G107), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n605), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n603), .A2(new_n358), .ZN(new_n631));
  INV_X1    g0431(.A(G190), .ZN(new_n632));
  AOI211_X1 g0432(.A(new_n632), .B(new_n594), .C1(new_n602), .C2(new_n302), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n624), .A2(new_n634), .A3(new_n628), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n587), .B1(new_n588), .B2(new_n301), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G200), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n637), .B(new_n590), .C1(new_n632), .C2(new_n636), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n592), .A2(new_n630), .A3(new_n635), .A4(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n451), .A2(new_n556), .A3(new_n639), .ZN(G372));
  NOR2_X1   g0440(.A1(new_n449), .A2(new_n355), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n330), .B1(new_n443), .B2(G169), .ZN(new_n642));
  AOI211_X1 g0442(.A(KEYINPUT14), .B(new_n328), .C1(new_n320), .C2(new_n310), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n322), .A2(new_n326), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n267), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n410), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n406), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n434), .A2(new_n437), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n424), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n547), .A2(new_n549), .ZN(new_n651));
  INV_X1    g0451(.A(new_n502), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n516), .B2(new_n517), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n546), .A2(G190), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n527), .A2(new_n551), .A3(new_n531), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n546), .A2(new_n358), .ZN(new_n657));
  OAI22_X1  g0457(.A1(new_n656), .A2(new_n657), .B1(new_n547), .B2(new_n549), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n651), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT26), .B1(new_n518), .B2(new_n658), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n584), .A2(new_n586), .A3(new_n591), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n635), .B1(new_n663), .B2(new_n629), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n661), .B(new_n662), .C1(new_n556), .C2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n650), .B1(new_n451), .B2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G343), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT91), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n590), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n663), .B(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(new_n638), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n629), .A2(new_n674), .ZN(new_n679));
  INV_X1    g0479(.A(new_n674), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n616), .A2(new_n621), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT24), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n616), .A2(new_n606), .A3(new_n621), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n261), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n628), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n686), .A2(new_n635), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n679), .B1(new_n687), .B2(new_n629), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n678), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n663), .A2(new_n674), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n629), .B2(new_n674), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n209), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n524), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n219), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n635), .A2(new_n638), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n702), .A2(new_n663), .A3(new_n629), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n513), .A2(new_n518), .A3(new_n555), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(new_n674), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n546), .A2(new_n603), .ZN(new_n706));
  INV_X1    g0506(.A(new_n589), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n707), .A4(new_n507), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n507), .A2(new_n546), .A3(new_n603), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n589), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n546), .A2(G179), .ZN(new_n712));
  INV_X1    g0512(.A(new_n603), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n510), .A3(new_n636), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n708), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT31), .B1(new_n715), .B2(new_n680), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT92), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n680), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n705), .A2(new_n718), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n502), .B(KEYINPUT83), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n510), .A2(G169), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n323), .B2(new_n510), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n555), .A2(new_n728), .A3(new_n660), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT26), .B1(new_n653), .B2(new_n658), .ZN(new_n732));
  INV_X1    g0532(.A(new_n651), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT93), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n592), .A2(new_n630), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n509), .A2(new_n512), .B1(new_n728), .B2(new_n730), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n737), .A2(new_n738), .A3(new_n555), .A4(new_n635), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT93), .A4(new_n733), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT29), .A3(new_n674), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n664), .A2(new_n556), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n555), .A2(new_n660), .A3(new_n730), .A4(new_n652), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n662), .A2(new_n733), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n674), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n742), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n727), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n701), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR2_X1   g0552(.A1(new_n213), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n205), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n696), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n678), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G330), .ZN(new_n759));
  INV_X1    g0559(.A(new_n677), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OR3_X1    g0563(.A1(new_n763), .A2(KEYINPUT95), .A3(G20), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT95), .B1(new_n763), .B2(G20), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n677), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n216), .B1(G20), .B2(new_n328), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(G20), .A2(G179), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT96), .Z(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n632), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G58), .A2(new_n774), .B1(new_n776), .B2(G77), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT97), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n206), .A2(G179), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n779), .A2(new_n632), .A3(G200), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n294), .B1(new_n523), .B2(new_n780), .C1(new_n480), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n775), .A2(new_n358), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G68), .B2(new_n783), .ZN(new_n784));
  OR3_X1    g0584(.A1(KEYINPUT98), .A2(G179), .A3(G200), .ZN(new_n785));
  OAI21_X1  g0585(.A(KEYINPUT98), .B1(G179), .B2(G200), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n632), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n206), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n773), .A2(new_n358), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G97), .A2(new_n789), .B1(new_n790), .B2(G50), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n206), .B(G190), .C1(new_n785), .C2(new_n786), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G159), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT32), .Z(new_n794));
  NAND4_X1  g0594(.A1(new_n778), .A2(new_n784), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  INV_X1    g0596(.A(new_n774), .ZN(new_n797));
  INV_X1    g0597(.A(new_n790), .ZN(new_n798));
  INV_X1    g0598(.A(G326), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n796), .A2(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G311), .B2(new_n776), .ZN(new_n801));
  INV_X1    g0601(.A(G303), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n333), .B1(new_n454), .B2(new_n781), .C1(new_n802), .C2(new_n780), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G329), .B2(new_n792), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT33), .B(G317), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n783), .A2(new_n805), .B1(new_n789), .B2(G294), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n801), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n770), .B1(new_n795), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n769), .A2(new_n766), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n695), .A2(new_n333), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n810), .A2(G355), .B1(new_n574), .B2(new_n695), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n241), .A2(G45), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT94), .Z(new_n813));
  NOR2_X1   g0613(.A1(new_n695), .A2(new_n389), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(G45), .B2(new_n219), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n811), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n757), .B(new_n808), .C1(new_n809), .C2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n761), .B1(new_n768), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  OAI21_X1  g0619(.A(new_n359), .B1(new_n357), .B2(new_n674), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n355), .ZN(new_n821));
  INV_X1    g0621(.A(new_n355), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n674), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n746), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n824), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n665), .A2(new_n674), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n756), .B1(new_n727), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n727), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n769), .A2(new_n762), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT99), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n757), .B1(new_n833), .B2(new_n202), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G283), .A2(new_n783), .B1(new_n774), .B2(G294), .ZN(new_n835));
  INV_X1    g0635(.A(new_n776), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n574), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n792), .ZN(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n333), .B1(new_n523), .B2(new_n781), .C1(new_n480), .C2(new_n780), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n798), .A2(new_n802), .B1(new_n478), .B2(new_n788), .ZN(new_n842));
  NOR4_X1   g0642(.A1(new_n837), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G137), .A2(new_n790), .B1(new_n774), .B2(G143), .ZN(new_n844));
  INV_X1    g0644(.A(G150), .ZN(new_n845));
  INV_X1    g0645(.A(new_n783), .ZN(new_n846));
  INV_X1    g0646(.A(G159), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n844), .B1(new_n845), .B2(new_n846), .C1(new_n847), .C2(new_n836), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT34), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n781), .A2(new_n247), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n380), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n419), .B2(new_n780), .C1(new_n838), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G58), .B2(new_n789), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n843), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n834), .B1(new_n770), .B2(new_n855), .C1(new_n826), .C2(new_n763), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n830), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NAND2_X1  g0658(.A1(new_n382), .A2(new_n254), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT16), .B1(new_n368), .B2(new_n370), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n388), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n404), .A2(new_n398), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(new_n409), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n861), .A2(new_n672), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n864), .A2(KEYINPUT103), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n863), .A2(new_n866), .A3(new_n409), .A4(new_n865), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT103), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n380), .A2(new_n363), .A3(new_n206), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n374), .A2(KEYINPUT7), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(G68), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT16), .B1(new_n874), .B2(new_n370), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n388), .B1(new_n859), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT102), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n878), .B(new_n388), .C1(new_n859), .C2(new_n875), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n672), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(new_n862), .A3(new_n879), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(new_n409), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n871), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n880), .B1(new_n406), .B2(new_n410), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n867), .A2(new_n870), .B1(new_n882), .B2(KEYINPUT37), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n885), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n887), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n864), .A2(new_n866), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n867), .A2(new_n870), .B1(new_n892), .B2(KEYINPUT37), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n866), .B1(new_n406), .B2(new_n410), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n888), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT39), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n268), .B(new_n674), .C1(new_n327), .C2(new_n331), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n646), .A2(KEYINPUT104), .A3(new_n674), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n406), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n897), .A2(new_n902), .B1(new_n903), .B2(new_n671), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n267), .A2(new_n674), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n332), .A2(new_n450), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n646), .B2(new_n449), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n907), .A2(new_n908), .B1(new_n827), .B2(new_n823), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n887), .A2(new_n890), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n410), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n447), .B(new_n445), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n822), .B1(new_n914), .B2(new_n442), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n913), .B1(new_n332), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n649), .B1(new_n916), .B2(new_n903), .ZN(new_n917));
  INV_X1    g0717(.A(new_n424), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n646), .A2(new_n439), .A3(new_n449), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n742), .A2(new_n920), .A3(new_n748), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n742), .A2(new_n920), .A3(KEYINPUT105), .A4(new_n748), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n912), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n887), .A2(new_n895), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n716), .A2(new_n717), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n824), .B1(new_n705), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n906), .B1(new_n332), .B2(new_n450), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n646), .A2(new_n449), .A3(new_n905), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n927), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT40), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT40), .B1(new_n887), .B2(new_n890), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n705), .A2(new_n928), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n920), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(G330), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n936), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n926), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n926), .A2(new_n941), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n942), .B(new_n943), .C1(new_n205), .C2(new_n753), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n494), .A2(new_n495), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT35), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(G116), .A3(new_n217), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT100), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n948), .A2(new_n949), .B1(new_n946), .B2(new_n945), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT36), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT36), .ZN(new_n953));
  INV_X1    g0753(.A(G58), .ZN(new_n954));
  OAI21_X1  g0754(.A(G77), .B1(new_n954), .B2(new_n247), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n955), .A2(new_n219), .B1(G50), .B2(new_n247), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n213), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT101), .Z(new_n958));
  NAND4_X1  g0758(.A1(new_n944), .A2(new_n952), .A3(new_n953), .A4(new_n958), .ZN(G367));
  OAI21_X1  g0759(.A(new_n809), .B1(new_n209), .B2(new_n346), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n236), .A2(new_n695), .A3(new_n389), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n756), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n419), .A2(new_n836), .B1(new_n846), .B2(new_n847), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n790), .A2(G143), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n789), .A2(G68), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(new_n797), .C2(new_n845), .ZN(new_n966));
  INV_X1    g0766(.A(new_n781), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n333), .B1(G77), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(G137), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n968), .B1(new_n954), .B2(new_n780), .C1(new_n969), .C2(new_n838), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n963), .A2(new_n966), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT110), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n454), .A2(new_n836), .B1(new_n798), .B2(new_n839), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n797), .A2(new_n802), .B1(new_n480), .B2(new_n788), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n389), .B1(G97), .B2(new_n967), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n780), .A2(new_n574), .ZN(new_n976));
  INV_X1    g0776(.A(G317), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n975), .B1(KEYINPUT46), .B2(new_n976), .C1(new_n838), .C2(new_n977), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n973), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n976), .A2(KEYINPUT46), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n783), .A2(G294), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n979), .B(new_n982), .C1(new_n980), .C2(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n972), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT47), .Z(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n770), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n680), .A2(new_n552), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n658), .B(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n962), .B(new_n986), .C1(new_n766), .C2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n692), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n738), .B1(new_n502), .B2(new_n674), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n730), .A2(new_n652), .A3(new_n680), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n990), .A2(KEYINPUT42), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n630), .ZN(new_n996));
  INV_X1    g0796(.A(new_n518), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n674), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT42), .B1(new_n990), .B2(new_n994), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT106), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n988), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n988), .A2(new_n1002), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1004), .A2(new_n689), .A3(new_n993), .A4(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT107), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n690), .B2(new_n994), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(KEYINPUT107), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n693), .A2(new_n993), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT44), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n990), .A2(new_n679), .A3(new_n993), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n689), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1014), .A2(new_n690), .A3(new_n1016), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT108), .B1(new_n688), .B2(new_n691), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n678), .B(new_n1021), .Z(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(new_n990), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n751), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n696), .B(KEYINPUT41), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n755), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n989), .B1(new_n1012), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT111), .ZN(G387));
  NOR2_X1   g0830(.A1(new_n1023), .A2(new_n750), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1023), .A2(new_n750), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n696), .B(KEYINPUT114), .Z(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n389), .B1(G116), .B2(new_n967), .ZN(new_n1036));
  INV_X1    g0836(.A(G294), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n788), .A2(new_n454), .B1(new_n1037), .B2(new_n780), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G317), .A2(new_n774), .B1(new_n790), .B2(G322), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n802), .B2(new_n836), .C1(new_n839), .C2(new_n846), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1036), .B1(new_n799), .B2(new_n838), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n774), .A2(G50), .B1(new_n789), .B2(new_n347), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT113), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n380), .B1(G97), .B2(new_n967), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n202), .B2(new_n780), .C1(new_n838), .C2(new_n845), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G68), .A2(new_n776), .B1(new_n790), .B2(G159), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n386), .B2(new_n846), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1048), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n769), .B1(new_n1046), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n698), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n810), .A2(new_n1055), .B1(new_n480), .B2(new_n695), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n233), .A2(new_n276), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n344), .A2(new_n419), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  AOI21_X1  g0861(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1060), .A2(new_n698), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n814), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1056), .B1(new_n1057), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n757), .B1(new_n1065), .B2(new_n809), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1054), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n688), .B2(new_n766), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1023), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n755), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1035), .A2(new_n1070), .ZN(G393));
  OAI21_X1  g0871(.A(new_n809), .B1(new_n478), .B2(new_n209), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n814), .A2(new_n244), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n756), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G311), .A2(new_n774), .B1(new_n790), .B2(G317), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n776), .A2(G294), .B1(new_n789), .B2(G116), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n802), .B2(new_n846), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n838), .A2(new_n796), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n333), .B1(new_n480), .B2(new_n781), .C1(new_n454), .C2(new_n780), .ZN(new_n1081));
  NOR4_X1   g0881(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT116), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G150), .A2(new_n790), .B1(new_n774), .B2(G159), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT51), .Z(new_n1086));
  OAI221_X1 g0886(.A(new_n389), .B1(new_n247), .B2(new_n780), .C1(new_n523), .C2(new_n781), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G143), .B2(new_n792), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n783), .A2(G50), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G77), .A2(new_n789), .B1(new_n776), .B2(new_n344), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1083), .A2(KEYINPUT116), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1084), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1074), .B1(new_n1093), .B2(new_n769), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n993), .B2(new_n767), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1020), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(new_n1031), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1034), .B1(new_n1020), .B2(new_n1032), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1095), .B1(new_n754), .B2(new_n1020), .C1(new_n1097), .C2(new_n1098), .ZN(G390));
  NAND3_X1  g0899(.A1(new_n741), .A2(new_n674), .A3(new_n821), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n823), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n907), .A2(new_n908), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n900), .A2(new_n927), .A3(new_n901), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT39), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n927), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n887), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n909), .B2(new_n902), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n725), .A2(G330), .A3(new_n826), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1102), .A2(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1106), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n759), .B(new_n824), .C1(new_n705), .C2(new_n928), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n930), .B2(new_n931), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n755), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G107), .A2(new_n783), .B1(new_n790), .B2(G283), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n574), .B2(new_n797), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n776), .A2(G97), .B1(new_n789), .B2(G77), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n780), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n294), .B(new_n850), .C1(G87), .C2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(new_n1037), .C2(new_n838), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT54), .B(G143), .Z(new_n1126));
  INV_X1    g0926(.A(KEYINPUT53), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n780), .B2(new_n845), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1123), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n776), .A2(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n294), .B1(new_n419), .B2(new_n781), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G125), .B2(new_n792), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(new_n969), .C2(new_n846), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n790), .A2(G128), .B1(new_n789), .B2(G159), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n852), .B2(new_n797), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1121), .A2(new_n1125), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n769), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n757), .B1(new_n833), .B2(new_n386), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(new_n897), .C2(new_n763), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1119), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n937), .A2(G330), .A3(new_n826), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n907), .A3(new_n908), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1101), .B1(new_n1102), .B2(new_n1112), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n725), .A2(G330), .A3(new_n826), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(new_n907), .A3(new_n908), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1116), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n827), .A2(new_n823), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1143), .A2(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n939), .A2(G330), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT29), .B1(new_n665), .B2(new_n674), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n451), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT105), .B1(new_n1152), .B2(new_n742), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n924), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n650), .B(new_n1150), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT117), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1145), .A2(new_n907), .A3(new_n908), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1142), .B1(new_n907), .B2(new_n908), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1148), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1113), .A2(new_n823), .A3(new_n1100), .A4(new_n1143), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT117), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1161), .A2(new_n925), .A3(new_n1162), .A4(new_n1150), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1148), .B1(new_n930), .B2(new_n931), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n900), .A2(new_n901), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1164), .A2(new_n1165), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1104), .B1(new_n1102), .B2(new_n1101), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1158), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1106), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1156), .A2(new_n1163), .A3(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(KEYINPUT118), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT118), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1156), .A2(new_n1163), .A3(new_n1173), .A4(new_n1170), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1034), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1149), .A2(new_n1155), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1118), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1141), .B1(new_n1172), .B2(new_n1178), .ZN(G378));
  AOI21_X1  g0979(.A(KEYINPUT122), .B1(new_n904), .B2(new_n911), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n422), .A2(new_n672), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT55), .Z(new_n1183));
  XNOR2_X1  g0983(.A(new_n438), .B(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1185));
  XOR2_X1   g0985(.A(new_n1184), .B(new_n1185), .Z(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n936), .B2(G330), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n639), .A2(new_n556), .A3(new_n680), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n721), .A2(new_n723), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n826), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n907), .B2(new_n908), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n932), .A2(KEYINPUT40), .B1(new_n1192), .B2(new_n934), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1193), .A2(new_n759), .A3(new_n1186), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1181), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1186), .B1(new_n1193), .B2(new_n759), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT40), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1192), .B2(new_n927), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n935), .ZN(new_n1199));
  OAI211_X1 g0999(.A(G330), .B(new_n1187), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(new_n1180), .A3(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1195), .A2(new_n755), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n757), .B1(new_n833), .B2(new_n419), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n965), .B1(new_n798), .B2(new_n574), .C1(new_n480), .C2(new_n797), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n838), .A2(new_n454), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n389), .A2(G41), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n781), .A2(new_n954), .B1(new_n780), .B2(new_n202), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G97), .A2(new_n783), .B1(new_n776), .B2(new_n347), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT119), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT120), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(G33), .A2(G41), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1206), .A2(G50), .A3(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G132), .A2(new_n783), .B1(new_n776), .B2(G137), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G125), .A2(new_n790), .B1(new_n774), .B2(G128), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n789), .A2(G150), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n792), .A2(G124), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1223), .B(new_n1216), .C1(new_n847), .C2(new_n781), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1221), .B2(KEYINPUT59), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1217), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1214), .A2(new_n1215), .A3(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1203), .B1(new_n770), .B2(new_n1227), .C1(new_n1187), .C2(new_n763), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1202), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1155), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1170), .B2(new_n1149), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT57), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n897), .A2(new_n902), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n903), .A2(new_n671), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1233), .A2(new_n911), .A3(new_n1234), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1196), .A2(new_n1235), .A3(new_n1200), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1034), .B1(new_n1232), .B2(new_n1238), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1196), .A2(new_n1180), .A3(new_n1200), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1180), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT57), .B1(new_n1242), .B2(new_n1231), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1229), .B1(new_n1239), .B2(new_n1243), .ZN(G375));
  NAND2_X1  g1044(.A1(new_n1149), .A2(new_n1155), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1156), .A2(new_n1163), .A3(new_n1026), .A4(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n907), .A2(new_n908), .A3(new_n762), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n574), .A2(new_n846), .B1(new_n798), .B2(new_n1037), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G283), .B2(new_n774), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n333), .B1(new_n202), .B2(new_n781), .C1(new_n478), .C2(new_n780), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G303), .B2(new_n792), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n776), .A2(G107), .B1(new_n789), .B2(new_n347), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G132), .A2(new_n790), .B1(new_n783), .B2(new_n1126), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n774), .A2(G137), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n389), .B1(new_n954), .B2(new_n781), .C1(new_n847), .C2(new_n780), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G128), .B2(new_n792), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n776), .A2(G150), .B1(new_n789), .B2(G50), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n770), .B1(new_n1253), .B2(new_n1259), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n757), .B(new_n1260), .C1(new_n247), .C2(new_n833), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1161), .A2(new_n755), .B1(new_n1247), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1246), .A2(new_n1262), .ZN(G381));
  NAND3_X1  g1063(.A1(new_n1035), .A2(new_n818), .A3(new_n1070), .ZN(new_n1264));
  OR4_X1    g1064(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1264), .ZN(new_n1265));
  OR4_X1    g1065(.A1(G387), .A2(new_n1265), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1066(.A1(new_n1202), .A2(new_n1228), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT57), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1230), .A2(new_n1169), .A3(new_n1168), .A4(new_n1161), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n1230), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n912), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1196), .A2(new_n1235), .A3(new_n1200), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1175), .B1(new_n1270), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1195), .A2(new_n1201), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1155), .B1(new_n1118), .B2(new_n1176), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1268), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1267), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1178), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1171), .A2(KEYINPUT118), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1140), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(G343), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(G213), .ZN(new_n1283));
  XOR2_X1   g1083(.A(new_n1283), .B(KEYINPUT123), .Z(new_n1284));
  NAND3_X1  g1084(.A1(new_n1278), .A2(new_n1281), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G407), .A2(G213), .A3(new_n1285), .ZN(G409));
  NAND2_X1  g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1264), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G390), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT111), .B1(new_n1287), .B2(new_n1264), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1289), .B1(G390), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1029), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n989), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(new_n1027), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1295), .B(new_n1289), .C1(G390), .C2(new_n1290), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT124), .B1(G375), .B2(new_n1281), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT124), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1278), .A2(new_n1300), .A3(G378), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n755), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT125), .B1(new_n1303), .B2(new_n1228), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1275), .A2(new_n1276), .A3(new_n1025), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1303), .A2(KEYINPUT125), .A3(new_n1228), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1305), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1281), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1284), .B1(new_n1302), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1245), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT60), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1245), .A2(new_n1312), .A3(KEYINPUT60), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1176), .A2(new_n1175), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G384), .B1(new_n1319), .B2(new_n1262), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1262), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n857), .B(new_n1321), .C1(new_n1317), .C2(new_n1318), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT63), .B1(new_n1311), .B2(new_n1323), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1325));
  AOI21_X1  g1125(.A(G378), .B1(new_n1325), .B2(new_n1308), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1323), .ZN(new_n1329));
  NOR4_X1   g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1329), .A4(new_n1284), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1298), .B1(new_n1324), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1284), .A2(G2897), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1320), .A2(new_n1322), .A3(new_n1333), .ZN(new_n1334));
  AOI211_X1 g1134(.A(new_n1175), .B(new_n1176), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n857), .B1(new_n1335), .B2(new_n1321), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1319), .A2(G384), .A3(new_n1262), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1332), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1334), .A2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1339), .B1(new_n1327), .B2(new_n1284), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT61), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT127), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1331), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1346));
  AND4_X1   g1146(.A1(new_n1300), .A2(new_n1346), .A3(G378), .A4(new_n1229), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1300), .B1(new_n1278), .B2(G378), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1310), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1284), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1349), .A2(new_n1350), .A3(new_n1323), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(KEYINPUT62), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT62), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1349), .A2(new_n1353), .A3(new_n1350), .A4(new_n1323), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1352), .A2(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(KEYINPUT127), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1297), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1345), .A2(new_n1357), .ZN(G405));
  AOI22_X1  g1158(.A1(new_n1299), .A2(new_n1301), .B1(new_n1281), .B2(G375), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1359), .B(new_n1329), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1360), .B(new_n1297), .ZN(G402));
endmodule


