

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(n522), .B(KEYINPUT69), .ZN(n646) );
  NAND2_X1 U551 ( .A1(n677), .A2(n767), .ZN(n723) );
  OR2_X1 U552 ( .A1(n693), .A2(n692), .ZN(n705) );
  NOR2_X1 U553 ( .A1(n921), .A2(n706), .ZN(n708) );
  INV_X1 U554 ( .A(KEYINPUT27), .ZN(n697) );
  INV_X1 U555 ( .A(KEYINPUT28), .ZN(n707) );
  INV_X1 U556 ( .A(n934), .ZN(n746) );
  AND2_X1 U557 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U558 ( .A1(n749), .A2(n748), .ZN(n752) );
  NOR2_X1 U559 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U560 ( .A(n592), .B(KEYINPUT78), .ZN(n695) );
  INV_X1 U561 ( .A(n695), .ZN(n891) );
  NOR2_X1 U562 ( .A1(n626), .A2(G651), .ZN(n640) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n519) );
  XNOR2_X1 U564 ( .A(n519), .B(KEYINPUT64), .ZN(n645) );
  NAND2_X1 U565 ( .A1(G89), .A2(n645), .ZN(n520) );
  XNOR2_X1 U566 ( .A(n520), .B(KEYINPUT4), .ZN(n524) );
  XOR2_X1 U567 ( .A(G651), .B(KEYINPUT68), .Z(n526) );
  XNOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .ZN(n521) );
  XNOR2_X1 U569 ( .A(n521), .B(KEYINPUT67), .ZN(n626) );
  OR2_X1 U570 ( .A1(n526), .A2(n626), .ZN(n522) );
  NAND2_X1 U571 ( .A1(G76), .A2(n646), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U573 ( .A(n525), .B(KEYINPUT5), .ZN(n532) );
  NOR2_X1 U574 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n527), .Z(n641) );
  NAND2_X1 U576 ( .A1(G63), .A2(n641), .ZN(n529) );
  NAND2_X1 U577 ( .A1(G51), .A2(n640), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U579 ( .A(KEYINPUT6), .B(n530), .Z(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U581 ( .A(n533), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U582 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U583 ( .A1(n640), .A2(G53), .ZN(n540) );
  NAND2_X1 U584 ( .A1(G65), .A2(n641), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G78), .A2(n646), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n538) );
  NAND2_X1 U587 ( .A1(n645), .A2(G91), .ZN(n536) );
  XOR2_X1 U588 ( .A(KEYINPUT72), .B(n536), .Z(n537) );
  NOR2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U591 ( .A(KEYINPUT73), .B(n541), .Z(G299) );
  INV_X1 U592 ( .A(G2105), .ZN(n543) );
  AND2_X1 U593 ( .A1(n543), .A2(G2104), .ZN(n864) );
  NAND2_X1 U594 ( .A1(G101), .A2(n864), .ZN(n542) );
  XOR2_X1 U595 ( .A(KEYINPUT23), .B(n542), .Z(n548) );
  NOR2_X1 U596 ( .A1(G2104), .A2(n543), .ZN(n868) );
  NAND2_X1 U597 ( .A1(G125), .A2(n868), .ZN(n546) );
  NAND2_X1 U598 ( .A1(G2105), .A2(G2104), .ZN(n544) );
  XNOR2_X2 U599 ( .A(n544), .B(KEYINPUT65), .ZN(n869) );
  NAND2_X1 U600 ( .A1(G113), .A2(n869), .ZN(n545) );
  AND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n676) );
  NOR2_X1 U603 ( .A1(G2104), .A2(G2105), .ZN(n549) );
  XOR2_X2 U604 ( .A(KEYINPUT17), .B(n549), .Z(n865) );
  NAND2_X1 U605 ( .A1(G137), .A2(n865), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n550), .B(KEYINPUT66), .ZN(n765) );
  AND2_X1 U607 ( .A1(n676), .A2(n765), .ZN(G160) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U609 ( .A(G57), .ZN(G237) );
  NAND2_X1 U610 ( .A1(G64), .A2(n641), .ZN(n552) );
  NAND2_X1 U611 ( .A1(G52), .A2(n640), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n646), .A2(G77), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G90), .A2(n645), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U618 ( .A(KEYINPUT71), .B(n558), .Z(G171) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  NAND2_X1 U620 ( .A1(n646), .A2(G75), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G88), .A2(n645), .ZN(n559) );
  NAND2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U623 ( .A1(G62), .A2(n641), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G50), .A2(n640), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U626 ( .A1(n564), .A2(n563), .ZN(G166) );
  NAND2_X1 U627 ( .A1(G102), .A2(n864), .ZN(n566) );
  NAND2_X1 U628 ( .A1(G138), .A2(n865), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G126), .A2(n868), .ZN(n568) );
  NAND2_X1 U631 ( .A1(G114), .A2(n869), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n570), .A2(n569), .ZN(G164) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n571), .B(KEYINPUT10), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT74), .B(n572), .ZN(G223) );
  XNOR2_X1 U637 ( .A(KEYINPUT75), .B(G223), .ZN(n818) );
  NAND2_X1 U638 ( .A1(n818), .A2(G567), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  NAND2_X1 U640 ( .A1(G81), .A2(n645), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G68), .A2(n646), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(KEYINPUT76), .Z(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n641), .A2(G56), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT14), .B(n579), .Z(n580) );
  NOR2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n640), .A2(G43), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n926) );
  INV_X1 U651 ( .A(G860), .ZN(n617) );
  OR2_X1 U652 ( .A1(n926), .A2(n617), .ZN(G153) );
  NAND2_X1 U653 ( .A1(n645), .A2(G92), .ZN(n590) );
  NAND2_X1 U654 ( .A1(G66), .A2(n641), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G54), .A2(n640), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G79), .A2(n646), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n586), .B(KEYINPUT77), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT15), .ZN(n592) );
  INV_X1 U661 ( .A(n891), .ZN(n925) );
  NOR2_X1 U662 ( .A1(G868), .A2(n925), .ZN(n593) );
  XNOR2_X1 U663 ( .A(n593), .B(KEYINPUT79), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(G284) );
  NOR2_X1 U666 ( .A1(G868), .A2(G299), .ZN(n596) );
  XNOR2_X1 U667 ( .A(n596), .B(KEYINPUT80), .ZN(n598) );
  INV_X1 U668 ( .A(G868), .ZN(n659) );
  NOR2_X1 U669 ( .A1(n659), .A2(G286), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U671 ( .A(KEYINPUT81), .B(n599), .Z(G297) );
  NAND2_X1 U672 ( .A1(n617), .A2(G559), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n600), .A2(n925), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U675 ( .A1(G868), .A2(n926), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n925), .A2(G868), .ZN(n602) );
  NOR2_X1 U677 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U678 ( .A1(n604), .A2(n603), .ZN(G282) );
  XOR2_X1 U679 ( .A(KEYINPUT82), .B(KEYINPUT18), .Z(n606) );
  NAND2_X1 U680 ( .A1(G123), .A2(n868), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n606), .B(n605), .ZN(n613) );
  NAND2_X1 U682 ( .A1(G99), .A2(n864), .ZN(n608) );
  NAND2_X1 U683 ( .A1(G111), .A2(n869), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT83), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G135), .A2(n865), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n996) );
  XNOR2_X1 U689 ( .A(G2096), .B(n996), .ZN(n615) );
  INV_X1 U690 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U692 ( .A1(n925), .A2(G559), .ZN(n616) );
  XOR2_X1 U693 ( .A(n926), .B(n616), .Z(n656) );
  NAND2_X1 U694 ( .A1(n617), .A2(n656), .ZN(n625) );
  NAND2_X1 U695 ( .A1(G55), .A2(n640), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G93), .A2(n645), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n646), .A2(G80), .ZN(n620) );
  XOR2_X1 U699 ( .A(KEYINPUT84), .B(n620), .Z(n621) );
  NOR2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n641), .A2(G67), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n658) );
  XNOR2_X1 U703 ( .A(n625), .B(n658), .ZN(G145) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G87), .A2(n626), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n641), .A2(n629), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G49), .A2(n640), .ZN(n630) );
  XOR2_X1 U709 ( .A(KEYINPUT85), .B(n630), .Z(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G48), .A2(n640), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G86), .A2(n645), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n646), .A2(G73), .ZN(n635) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n635), .Z(n636) );
  NOR2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n641), .A2(G61), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n639), .A2(n638), .ZN(G305) );
  NAND2_X1 U719 ( .A1(n640), .A2(G47), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n641), .A2(G60), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U722 ( .A(KEYINPUT70), .B(n644), .Z(n650) );
  NAND2_X1 U723 ( .A1(n645), .A2(G85), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n646), .A2(G72), .ZN(n647) );
  AND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(G290) );
  XNOR2_X1 U727 ( .A(KEYINPUT19), .B(G288), .ZN(n655) );
  INV_X1 U728 ( .A(G299), .ZN(n921) );
  XNOR2_X1 U729 ( .A(n921), .B(G305), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(n658), .ZN(n652) );
  XNOR2_X1 U731 ( .A(G166), .B(n652), .ZN(n653) );
  XNOR2_X1 U732 ( .A(n653), .B(G290), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(n894) );
  XNOR2_X1 U734 ( .A(n656), .B(n894), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U740 ( .A1(n663), .A2(G2090), .ZN(n664) );
  XNOR2_X1 U741 ( .A(n664), .B(KEYINPUT86), .ZN(n665) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U743 ( .A1(G2072), .A2(n666), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U745 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n668) );
  NAND2_X1 U746 ( .A1(G132), .A2(G82), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U748 ( .A1(n669), .A2(G218), .ZN(n670) );
  NAND2_X1 U749 ( .A1(G96), .A2(n670), .ZN(n822) );
  NAND2_X1 U750 ( .A1(n822), .A2(G2106), .ZN(n674) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n671) );
  NOR2_X1 U752 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G108), .A2(n672), .ZN(n823) );
  NAND2_X1 U754 ( .A1(n823), .A2(G567), .ZN(n673) );
  NAND2_X1 U755 ( .A1(n674), .A2(n673), .ZN(n824) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U757 ( .A1(n824), .A2(n675), .ZN(n821) );
  NAND2_X1 U758 ( .A1(n821), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G166), .ZN(G303) );
  AND2_X1 U760 ( .A1(n676), .A2(G40), .ZN(n764) );
  AND2_X1 U761 ( .A1(n765), .A2(n764), .ZN(n677) );
  NOR2_X1 U762 ( .A1(G164), .A2(G1384), .ZN(n767) );
  NAND2_X1 U763 ( .A1(G8), .A2(n723), .ZN(n758) );
  NOR2_X1 U764 ( .A1(G1981), .A2(G305), .ZN(n678) );
  XOR2_X1 U765 ( .A(n678), .B(KEYINPUT92), .Z(n679) );
  XNOR2_X1 U766 ( .A(KEYINPUT24), .B(n679), .ZN(n680) );
  NOR2_X1 U767 ( .A1(n758), .A2(n680), .ZN(n763) );
  XNOR2_X1 U768 ( .A(G1961), .B(KEYINPUT93), .ZN(n964) );
  NAND2_X1 U769 ( .A1(n964), .A2(n723), .ZN(n682) );
  INV_X1 U770 ( .A(n723), .ZN(n687) );
  XNOR2_X1 U771 ( .A(KEYINPUT25), .B(G2078), .ZN(n953) );
  NAND2_X1 U772 ( .A1(n687), .A2(n953), .ZN(n681) );
  NAND2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U774 ( .A(n683), .B(KEYINPUT94), .ZN(n717) );
  NAND2_X1 U775 ( .A1(G171), .A2(n717), .ZN(n713) );
  NAND2_X1 U776 ( .A1(G1348), .A2(n723), .ZN(n685) );
  NAND2_X1 U777 ( .A1(G2067), .A2(n687), .ZN(n684) );
  NAND2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U779 ( .A(KEYINPUT97), .B(n686), .ZN(n694) );
  NOR2_X1 U780 ( .A1(n695), .A2(n694), .ZN(n693) );
  XNOR2_X1 U781 ( .A(G1996), .B(KEYINPUT96), .ZN(n948) );
  NAND2_X1 U782 ( .A1(n948), .A2(n687), .ZN(n688) );
  XNOR2_X1 U783 ( .A(n688), .B(KEYINPUT26), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n723), .A2(G1341), .ZN(n689) );
  NAND2_X1 U785 ( .A1(n690), .A2(n689), .ZN(n691) );
  OR2_X1 U786 ( .A1(n926), .A2(n691), .ZN(n692) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n703) );
  INV_X1 U788 ( .A(G2072), .ZN(n696) );
  OR2_X1 U789 ( .A1(n723), .A2(n696), .ZN(n698) );
  XNOR2_X1 U790 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n723), .A2(G1956), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U793 ( .A(n701), .B(KEYINPUT95), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n921), .A2(n706), .ZN(n702) );
  AND2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n710) );
  XNOR2_X1 U797 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U798 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U799 ( .A(KEYINPUT29), .B(n711), .Z(n712) );
  NAND2_X1 U800 ( .A1(n713), .A2(n712), .ZN(n722) );
  NOR2_X1 U801 ( .A1(G1966), .A2(n758), .ZN(n735) );
  NOR2_X1 U802 ( .A1(G2084), .A2(n723), .ZN(n731) );
  NOR2_X1 U803 ( .A1(n735), .A2(n731), .ZN(n714) );
  NAND2_X1 U804 ( .A1(G8), .A2(n714), .ZN(n715) );
  XNOR2_X1 U805 ( .A(KEYINPUT30), .B(n715), .ZN(n716) );
  NOR2_X1 U806 ( .A1(G168), .A2(n716), .ZN(n719) );
  NOR2_X1 U807 ( .A1(G171), .A2(n717), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U809 ( .A(KEYINPUT31), .B(n720), .Z(n721) );
  NAND2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n733) );
  NAND2_X1 U811 ( .A1(n733), .A2(G286), .ZN(n728) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n758), .ZN(n725) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n723), .ZN(n724) );
  NOR2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U815 ( .A1(n726), .A2(G303), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U817 ( .A1(n729), .A2(G8), .ZN(n730) );
  XNOR2_X1 U818 ( .A(n730), .B(KEYINPUT32), .ZN(n737) );
  NAND2_X1 U819 ( .A1(G8), .A2(n731), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n734) );
  OR2_X1 U821 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U822 ( .A1(n737), .A2(n736), .ZN(n756) );
  NOR2_X1 U823 ( .A1(G1971), .A2(G303), .ZN(n738) );
  XNOR2_X1 U824 ( .A(n738), .B(KEYINPUT99), .ZN(n740) );
  NOR2_X1 U825 ( .A1(G288), .A2(G1976), .ZN(n739) );
  XOR2_X1 U826 ( .A(n739), .B(KEYINPUT98), .Z(n920) );
  AND2_X1 U827 ( .A1(n740), .A2(n920), .ZN(n742) );
  INV_X1 U828 ( .A(KEYINPUT33), .ZN(n741) );
  AND2_X1 U829 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U830 ( .A1(n756), .A2(n743), .ZN(n749) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n915) );
  INV_X1 U832 ( .A(n915), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n744), .A2(n758), .ZN(n745) );
  OR2_X1 U834 ( .A1(KEYINPUT33), .A2(n745), .ZN(n747) );
  XNOR2_X1 U835 ( .A(G1981), .B(G305), .ZN(n934) );
  NOR2_X1 U836 ( .A1(n758), .A2(n920), .ZN(n750) );
  NAND2_X1 U837 ( .A1(KEYINPUT33), .A2(n750), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U839 ( .A(n753), .B(KEYINPUT100), .ZN(n761) );
  NAND2_X1 U840 ( .A1(G8), .A2(G166), .ZN(n754) );
  NOR2_X1 U841 ( .A1(G2090), .A2(n754), .ZN(n755) );
  XNOR2_X1 U842 ( .A(n755), .B(KEYINPUT101), .ZN(n757) );
  NAND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U845 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U846 ( .A1(n763), .A2(n762), .ZN(n797) );
  NAND2_X1 U847 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U848 ( .A1(n767), .A2(n766), .ZN(n813) );
  XOR2_X1 U849 ( .A(n813), .B(KEYINPUT91), .Z(n785) );
  NAND2_X1 U850 ( .A1(G141), .A2(n865), .ZN(n768) );
  XNOR2_X1 U851 ( .A(n768), .B(KEYINPUT90), .ZN(n775) );
  NAND2_X1 U852 ( .A1(G129), .A2(n868), .ZN(n770) );
  NAND2_X1 U853 ( .A1(G117), .A2(n869), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U855 ( .A1(n864), .A2(G105), .ZN(n771) );
  XOR2_X1 U856 ( .A(KEYINPUT38), .B(n771), .Z(n772) );
  NOR2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U858 ( .A1(n775), .A2(n774), .ZN(n881) );
  NAND2_X1 U859 ( .A1(G1996), .A2(n881), .ZN(n784) );
  NAND2_X1 U860 ( .A1(G95), .A2(n864), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G131), .A2(n865), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U863 ( .A(KEYINPUT89), .B(n778), .ZN(n782) );
  NAND2_X1 U864 ( .A1(G119), .A2(n868), .ZN(n780) );
  NAND2_X1 U865 ( .A1(G107), .A2(n869), .ZN(n779) );
  AND2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n875) );
  NAND2_X1 U868 ( .A1(G1991), .A2(n875), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n994) );
  NAND2_X1 U870 ( .A1(n785), .A2(n994), .ZN(n803) );
  NAND2_X1 U871 ( .A1(G104), .A2(n864), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G140), .A2(n865), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U874 ( .A(KEYINPUT34), .B(n788), .ZN(n793) );
  NAND2_X1 U875 ( .A1(G128), .A2(n868), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G116), .A2(n869), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U878 ( .A(n791), .B(KEYINPUT35), .Z(n792) );
  NOR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U880 ( .A(KEYINPUT36), .B(n794), .Z(n795) );
  XOR2_X1 U881 ( .A(KEYINPUT88), .B(n795), .Z(n889) );
  XNOR2_X1 U882 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  NOR2_X1 U883 ( .A1(n889), .A2(n811), .ZN(n997) );
  NAND2_X1 U884 ( .A1(n813), .A2(n997), .ZN(n809) );
  NAND2_X1 U885 ( .A1(n803), .A2(n809), .ZN(n796) );
  NOR2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n798), .B(KEYINPUT102), .ZN(n800) );
  XNOR2_X1 U888 ( .A(G1986), .B(G290), .ZN(n918) );
  NAND2_X1 U889 ( .A1(n918), .A2(n813), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n816) );
  XOR2_X1 U891 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n808) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n881), .ZN(n1009) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U894 ( .A1(G1991), .A2(n875), .ZN(n1001) );
  NOR2_X1 U895 ( .A1(n801), .A2(n1001), .ZN(n802) );
  XNOR2_X1 U896 ( .A(n802), .B(KEYINPUT103), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U898 ( .A(KEYINPUT104), .B(n805), .Z(n806) );
  NOR2_X1 U899 ( .A1(n1009), .A2(n806), .ZN(n807) );
  XNOR2_X1 U900 ( .A(n808), .B(n807), .ZN(n810) );
  NAND2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U902 ( .A1(n889), .A2(n811), .ZN(n993) );
  NAND2_X1 U903 ( .A1(n812), .A2(n993), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U906 ( .A(n817), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n818), .ZN(G217) );
  AND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U909 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(G188) );
  INV_X1 U913 ( .A(G132), .ZN(G219) );
  INV_X1 U914 ( .A(G120), .ZN(G236) );
  INV_X1 U915 ( .A(G96), .ZN(G221) );
  INV_X1 U916 ( .A(G82), .ZN(G220) );
  INV_X1 U917 ( .A(G69), .ZN(G235) );
  NOR2_X1 U918 ( .A1(n823), .A2(n822), .ZN(G325) );
  INV_X1 U919 ( .A(G325), .ZN(G261) );
  INV_X1 U920 ( .A(n824), .ZN(G319) );
  XOR2_X1 U921 ( .A(G2474), .B(G1981), .Z(n826) );
  XNOR2_X1 U922 ( .A(G1996), .B(G1991), .ZN(n825) );
  XNOR2_X1 U923 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U924 ( .A(n827), .B(KEYINPUT110), .Z(n829) );
  XNOR2_X1 U925 ( .A(G1971), .B(G1976), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U927 ( .A(G1956), .B(G1961), .Z(n831) );
  XNOR2_X1 U928 ( .A(G1986), .B(G1966), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U930 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U931 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(G229) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2078), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n836), .B(KEYINPUT43), .ZN(n846) );
  XOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .Z(n838) );
  XNOR2_X1 U936 ( .A(KEYINPUT107), .B(G2096), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U938 ( .A(G2100), .B(G2090), .Z(n840) );
  XNOR2_X1 U939 ( .A(G2072), .B(G2084), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U942 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(G227) );
  NAND2_X1 U945 ( .A1(G124), .A2(n868), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n847), .B(KEYINPUT112), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U948 ( .A1(G100), .A2(n864), .ZN(n849) );
  NAND2_X1 U949 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U950 ( .A1(G136), .A2(n865), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G112), .A2(n869), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U953 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U954 ( .A(KEYINPUT113), .B(n855), .Z(G162) );
  NAND2_X1 U955 ( .A1(G130), .A2(n868), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G118), .A2(n869), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G106), .A2(n864), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G142), .A2(n865), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U961 ( .A(KEYINPUT45), .B(n860), .Z(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n996), .B(n863), .ZN(n877) );
  NAND2_X1 U964 ( .A1(G103), .A2(n864), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G139), .A2(n865), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n874) );
  NAND2_X1 U967 ( .A1(G127), .A2(n868), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G115), .A2(n869), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n1004) );
  XNOR2_X1 U972 ( .A(n875), .B(n1004), .ZN(n876) );
  XNOR2_X1 U973 ( .A(n877), .B(n876), .ZN(n885) );
  XOR2_X1 U974 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n879) );
  XNOR2_X1 U975 ( .A(G164), .B(KEYINPUT115), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U977 ( .A(KEYINPUT114), .B(n880), .ZN(n883) );
  XNOR2_X1 U978 ( .A(n881), .B(KEYINPUT46), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U980 ( .A(n885), .B(n884), .Z(n887) );
  XNOR2_X1 U981 ( .A(G160), .B(G162), .ZN(n886) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U983 ( .A(n889), .B(n888), .Z(n890) );
  NOR2_X1 U984 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U985 ( .A(n926), .B(KEYINPUT117), .ZN(n893) );
  XNOR2_X1 U986 ( .A(G171), .B(n891), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n893), .B(n892), .ZN(n896) );
  XNOR2_X1 U988 ( .A(G286), .B(n894), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U990 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2438), .B(KEYINPUT106), .Z(n899) );
  XNOR2_X1 U992 ( .A(G2443), .B(G2430), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U994 ( .A(n900), .B(G2435), .Z(n902) );
  XNOR2_X1 U995 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U997 ( .A(G2451), .B(G2427), .Z(n904) );
  XNOR2_X1 U998 ( .A(G2454), .B(G2446), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1000 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n907), .ZN(n913) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  INV_X1 U1010 ( .A(n913), .ZN(G401) );
  XOR2_X1 U1011 ( .A(G16), .B(KEYINPUT118), .Z(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT56), .B(n914), .ZN(n941) );
  XNOR2_X1 U1013 ( .A(G166), .B(G1971), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n923) );
  XOR2_X1 U1017 ( .A(G1956), .B(n921), .Z(n922) );
  NOR2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1019 ( .A(KEYINPUT120), .B(n924), .Z(n939) );
  XNOR2_X1 U1020 ( .A(n925), .B(G1348), .ZN(n929) );
  XNOR2_X1 U1021 ( .A(G1341), .B(KEYINPUT121), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(n927), .B(n926), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n932) );
  XOR2_X1 U1024 ( .A(G1961), .B(G301), .Z(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT119), .B(n930), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n937) );
  XOR2_X1 U1027 ( .A(G168), .B(G1966), .Z(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1029 ( .A(KEYINPUT57), .B(n935), .Z(n936) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1031 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n962) );
  XOR2_X1 U1033 ( .A(G2090), .B(G35), .Z(n944) );
  XOR2_X1 U1034 ( .A(KEYINPUT54), .B(G34), .Z(n942) );
  XNOR2_X1 U1035 ( .A(G2084), .B(n942), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n958) );
  XNOR2_X1 U1037 ( .A(G1991), .B(G25), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(G33), .B(G2072), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n952) );
  XOR2_X1 U1040 ( .A(G2067), .B(G26), .Z(n947) );
  NAND2_X1 U1041 ( .A1(n947), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G32), .B(n948), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G27), .B(n953), .Z(n954) );
  NOR2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(n956), .B(KEYINPUT53), .ZN(n957) );
  NOR2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1049 ( .A(KEYINPUT55), .B(n959), .Z(n960) );
  NOR2_X1 U1050 ( .A1(G29), .A2(n960), .ZN(n961) );
  NOR2_X1 U1051 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n963), .ZN(n991) );
  XOR2_X1 U1053 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n988) );
  XOR2_X1 U1054 ( .A(G1966), .B(G21), .Z(n966) );
  XNOR2_X1 U1055 ( .A(n964), .B(G5), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n978) );
  XOR2_X1 U1057 ( .A(G1956), .B(G20), .Z(n970) );
  XNOR2_X1 U1058 ( .A(G1341), .B(G19), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G1981), .B(G6), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1062 ( .A(KEYINPUT122), .B(n971), .Z(n975) );
  XOR2_X1 U1063 ( .A(G4), .B(KEYINPUT123), .Z(n973) );
  XNOR2_X1 U1064 ( .A(G1348), .B(KEYINPUT59), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n973), .B(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(KEYINPUT60), .B(n976), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n986) );
  XOR2_X1 U1069 ( .A(G1986), .B(KEYINPUT124), .Z(n979) );
  XNOR2_X1 U1070 ( .A(G24), .B(n979), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(G1971), .B(G22), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G23), .B(G1976), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1075 ( .A(KEYINPUT58), .B(n984), .Z(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(n988), .B(n987), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n989), .ZN(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(KEYINPUT126), .B(n992), .ZN(n1020) );
  INV_X1 U1081 ( .A(n993), .ZN(n995) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n1003) );
  XNOR2_X1 U1083 ( .A(G160), .B(G2084), .ZN(n999) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1014) );
  XOR2_X1 U1088 ( .A(G2072), .B(n1004), .Z(n1006) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n1005) );
  NOR2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(KEYINPUT50), .B(n1007), .ZN(n1012) );
  XOR2_X1 U1092 ( .A(G2090), .B(G162), .Z(n1008) );
  NOR2_X1 U1093 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(KEYINPUT51), .B(n1010), .Z(n1011) );
  NAND2_X1 U1095 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1096 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1097 ( .A(KEYINPUT52), .B(n1015), .ZN(n1017) );
  INV_X1 U1098 ( .A(KEYINPUT55), .ZN(n1016) );
  NAND2_X1 U1099 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1100 ( .A1(n1018), .A2(G29), .ZN(n1019) );
  NAND2_X1 U1101 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1102 ( .A(n1021), .B(KEYINPUT62), .ZN(n1022) );
  XNOR2_X1 U1103 ( .A(KEYINPUT127), .B(n1022), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

