//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G107), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n189), .A2(new_n192), .A3(new_n193), .A4(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n191), .A2(G104), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n188), .A2(G107), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT78), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(KEYINPUT1), .A3(G146), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n207), .B(new_n208), .C1(G128), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n195), .A2(new_n198), .A3(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n200), .A2(KEYINPUT10), .A3(new_n210), .A4(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n214));
  OR2_X1    g028(.A1(new_n214), .A2(KEYINPUT10), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(KEYINPUT10), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n202), .A2(new_n204), .A3(new_n206), .ZN(new_n217));
  AOI21_X1  g031(.A(G128), .B1(new_n204), .B2(new_n206), .ZN(new_n218));
  INV_X1    g032(.A(new_n208), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n215), .B(new_n216), .C1(new_n220), .C2(new_n199), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n189), .A2(new_n192), .A3(new_n194), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n195), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT0), .B(G128), .Z(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n209), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n222), .A2(new_n229), .A3(G101), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n213), .A2(new_n221), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G134), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT11), .B1(new_n235), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n233), .A3(G134), .ZN(new_n238));
  AOI211_X1 g052(.A(G131), .B(new_n234), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(G137), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n232), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n213), .A2(new_n221), .A3(new_n231), .A4(new_n244), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT68), .B(G953), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G227), .ZN(new_n249));
  XNOR2_X1  g063(.A(G110), .B(G140), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n247), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n210), .B1(new_n200), .B2(new_n212), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n220), .A2(new_n199), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n245), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT79), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n244), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n195), .A2(new_n198), .A3(new_n211), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n211), .B1(new_n195), .B2(new_n198), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n220), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n199), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n210), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n245), .A3(new_n259), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n253), .B1(new_n261), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n252), .B1(new_n269), .B2(new_n251), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n187), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n247), .A2(new_n251), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT80), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n261), .A2(new_n268), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n247), .A2(new_n277), .A3(new_n251), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n246), .A2(new_n247), .ZN(new_n280));
  INV_X1    g094(.A(new_n251), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(G902), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n283), .A2(KEYINPUT81), .A3(new_n187), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT81), .B1(new_n283), .B2(new_n187), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n273), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT9), .B(G234), .ZN(new_n287));
  OAI21_X1  g101(.A(G221), .B1(new_n287), .B2(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G214), .B1(G237), .B2(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n228), .A2(G125), .ZN(new_n291));
  INV_X1    g105(.A(G125), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n210), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G224), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G953), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n296), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n291), .B2(new_n293), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT6), .ZN(new_n301));
  INV_X1    g115(.A(G119), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G116), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n304));
  INV_X1    g118(.A(G116), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(G119), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n302), .A2(KEYINPUT66), .A3(G116), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT2), .B(G113), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G113), .ZN(new_n312));
  INV_X1    g126(.A(G113), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(KEYINPUT2), .ZN(new_n314));
  OAI221_X1 g128(.A(new_n303), .B1(new_n312), .B2(new_n314), .C1(new_n306), .C2(new_n307), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n224), .A3(new_n230), .ZN(new_n317));
  OAI211_X1 g131(.A(KEYINPUT5), .B(new_n303), .C1(new_n306), .C2(new_n307), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n303), .A2(KEYINPUT5), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(G113), .A3(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n200), .A2(new_n320), .A3(new_n315), .A4(new_n212), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT82), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g138(.A(G110), .B(G122), .Z(new_n325));
  NAND3_X1  g139(.A1(new_n317), .A2(new_n321), .A3(KEYINPUT82), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n322), .A2(new_n325), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n301), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n317), .A2(new_n321), .A3(KEYINPUT82), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT82), .B1(new_n317), .B2(new_n321), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT6), .B1(new_n333), .B2(new_n325), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n300), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G210), .B1(G237), .B2(G902), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n296), .A2(KEYINPUT7), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n297), .A2(new_n299), .A3(new_n337), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n294), .A2(KEYINPUT7), .A3(new_n296), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n325), .B(KEYINPUT8), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n320), .A2(new_n315), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n199), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n341), .B1(new_n343), .B2(new_n321), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n328), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(G902), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n335), .A2(new_n336), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n336), .B1(new_n335), .B2(new_n346), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n290), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n290), .ZN(new_n352));
  INV_X1    g166(.A(new_n336), .ZN(new_n353));
  INV_X1    g167(.A(new_n300), .ZN(new_n354));
  INV_X1    g168(.A(new_n325), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n331), .A2(new_n332), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT6), .B1(new_n356), .B2(new_n328), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n327), .A2(new_n301), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n346), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n353), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n335), .A2(new_n336), .A3(new_n346), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n352), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT83), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n289), .B1(new_n351), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n248), .A2(G221), .A3(G234), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n366), .A2(G137), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(G137), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n367), .B2(new_n369), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT23), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n302), .B2(G128), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n374), .B(new_n375), .C1(G119), .C2(new_n201), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G110), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT72), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT16), .ZN(new_n380));
  INV_X1    g194(.A(G140), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G125), .ZN(new_n382));
  XOR2_X1   g196(.A(G125), .B(G140), .Z(new_n383));
  OAI211_X1 g197(.A(G146), .B(new_n382), .C1(new_n383), .C2(new_n380), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT73), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n292), .A2(new_n381), .ZN(new_n386));
  NAND2_X1  g200(.A1(G125), .A2(G140), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n382), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n203), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT73), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n389), .A2(new_n392), .A3(G146), .A4(new_n382), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT24), .B(G110), .Z(new_n395));
  XNOR2_X1  g209(.A(G119), .B(G128), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n379), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n388), .A2(KEYINPUT74), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT74), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(new_n386), .B2(new_n387), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n203), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n376), .A2(G110), .B1(new_n396), .B2(new_n395), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n384), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n372), .A2(new_n398), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n372), .B1(new_n398), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n271), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT25), .ZN(new_n408));
  INV_X1    g222(.A(G234), .ZN(new_n409));
  OAI21_X1  g223(.A(G217), .B1(new_n409), .B2(G902), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT71), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT25), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n412), .B(new_n271), .C1(new_n405), .C2(new_n406), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n408), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n405), .A2(new_n406), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n411), .A2(G902), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT76), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n228), .B1(new_n239), .B2(new_n243), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT65), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n233), .B2(G134), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n233), .A2(G134), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n242), .A2(new_n421), .ZN(new_n425));
  OAI21_X1  g239(.A(G131), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n241), .A2(new_n240), .A3(new_n242), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n210), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n420), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT30), .B1(new_n429), .B2(KEYINPUT64), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT64), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT30), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n431), .B(new_n432), .C1(new_n420), .C2(new_n428), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n316), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT67), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT67), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n436), .B(new_n316), .C1(new_n430), .C2(new_n433), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G237), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n248), .A2(G210), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT70), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n440), .A2(KEYINPUT70), .ZN(new_n444));
  INV_X1    g258(.A(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(KEYINPUT70), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT26), .B(G101), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n443), .A2(new_n447), .A3(new_n449), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n316), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n420), .A3(new_n428), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n438), .A2(KEYINPUT31), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n435), .A2(new_n454), .A3(new_n456), .A4(new_n437), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n429), .A2(new_n316), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n455), .B1(new_n420), .B2(new_n428), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT28), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT28), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT31), .B1(new_n464), .B2(new_n453), .ZN(new_n465));
  AOI21_X1  g279(.A(G902), .B1(new_n458), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G472), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n457), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT32), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT32), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n457), .A2(new_n466), .A3(new_n470), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n435), .A2(new_n456), .A3(new_n437), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n453), .ZN(new_n474));
  INV_X1    g288(.A(new_n464), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT29), .B1(new_n475), .B2(new_n454), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(KEYINPUT29), .A3(new_n454), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n271), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G472), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n419), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(KEYINPUT68), .A2(G953), .ZN(new_n482));
  NOR2_X1   g296(.A1(KEYINPUT68), .A2(G953), .ZN(new_n483));
  OAI211_X1 g297(.A(G214), .B(new_n439), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n205), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n248), .A2(G143), .A3(G214), .A4(new_n439), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G131), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT85), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n385), .A2(new_n391), .A3(new_n393), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n486), .A3(new_n240), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n240), .B1(new_n485), .B2(new_n486), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT17), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n490), .A2(new_n491), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G113), .B(G122), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n188), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT84), .B1(new_n388), .B2(new_n203), .ZN(new_n500));
  OR3_X1    g314(.A1(new_n388), .A2(KEYINPUT84), .A3(new_n203), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n402), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n485), .B(new_n486), .C1(new_n503), .C2(new_n240), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n502), .B(new_n504), .C1(new_n503), .C2(new_n488), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n497), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n499), .B1(new_n497), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n271), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G475), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n499), .A3(new_n505), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT19), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n399), .B2(new_n401), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n383), .A2(KEYINPUT19), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n203), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n492), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n514), .B(new_n384), .C1(new_n494), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n499), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n521), .B(KEYINPUT86), .Z(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(KEYINPUT20), .A3(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n509), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G953), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n528), .A2(G952), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n409), .B2(new_n439), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI211_X1 g345(.A(new_n271), .B(new_n248), .C1(G234), .C2(G237), .ZN(new_n532));
  XOR2_X1   g346(.A(KEYINPUT21), .B(G898), .Z(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n205), .A2(G128), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n201), .A2(G143), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G134), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n235), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G122), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G116), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n305), .A2(G122), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G107), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n305), .A2(KEYINPUT14), .A3(G122), .ZN(new_n548));
  OAI211_X1 g362(.A(G107), .B(new_n548), .C1(new_n545), .C2(KEYINPUT14), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n541), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT13), .ZN(new_n551));
  OR3_X1    g365(.A1(new_n201), .A2(KEYINPUT13), .A3(G143), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(G134), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n191), .B1(new_n543), .B2(new_n544), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n553), .B(new_n540), .C1(new_n546), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n287), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(G217), .A3(new_n528), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT87), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n556), .A2(new_n558), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n556), .A2(KEYINPUT87), .A3(new_n558), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n271), .ZN(new_n565));
  INV_X1    g379(.A(G478), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n565), .B(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n527), .A2(new_n535), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n365), .A2(new_n481), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  INV_X1    g385(.A(KEYINPUT90), .ZN(new_n572));
  INV_X1    g386(.A(new_n535), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n573), .B(new_n290), .C1(new_n347), .C2(new_n348), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n556), .A2(KEYINPUT88), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n558), .ZN(new_n577));
  INV_X1    g391(.A(new_n558), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n556), .A2(KEYINPUT88), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n575), .B2(new_n564), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT89), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n581), .A2(new_n582), .A3(G478), .A4(new_n271), .ZN(new_n583));
  INV_X1    g397(.A(new_n579), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n578), .B1(new_n556), .B2(KEYINPUT88), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT33), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT87), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n587), .B(new_n578), .C1(new_n550), .C2(new_n555), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n559), .A2(new_n588), .A3(new_n561), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n586), .B(G478), .C1(new_n589), .C2(KEYINPUT33), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT89), .B1(new_n590), .B2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n565), .A2(new_n566), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n583), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n527), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n572), .B1(new_n574), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n596), .A2(new_n363), .A3(KEYINPUT90), .A4(new_n573), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n288), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n419), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n457), .A2(new_n466), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G472), .ZN(new_n602));
  AND4_X1   g416(.A1(new_n468), .A2(new_n286), .A3(new_n600), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT34), .B(G104), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G6));
  AND3_X1   g420(.A1(new_n509), .A2(new_n525), .A3(new_n526), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n568), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n574), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G107), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  NOR2_X1   g426(.A1(new_n372), .A2(KEYINPUT36), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n398), .A2(new_n404), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n417), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n414), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n602), .A2(new_n468), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT91), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT91), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n602), .A2(new_n620), .A3(new_n468), .A4(new_n617), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n365), .A2(new_n569), .A3(new_n619), .A4(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT37), .B(G110), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G12));
  INV_X1    g438(.A(new_n617), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n472), .B2(new_n480), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n279), .A2(new_n282), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n187), .A3(new_n271), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT81), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n283), .A2(KEYINPUT81), .A3(new_n187), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n599), .B1(new_n632), .B2(new_n273), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT92), .B(G900), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n531), .B1(new_n532), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n608), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n626), .A2(new_n633), .A3(new_n363), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  NAND2_X1  g452(.A1(new_n361), .A2(new_n362), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT94), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n527), .A2(new_n568), .A3(new_n290), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n635), .B(KEYINPUT39), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n633), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT95), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT40), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n648), .B(KEYINPUT95), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n473), .A2(new_n454), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n459), .A2(new_n460), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(G902), .B1(new_n656), .B2(new_n453), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n467), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n469), .B2(new_n471), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n617), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n645), .A2(new_n650), .A3(new_n653), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n205), .ZN(G45));
  INV_X1    g476(.A(new_n635), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n593), .A2(new_n527), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n626), .A2(new_n633), .A3(new_n363), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  OR2_X1    g481(.A1(new_n283), .A2(new_n187), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n288), .B(new_n668), .C1(new_n284), .C2(new_n285), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT96), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n283), .A2(new_n187), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n630), .B2(new_n631), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT96), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n673), .A3(new_n288), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n598), .A2(new_n481), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT41), .B(G113), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  NAND3_X1  g492(.A1(new_n481), .A2(new_n675), .A3(new_n609), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  INV_X1    g494(.A(KEYINPUT97), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n669), .B2(new_n349), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n363), .A2(new_n672), .A3(KEYINPUT97), .A4(new_n288), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n569), .A3(new_n626), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT98), .B(G119), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G21));
  NAND2_X1  g501(.A1(new_n643), .A2(new_n639), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n535), .ZN(new_n689));
  INV_X1    g503(.A(new_n419), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n458), .A2(new_n465), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n271), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT31), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n458), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n691), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n602), .A2(new_n696), .A3(new_n468), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n601), .A2(new_n691), .A3(G472), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n675), .A2(new_n689), .A3(new_n690), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT100), .B(G122), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G24));
  NAND2_X1  g516(.A1(new_n664), .A2(KEYINPUT101), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n593), .A2(new_n527), .A3(new_n704), .A4(new_n663), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n697), .A2(new_n698), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n684), .A2(new_n706), .A3(new_n617), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G125), .ZN(G27));
  NOR2_X1   g522(.A1(new_n639), .A2(new_n352), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n267), .A2(new_n245), .A3(new_n259), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n259), .B1(new_n267), .B2(new_n245), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n247), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n281), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n187), .A2(KEYINPUT102), .A3(G902), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n252), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n716), .B1(new_n272), .B2(new_n717), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n710), .B(new_n599), .C1(new_n632), .C2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n284), .B2(new_n285), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT103), .B1(new_n720), .B2(new_n288), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n709), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n472), .A2(new_n480), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n703), .A2(new_n705), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n690), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT104), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n709), .ZN(new_n727));
  AOI21_X1  g541(.A(G902), .B1(new_n714), .B2(new_n252), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT102), .B1(new_n728), .B2(new_n187), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n630), .A2(new_n631), .B1(new_n729), .B2(new_n716), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n710), .B1(new_n730), .B2(new_n599), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n720), .A2(KEYINPUT103), .A3(new_n288), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n481), .A4(new_n724), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n726), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n733), .A2(KEYINPUT42), .A3(new_n481), .A4(new_n724), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n726), .A2(new_n735), .A3(new_n740), .A4(new_n736), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  OAI211_X1 g557(.A(new_n636), .B(new_n709), .C1(new_n719), .C2(new_n721), .ZN(new_n744));
  INV_X1    g558(.A(new_n481), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT106), .B(G134), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G36));
  NAND2_X1  g562(.A1(new_n607), .A2(new_n593), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT108), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n753), .B2(new_n749), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(KEYINPUT109), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n754), .A2(KEYINPUT109), .B1(new_n468), .B2(new_n602), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n756), .A3(new_n617), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n727), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n270), .B(KEYINPUT45), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n761), .B(G469), .C1(new_n762), .C2(G902), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(G469), .ZN(new_n764));
  NAND2_X1  g578(.A1(G469), .A2(G902), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n632), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n288), .A3(new_n647), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n757), .B2(new_n758), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n760), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  NAND2_X1  g585(.A1(new_n767), .A2(new_n288), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT47), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n723), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n727), .A2(new_n690), .A3(new_n664), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  AND2_X1   g592(.A1(new_n754), .A2(new_n531), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n727), .A2(new_n669), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n481), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT48), .ZN(new_n782));
  INV_X1    g596(.A(new_n699), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n419), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n684), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n529), .A3(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n642), .A2(new_n352), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n779), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n669), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT50), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(KEYINPUT50), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n790), .A2(new_n791), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n779), .A2(new_n784), .A3(new_n789), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n792), .B(KEYINPUT50), .C1(new_n796), .C2(new_n669), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n690), .A2(new_n780), .A3(new_n531), .A4(new_n659), .ZN(new_n799));
  INV_X1    g613(.A(new_n593), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n607), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n754), .A2(new_n531), .A3(new_n617), .A4(new_n780), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n783), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n798), .A2(new_n806), .A3(KEYINPUT116), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n672), .A2(new_n599), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n727), .B1(new_n773), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n786), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n795), .A2(new_n804), .A3(new_n797), .A4(new_n805), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n807), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT51), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n803), .B1(new_n786), .B2(new_n809), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n798), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n788), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n799), .A2(new_n596), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n676), .A2(new_n685), .A3(new_n700), .A4(new_n679), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n363), .A2(KEYINPUT83), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n350), .B(new_n352), .C1(new_n361), .C2(new_n362), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n569), .B(new_n633), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n619), .A2(new_n621), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n745), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n351), .A2(new_n364), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n608), .A2(new_n594), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n573), .A2(new_n603), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n823), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n603), .A2(new_n829), .A3(new_n573), .A4(new_n830), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n622), .A2(new_n570), .A3(KEYINPUT111), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n822), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n706), .B1(new_n721), .B2(new_n719), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n527), .A2(new_n568), .A3(new_n635), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n723), .A2(new_n633), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n625), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n746), .B1(new_n839), .B2(new_n709), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n720), .A2(new_n288), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n659), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT112), .B1(new_n617), .B2(new_n635), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n414), .A2(new_n616), .A3(new_n844), .A4(new_n663), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n639), .A2(new_n843), .A3(new_n643), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n842), .A2(KEYINPUT113), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT113), .B1(new_n842), .B2(new_n846), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n707), .A2(new_n637), .A3(new_n666), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n707), .A2(new_n637), .A3(new_n666), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n842), .A2(new_n846), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n847), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n835), .B(new_n840), .C1(new_n853), .C2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n821), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n832), .A2(new_n834), .ZN(new_n863));
  INV_X1    g677(.A(new_n822), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n863), .A2(new_n864), .A3(new_n840), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n852), .B1(new_n850), .B2(new_n851), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n854), .A2(KEYINPUT52), .A3(new_n858), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n742), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT54), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n862), .A2(KEYINPUT54), .A3(new_n869), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n819), .B(new_n820), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(G952), .B2(G953), .ZN(new_n873));
  INV_X1    g687(.A(new_n672), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n607), .B(new_n593), .C1(new_n874), .C2(KEYINPUT49), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(KEYINPUT49), .B2(new_n874), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n600), .A2(new_n290), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT110), .Z(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n878), .A3(new_n642), .A4(new_n659), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(G75));
  AOI21_X1  g694(.A(new_n271), .B1(new_n862), .B2(new_n869), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT56), .B1(new_n881), .B2(G210), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n330), .A2(new_n334), .A3(new_n300), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n359), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT55), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n882), .A2(new_n885), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n248), .A2(G952), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G51));
  XOR2_X1   g703(.A(new_n765), .B(KEYINPUT57), .Z(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n871), .A2(new_n870), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n627), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT117), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n881), .A2(G469), .A3(new_n762), .ZN(new_n895));
  INV_X1    g709(.A(new_n870), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n862), .A2(KEYINPUT54), .A3(new_n869), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n897), .A3(new_n890), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT117), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n899), .A3(new_n627), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n894), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n888), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n901), .A2(KEYINPUT118), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(new_n520), .Z(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n888), .ZN(G60));
  NAND2_X1  g724(.A1(G478), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT59), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n896), .A2(new_n897), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n581), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT119), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT119), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n888), .B(new_n915), .C1(new_n917), .C2(new_n918), .ZN(G63));
  NAND2_X1  g733(.A1(new_n862), .A2(new_n869), .ZN(new_n920));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT60), .Z(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT120), .ZN(new_n924));
  INV_X1    g738(.A(new_n415), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n923), .B(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n615), .B(KEYINPUT121), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n926), .A2(new_n930), .A3(new_n902), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n926), .A2(new_n930), .A3(KEYINPUT61), .A4(new_n902), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(G66));
  INV_X1    g749(.A(new_n835), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n528), .B1(new_n533), .B2(G224), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n936), .A2(new_n248), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n357), .B(new_n358), .C1(G898), .C2(new_n248), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G69));
  INV_X1    g756(.A(new_n777), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n760), .B2(new_n769), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n744), .B1(new_n768), .B2(new_n688), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n851), .B1(new_n945), .B2(new_n481), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n742), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n944), .A2(KEYINPUT124), .A3(new_n742), .A4(new_n946), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n949), .A2(new_n248), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n430), .A2(new_n433), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n512), .A2(new_n513), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(G900), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n951), .B(new_n954), .C1(new_n955), .C2(new_n248), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n661), .A2(new_n851), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  INV_X1    g772(.A(new_n648), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n959), .A2(new_n481), .A3(new_n709), .A4(new_n830), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT123), .Z(new_n961));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n944), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n962), .A2(new_n248), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(new_n954), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n248), .B1(G227), .B2(G900), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n956), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n956), .B2(new_n964), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(G72));
  XNOR2_X1  g782(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n467), .A2(new_n271), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n962), .B2(new_n936), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n974), .B(new_n971), .C1(new_n962), .C2(new_n936), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n971), .B1(new_n474), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n474), .A2(new_n977), .A3(new_n458), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n920), .A2(new_n979), .ZN(new_n980));
  OAI22_X1  g794(.A1(new_n976), .A2(new_n654), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n949), .A2(new_n835), .A3(new_n950), .ZN(new_n982));
  AOI211_X1 g796(.A(new_n454), .B(new_n473), .C1(new_n982), .C2(new_n971), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n981), .A2(new_n983), .A3(new_n888), .ZN(G57));
endmodule


