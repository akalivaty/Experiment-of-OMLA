//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  NAND2_X1  g002(.A1(G234), .A2(G237), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT21), .B(G898), .Z(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(G902), .A3(G953), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT67), .A2(G116), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT67), .A2(G116), .ZN(new_n195));
  OAI21_X1  g009(.A(G119), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G116), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT2), .A2(G113), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT2), .A2(G113), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n198), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT68), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n196), .A2(new_n204), .A3(new_n201), .A4(new_n198), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n206), .A2(G113), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n196), .A2(KEYINPUT5), .A3(new_n198), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n203), .A2(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G104), .B(G107), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT84), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT84), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G101), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n213), .B2(G104), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n221), .A2(new_n214), .B1(new_n222), .B2(new_n213), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT82), .B(G101), .Z(new_n224));
  AOI22_X1  g038(.A1(new_n212), .A2(new_n219), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n220), .A2(new_n213), .A3(G104), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n215), .A2(G107), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT83), .A2(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n221), .A2(new_n214), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n224), .A2(new_n233), .A3(new_n227), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT4), .B1(new_n230), .B2(new_n231), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n196), .A2(new_n198), .ZN(new_n238));
  INV_X1    g052(.A(new_n201), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n203), .A2(new_n205), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n226), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(G110), .B(G122), .Z(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(KEYINPUT90), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT90), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n203), .A2(new_n205), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n239), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n230), .A2(new_n231), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n234), .A3(new_n232), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n247), .A2(new_n251), .B1(new_n209), .B2(new_n225), .ZN(new_n252));
  INV_X1    g066(.A(new_n242), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n244), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n253), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n243), .A2(new_n254), .A3(KEYINPUT6), .A4(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT91), .B(KEYINPUT6), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n237), .A2(new_n240), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n207), .A2(new_n208), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n245), .A2(new_n225), .A3(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n242), .B(new_n257), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT92), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n241), .A2(KEYINPUT92), .A3(new_n242), .A4(new_n257), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G143), .B(G146), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT0), .A3(G128), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G128), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n267), .B(G125), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n270));
  NOR2_X1   g084(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n271));
  OAI21_X1  g085(.A(G128), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n266), .ZN(new_n273));
  INV_X1    g087(.A(G146), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G143), .ZN(new_n275));
  INV_X1    g089(.A(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G146), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G128), .ZN(new_n279));
  INV_X1    g093(.A(new_n277), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n270), .A2(new_n271), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n273), .A2(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n269), .B1(new_n282), .B2(G125), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n187), .A2(G224), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n256), .A2(new_n265), .A3(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n242), .B(KEYINPUT8), .Z(new_n287));
  NOR2_X1   g101(.A1(new_n209), .A2(new_n225), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(new_n260), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n284), .A2(KEYINPUT7), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n283), .B(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n255), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT93), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT93), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n296), .A3(new_n293), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n286), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  XOR2_X1   g113(.A(new_n299), .B(KEYINPUT94), .Z(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G214), .B1(G237), .B2(G902), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n286), .A2(new_n295), .A3(new_n300), .A4(new_n297), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n193), .B1(new_n306), .B2(KEYINPUT95), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT95), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G472), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n273), .A2(new_n279), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n281), .A2(new_n280), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT65), .B(G137), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT11), .ZN(new_n317));
  INV_X1    g131(.A(G134), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n316), .A2(new_n319), .B1(new_n318), .B2(G137), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n317), .B1(new_n318), .B2(G137), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT64), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT64), .B(new_n317), .C1(new_n318), .C2(G137), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G137), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n316), .B2(G134), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G131), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n315), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n267), .B1(new_n266), .B2(new_n268), .ZN(new_n333));
  INV_X1    g147(.A(new_n324), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT64), .B1(new_n329), .B2(new_n317), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(KEYINPUT65), .A2(G137), .ZN(new_n337));
  AND2_X1   g151(.A1(KEYINPUT65), .A2(G137), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n319), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n318), .A2(G137), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G131), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n333), .B1(new_n342), .B2(new_n327), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n312), .B1(new_n332), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n333), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n320), .A2(new_n326), .A3(new_n325), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n326), .B1(new_n320), .B2(new_n325), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n315), .A2(new_n327), .A3(new_n331), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(KEYINPUT30), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n344), .A2(new_n247), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n240), .A3(new_n349), .ZN(new_n352));
  INV_X1    g166(.A(G237), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT69), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT69), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G237), .ZN(new_n356));
  AOI21_X1  g170(.A(G953), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G210), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT26), .B(G101), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n351), .A2(new_n352), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT31), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n351), .A2(new_n365), .A3(new_n352), .A4(new_n362), .ZN(new_n366));
  INV_X1    g180(.A(new_n362), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n247), .B1(new_n332), .B2(new_n343), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n352), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n352), .A2(new_n368), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n367), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n364), .A2(new_n366), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT71), .B1(new_n363), .B2(KEYINPUT31), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n311), .B(new_n293), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT32), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n348), .A2(new_n240), .A3(new_n349), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n240), .B1(new_n348), .B2(new_n349), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT28), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n381), .A2(KEYINPUT29), .A3(new_n362), .A4(new_n371), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n293), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT73), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT73), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n385), .A3(new_n293), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n351), .A2(new_n352), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n367), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n370), .A2(new_n372), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n388), .A2(KEYINPUT72), .B1(new_n389), .B2(new_n362), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n381), .A2(KEYINPUT72), .A3(new_n362), .A4(new_n371), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n384), .B(new_n386), .C1(new_n390), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G472), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n363), .A2(KEYINPUT31), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT71), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n398), .A2(new_n364), .A3(new_n366), .A4(new_n373), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n399), .A2(KEYINPUT32), .A3(new_n311), .A4(new_n293), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n378), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT77), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT22), .B(G137), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT16), .ZN(new_n406));
  INV_X1    g220(.A(G140), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(G125), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(G125), .ZN(new_n409));
  INV_X1    g223(.A(G125), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n408), .B1(new_n412), .B2(new_n406), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n274), .ZN(new_n414));
  OAI211_X1 g228(.A(G146), .B(new_n408), .C1(new_n412), .C2(new_n406), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(KEYINPUT75), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT74), .B1(new_n197), .B2(G128), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n417), .A2(KEYINPUT23), .B1(new_n197), .B2(G128), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT23), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT74), .B(new_n419), .C1(new_n197), .C2(G128), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G119), .B(G128), .ZN(new_n422));
  XOR2_X1   g236(.A(KEYINPUT24), .B(G110), .Z(new_n423));
  AOI22_X1  g237(.A1(new_n421), .A2(G110), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n413), .A2(new_n425), .A3(new_n274), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n416), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  OAI22_X1  g241(.A1(new_n421), .A2(G110), .B1(new_n422), .B2(new_n423), .ZN(new_n428));
  XNOR2_X1  g242(.A(G125), .B(G140), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n274), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT76), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n432), .A3(new_n415), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT78), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n427), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n427), .B2(new_n433), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n405), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n427), .A2(new_n433), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT78), .ZN(new_n439));
  INV_X1    g253(.A(new_n405), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n293), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT79), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT25), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G217), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(G234), .B2(new_n293), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n442), .A2(new_n444), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n437), .A2(KEYINPUT25), .A3(new_n441), .A4(new_n293), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n437), .A2(new_n441), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT80), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n447), .A2(G902), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n449), .A2(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n401), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT9), .B(G234), .Z(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G221), .B1(new_n460), .B2(G902), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G469), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n187), .A2(G227), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT81), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G140), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n342), .A2(new_n327), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT10), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n313), .B2(new_n314), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n251), .A2(new_n345), .B1(new_n472), .B2(new_n225), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n218), .B1(new_n217), .B2(G101), .ZN(new_n475));
  AOI211_X1 g289(.A(KEYINPUT84), .B(new_n211), .C1(new_n214), .C2(new_n216), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n234), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n280), .A2(KEYINPUT1), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n273), .B2(new_n279), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n474), .B(new_n471), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n212), .A2(new_n219), .ZN(new_n482));
  INV_X1    g296(.A(G128), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n275), .B2(new_n277), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n266), .B2(new_n272), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n482), .B(new_n234), .C1(new_n485), .C2(new_n478), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n474), .B1(new_n486), .B2(new_n471), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n470), .B(new_n473), .C1(new_n481), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n477), .A2(new_n479), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT85), .B1(new_n491), .B2(KEYINPUT10), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n480), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n493), .A2(KEYINPUT86), .A3(new_n470), .A4(new_n473), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n468), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n486), .B1(new_n315), .B2(new_n225), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT87), .A3(new_n469), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT12), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n345), .B1(new_n235), .B2(new_n236), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n315), .A2(new_n225), .A3(KEYINPUT10), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n492), .B2(new_n480), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT88), .B1(new_n504), .B2(new_n470), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n473), .B1(new_n481), .B2(new_n487), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n469), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n490), .A2(new_n494), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n467), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n500), .B1(new_n511), .B2(KEYINPUT89), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n505), .A2(new_n508), .B1(new_n490), .B2(new_n494), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n513), .A2(new_n514), .A3(new_n467), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n463), .B(new_n293), .C1(new_n512), .C2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n463), .A2(new_n293), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n510), .A2(new_n499), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n518), .A2(new_n468), .B1(new_n495), .B2(new_n509), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n519), .B2(G469), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n462), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT96), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n355), .A2(G237), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n353), .A2(KEYINPUT69), .ZN(new_n525));
  OAI211_X1 g339(.A(G214), .B(new_n187), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n276), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n357), .A2(G143), .A3(G214), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n523), .B1(new_n529), .B2(G131), .ZN(new_n530));
  AOI211_X1 g344(.A(KEYINPUT96), .B(new_n326), .C1(new_n527), .C2(new_n528), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT17), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT98), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n416), .A2(new_n426), .ZN(new_n535));
  INV_X1    g349(.A(new_n530), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n537));
  INV_X1    g351(.A(new_n529), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n326), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n529), .A2(new_n523), .A3(G131), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT98), .B(KEYINPUT17), .C1(new_n530), .C2(new_n531), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n534), .A2(new_n535), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(G113), .B(G122), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT97), .B(G104), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n538), .B1(new_n547), .B2(new_n326), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n432), .B1(new_n274), .B2(new_n429), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n529), .A2(G131), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(new_n547), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n543), .A2(new_n546), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n546), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n412), .B(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n415), .B1(new_n557), .B2(G146), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n530), .A2(new_n531), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n559), .B2(new_n539), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n556), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G475), .A2(G902), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n522), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n563), .ZN(new_n565));
  AOI211_X1 g379(.A(KEYINPUT20), .B(new_n565), .C1(new_n555), .C2(new_n561), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n543), .A2(new_n554), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n556), .ZN(new_n568));
  AOI21_X1  g382(.A(G902), .B1(new_n568), .B2(new_n555), .ZN(new_n569));
  INV_X1    g383(.A(G475), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n564), .A2(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT67), .B(G116), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G122), .ZN(new_n573));
  INV_X1    g387(.A(G116), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT99), .B(G122), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n213), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT13), .B1(new_n483), .B2(G143), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n318), .ZN(new_n579));
  XNOR2_X1  g393(.A(G128), .B(G143), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n573), .B(G107), .C1(new_n574), .C2(new_n575), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(KEYINPUT14), .B(G107), .C1(new_n575), .C2(new_n574), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n577), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n580), .B(new_n318), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n576), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n460), .A2(new_n446), .A3(G953), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n590), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n588), .A2(KEYINPUT100), .A3(new_n590), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n293), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G478), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(KEYINPUT15), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n571), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n310), .A2(new_n458), .A3(new_n521), .A4(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT101), .B(KEYINPUT102), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n224), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n601), .B(new_n603), .ZN(G3));
  OAI21_X1  g418(.A(new_n293), .B1(new_n374), .B2(new_n375), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G472), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n606), .A2(new_n376), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n521), .A2(new_n456), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n521), .A2(KEYINPUT103), .A3(new_n456), .A4(new_n607), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n193), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n594), .A2(new_n615), .A3(new_n595), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n591), .A2(KEYINPUT33), .A3(new_n593), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(G478), .A3(new_n293), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n596), .A2(new_n597), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n613), .A2(new_n614), .A3(new_n571), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n571), .A2(new_n620), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT104), .B1(new_n622), .B2(new_n612), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n610), .A2(new_n611), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  INV_X1    g441(.A(new_n599), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n612), .A2(new_n628), .A3(new_n571), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n610), .A2(new_n611), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n405), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n438), .B(new_n633), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n449), .A2(new_n452), .B1(new_n455), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n635), .A2(new_n571), .A3(new_n599), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n310), .A2(new_n521), .A3(new_n607), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  NAND2_X1  g453(.A1(new_n562), .A2(new_n563), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT20), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n562), .A2(new_n522), .A3(new_n563), .ZN(new_n642));
  INV_X1    g456(.A(new_n555), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n546), .B1(new_n543), .B2(new_n554), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n293), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n641), .A2(new_n642), .B1(G475), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n190), .B(KEYINPUT105), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(G900), .B2(new_n192), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n646), .A2(new_n599), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n305), .A2(new_n635), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n650), .A2(new_n521), .A3(new_n401), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XOR2_X1   g467(.A(new_n649), .B(KEYINPUT39), .Z(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n521), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n367), .B1(new_n379), .B2(new_n380), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(G472), .A3(new_n363), .ZN(new_n661));
  NAND2_X1  g475(.A1(G472), .A2(G902), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT108), .Z(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n378), .A3(new_n400), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n635), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n302), .A2(new_n304), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT107), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n667), .B(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n303), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n571), .A2(new_n599), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n666), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n658), .A2(new_n659), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n276), .ZN(G45));
  NAND3_X1  g489(.A1(new_n571), .A2(new_n620), .A3(new_n649), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n521), .A2(new_n677), .A3(new_n401), .A4(new_n651), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  NAND2_X1  g493(.A1(new_n509), .A2(new_n510), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(KEYINPUT89), .A3(new_n468), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n514), .B1(new_n513), .B2(new_n467), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n500), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n293), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n461), .A3(new_n516), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n457), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n624), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n629), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NOR2_X1   g506(.A1(new_n686), .A2(new_n305), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(new_n401), .A3(new_n193), .A4(new_n636), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  NAND3_X1  g509(.A1(new_n396), .A2(new_n366), .A3(new_n373), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n311), .A3(new_n293), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n606), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n456), .A3(new_n193), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n686), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n646), .B2(new_n628), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n571), .A2(new_n599), .A3(KEYINPUT109), .ZN(new_n703));
  AND4_X1   g517(.A1(KEYINPUT110), .A2(new_n702), .A3(new_n306), .A4(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n305), .B1(new_n672), .B2(new_n701), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT110), .B1(new_n705), .B2(new_n703), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n700), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  AND3_X1   g522(.A1(new_n683), .A2(new_n463), .A3(new_n293), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n463), .B1(new_n683), .B2(new_n293), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n709), .A2(new_n710), .A3(new_n462), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n634), .A2(new_n455), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n451), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n712), .B1(new_n713), .B2(new_n448), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n606), .A2(new_n714), .A3(new_n697), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n676), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n711), .A2(new_n716), .A3(new_n306), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT111), .B(G125), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G27));
  XOR2_X1   g533(.A(KEYINPUT112), .B(KEYINPUT42), .Z(new_n720));
  AOI21_X1  g534(.A(new_n671), .B1(new_n302), .B2(new_n304), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n521), .A2(new_n456), .A3(new_n401), .A4(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n720), .B1(new_n722), .B2(new_n676), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n516), .A2(new_n520), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n721), .A3(new_n461), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n457), .A3(new_n676), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n723), .A2(new_n724), .B1(new_n727), .B2(KEYINPUT42), .ZN(new_n728));
  OAI211_X1 g542(.A(KEYINPUT113), .B(new_n720), .C1(new_n722), .C2(new_n676), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G131), .ZN(G33));
  INV_X1    g545(.A(new_n722), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n650), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(KEYINPUT114), .A3(new_n650), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  NAND2_X1  g552(.A1(new_n646), .A2(new_n620), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n646), .A2(KEYINPUT43), .A3(new_n620), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n607), .A2(new_n635), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT44), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n519), .A2(KEYINPUT45), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n519), .A2(KEYINPUT45), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(G469), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n517), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n516), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT46), .B1(new_n749), .B2(new_n750), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n461), .B(new_n655), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n743), .A2(KEYINPUT44), .A3(new_n744), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n746), .A2(new_n721), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT115), .B(G137), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G39));
  OAI21_X1  g573(.A(new_n461), .B1(new_n752), .B2(new_n753), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(KEYINPUT116), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n456), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n721), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n765), .A2(new_n401), .A3(new_n676), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n761), .A2(KEYINPUT116), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n760), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n763), .B(new_n766), .C1(new_n768), .C2(new_n762), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  NOR2_X1   g584(.A1(new_n709), .A2(new_n710), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT49), .ZN(new_n772));
  INV_X1    g586(.A(new_n670), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n456), .A2(new_n461), .A3(new_n303), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n774), .A3(new_n739), .ZN(new_n775));
  INV_X1    g589(.A(new_n665), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n772), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n711), .A2(new_n721), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n648), .B1(new_n741), .B2(new_n742), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n714), .A3(new_n698), .A4(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n665), .A2(new_n764), .A3(new_n190), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n646), .A3(new_n619), .A4(new_n618), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n780), .A2(new_n456), .A3(new_n698), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n773), .A2(new_n686), .A3(new_n303), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(KEYINPUT50), .A3(new_n786), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n789), .A2(KEYINPUT117), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT117), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n781), .B(new_n784), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n771), .A2(new_n462), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n768), .A2(new_n762), .ZN(new_n795));
  INV_X1    g609(.A(new_n763), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n785), .A2(new_n721), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n778), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n779), .A2(new_n782), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n188), .B1(new_n801), .B2(new_n622), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n785), .A2(new_n693), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT119), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT119), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n779), .A2(new_n780), .A3(new_n458), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT48), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT120), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n797), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(KEYINPUT118), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n798), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n784), .A2(new_n781), .A3(KEYINPUT51), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n789), .B2(new_n790), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n806), .A2(new_n818), .A3(new_n808), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n800), .A2(new_n810), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n636), .A2(new_n401), .A3(new_n721), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n521), .A2(new_n649), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n725), .A2(new_n721), .A3(new_n461), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n716), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n687), .B1(new_n624), .B2(new_n629), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n707), .A2(new_n824), .A3(new_n825), .A4(new_n694), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n610), .A2(new_n611), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n622), .B1(new_n628), .B2(new_n571), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n310), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n601), .B(new_n637), .C1(new_n827), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n728), .A2(new_n729), .B1(new_n735), .B2(new_n736), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n717), .A2(new_n652), .A3(new_n678), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n521), .A2(new_n665), .A3(new_n635), .A4(new_n649), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n704), .B2(new_n706), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n836), .A3(KEYINPUT52), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n702), .A2(new_n306), .A3(new_n703), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n705), .A2(KEYINPUT110), .A3(new_n703), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n834), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n717), .A2(new_n652), .A3(new_n678), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n837), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n831), .A2(new_n832), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n831), .A2(new_n832), .A3(new_n846), .A4(KEYINPUT53), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n820), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(G952), .A2(G953), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n777), .B1(new_n856), .B2(new_n857), .ZN(G75));
  NAND3_X1  g672(.A1(new_n851), .A2(G902), .A3(new_n300), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n256), .A2(new_n265), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(new_n285), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT55), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n187), .A2(G952), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n293), .B1(new_n849), .B2(new_n850), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n869), .B2(new_n300), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n860), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n864), .B1(new_n870), .B2(new_n860), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(G51));
  XNOR2_X1  g687(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n517), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n855), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n683), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n749), .B(KEYINPUT123), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n869), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n866), .B1(new_n877), .B2(new_n879), .ZN(G54));
  NAND3_X1  g694(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .ZN(new_n881));
  INV_X1    g695(.A(new_n562), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n867), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT124), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n886), .A3(new_n882), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(G60));
  AND2_X1   g702(.A1(new_n616), .A2(new_n617), .ZN(new_n889));
  NAND2_X1  g703(.A1(G478), .A2(G902), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT59), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n855), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n867), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n889), .B1(new_n855), .B2(new_n891), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(G63));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n896));
  XNOR2_X1  g710(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n446), .A2(new_n293), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n851), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n454), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n867), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n634), .B(KEYINPUT126), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n896), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n866), .B1(new_n900), .B2(new_n901), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n907), .B(KEYINPUT61), .C1(new_n900), .C2(new_n904), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(G66));
  NAND2_X1  g723(.A1(new_n191), .A2(G224), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G953), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n707), .A2(new_n694), .A3(new_n825), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n830), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n915), .A3(new_n187), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n914), .B2(new_n187), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n911), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n862), .B1(G898), .B2(new_n187), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  NAND2_X1  g735(.A1(G900), .A2(G953), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n755), .B(new_n458), .C1(new_n706), .C2(new_n704), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n757), .A2(new_n769), .A3(new_n833), .A4(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n832), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n923), .B1(new_n927), .B2(new_n187), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n344), .A2(new_n350), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n557), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n674), .A2(new_n844), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n656), .A2(new_n458), .A3(new_n721), .A4(new_n828), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n757), .A2(new_n769), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n931), .A2(new_n187), .ZN(new_n938));
  OAI22_X1  g752(.A1(new_n928), .A2(new_n931), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(G227), .A2(G900), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(G953), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G72));
  NAND2_X1  g756(.A1(new_n388), .A2(new_n363), .ZN(new_n943));
  INV_X1    g757(.A(new_n387), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n925), .B2(new_n926), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n913), .B(new_n945), .C1(new_n937), .C2(new_n944), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n662), .B(KEYINPUT63), .Z(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n851), .A2(new_n943), .A3(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n866), .A3(new_n949), .ZN(G57));
endmodule


