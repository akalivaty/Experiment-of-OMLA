//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1174, new_n1175, new_n1176,
    new_n1178, new_n1179, new_n1180, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT66), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n211), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n235), .A2(new_n209), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n231), .B(new_n237), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n227), .A2(new_n238), .ZN(G361));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G238), .B(G244), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT2), .B(G226), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n243), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XOR2_X1   g0051(.A(new_n251), .B(KEYINPUT68), .Z(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G68), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G58), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  AOI21_X1  g0056(.A(new_n235), .B1(G33), .B2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G222), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(G1698), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n265), .B1(new_n219), .B2(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n258), .B1(new_n269), .B2(KEYINPUT70), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(KEYINPUT70), .B2(new_n269), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n208), .A2(G274), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT69), .B(G45), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n257), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(G226), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT74), .B1(new_n280), .B2(G169), .ZN(new_n281));
  INV_X1    g0081(.A(G179), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n202), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n235), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n208), .B2(G20), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n289), .B2(new_n202), .ZN(new_n290));
  XOR2_X1   g0090(.A(new_n290), .B(KEYINPUT73), .Z(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT8), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G58), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT72), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT71), .B(G58), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n294), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n209), .A2(G33), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n293), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n288), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT74), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n284), .B(new_n303), .C1(new_n304), .C2(new_n283), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n280), .A2(G190), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n280), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n303), .A2(new_n306), .ZN(new_n310));
  XOR2_X1   g0110(.A(new_n310), .B(KEYINPUT77), .Z(new_n311));
  NOR2_X1   g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT10), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n305), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n266), .A2(G232), .A3(G1698), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G97), .ZN(new_n318));
  INV_X1    g0118(.A(G1698), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n266), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G226), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n317), .B(new_n318), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n257), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n275), .B1(G238), .B2(new_n278), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT13), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT14), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n326), .A2(new_n330), .A3(G169), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n329), .B(new_n331), .C1(new_n282), .C2(new_n326), .ZN(new_n332));
  INV_X1    g0132(.A(new_n292), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n333), .A2(new_n202), .B1(new_n209), .B2(G68), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n300), .A2(new_n219), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n288), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT11), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n289), .A2(G68), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT12), .ZN(new_n341));
  INV_X1    g0141(.A(new_n285), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n213), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n336), .A2(new_n337), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n339), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n332), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n327), .A2(G190), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n326), .A2(G200), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G20), .A2(G77), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT8), .B(G58), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n354), .B1(new_n355), .B2(new_n300), .C1(new_n333), .C2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n357), .A2(new_n288), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n289), .A2(G77), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G77), .B2(new_n285), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n266), .A2(G232), .A3(new_n319), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n362), .B1(new_n221), .B2(new_n266), .C1(new_n268), .C2(new_n214), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n257), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n275), .B1(G244), .B2(new_n278), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n361), .B1(new_n367), .B2(new_n308), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT76), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n369), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(G190), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n372), .A2(KEYINPUT75), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(KEYINPUT75), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n370), .A2(new_n371), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n361), .B1(new_n328), .B2(new_n366), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(G179), .B2(new_n366), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n316), .A2(new_n353), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n299), .A2(new_n289), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n299), .B2(new_n285), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  INV_X1    g0183(.A(G159), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n333), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n201), .B1(new_n297), .B2(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n209), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n266), .B2(G20), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n261), .A2(G33), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT7), .B(new_n209), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n213), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n383), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n288), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT79), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT16), .B(new_n386), .C1(new_n387), .C2(new_n209), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT78), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n263), .A2(new_n400), .A3(KEYINPUT7), .A4(new_n209), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n401), .A3(new_n390), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n398), .B1(new_n402), .B2(G68), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n396), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n288), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n263), .B2(new_n209), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n389), .B(G20), .C1(new_n260), .C2(new_n262), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(KEYINPUT71), .A2(G58), .ZN(new_n409));
  NOR2_X1   g0209(.A1(KEYINPUT71), .A2(G58), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n209), .B1(new_n411), .B2(new_n232), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n385), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n405), .B1(new_n414), .B2(new_n383), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n402), .A2(G68), .ZN(new_n416));
  INV_X1    g0216(.A(new_n398), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT79), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n382), .B1(new_n404), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT80), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n397), .B1(new_n396), .B2(new_n403), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n418), .A2(KEYINPUT79), .A3(new_n288), .A4(new_n395), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n381), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT80), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n320), .A2(new_n267), .B1(new_n259), .B2(new_n215), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n268), .A2(new_n321), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n257), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n275), .B1(G232), .B2(new_n278), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n282), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(G169), .B2(new_n431), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n421), .A2(new_n426), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n308), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(G190), .B2(new_n431), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n424), .A2(KEYINPUT81), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT81), .B1(new_n424), .B2(new_n438), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT17), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT17), .B1(new_n424), .B2(new_n438), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n421), .A2(new_n426), .A3(new_n444), .A4(new_n434), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n436), .A2(new_n441), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n379), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT82), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT6), .ZN(new_n450));
  INV_X1    g0250(.A(G97), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n221), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n452), .B2(new_n205), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n221), .A2(KEYINPUT6), .A3(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n455), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n456));
  OAI21_X1  g0256(.A(G107), .B1(new_n406), .B2(new_n407), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n449), .B1(new_n458), .B2(new_n288), .ZN(new_n459));
  AOI211_X1 g0259(.A(KEYINPUT82), .B(new_n405), .C1(new_n456), .C2(new_n457), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n285), .A2(G97), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT83), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n259), .B2(G1), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n208), .A2(KEYINPUT83), .A3(G33), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n285), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n288), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n462), .B1(new_n467), .B2(G97), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n461), .A2(KEYINPUT84), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n459), .B2(new_n460), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT84), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT4), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n320), .B2(new_n220), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G283), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n473), .A2(new_n475), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n208), .B(G45), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n258), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n478), .A2(new_n257), .B1(G257), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G274), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G200), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n484), .A2(new_n486), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G190), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n469), .A2(new_n472), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(G179), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(G169), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n470), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n266), .A2(new_n209), .A3(G87), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n496), .B(KEYINPUT22), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT23), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n209), .B2(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n221), .A2(KEYINPUT23), .A3(G20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n499), .A2(new_n500), .B1(new_n502), .B2(new_n209), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT24), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n288), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n486), .B1(new_n222), .B2(new_n482), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n266), .A2(G257), .A3(G1698), .ZN(new_n508));
  INV_X1    g0308(.A(G294), .ZN(new_n509));
  OAI221_X1 g0309(.A(new_n508), .B1(new_n259), .B2(new_n509), .C1(new_n320), .C2(new_n216), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n257), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G190), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT25), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n285), .B2(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n342), .A2(KEYINPUT25), .A3(new_n221), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n467), .A2(G107), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g0316(.A1(new_n511), .A2(new_n308), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n506), .A2(new_n512), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n491), .A2(new_n495), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n486), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(G270), .B2(new_n483), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n266), .A2(G257), .A3(new_n319), .ZN(new_n522));
  INV_X1    g0322(.A(G303), .ZN(new_n523));
  OAI221_X1 g0323(.A(new_n522), .B1(new_n523), .B2(new_n266), .C1(new_n268), .C2(new_n222), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n257), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(G179), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n477), .B(new_n209), .C1(G33), .C2(new_n451), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(new_n288), .C1(new_n209), .C2(G116), .ZN(new_n529));
  XOR2_X1   g0329(.A(new_n529), .B(KEYINPUT20), .Z(new_n530));
  NOR2_X1   g0330(.A1(new_n285), .A2(G116), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n467), .B2(G116), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n521), .A2(new_n525), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(new_n533), .A3(KEYINPUT21), .A4(G169), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n533), .A3(G169), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT21), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n533), .B1(G200), .B2(new_n535), .ZN(new_n541));
  INV_X1    g0341(.A(G190), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n535), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n537), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(G250), .B1(new_n276), .B2(G1), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n257), .A2(new_n545), .B1(new_n276), .B2(new_n272), .ZN(new_n546));
  OAI221_X1 g0346(.A(new_n501), .B1(new_n268), .B2(new_n220), .C1(new_n214), .C2(new_n320), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n257), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G179), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n328), .B2(new_n548), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT85), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT85), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n549), .B(new_n552), .C1(new_n328), .C2(new_n548), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n266), .A2(new_n209), .A3(G68), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n209), .B1(new_n318), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G87), .B2(new_n206), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n300), .B2(new_n451), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n288), .B1(new_n342), .B2(new_n355), .ZN(new_n561));
  INV_X1    g0361(.A(new_n467), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n355), .B(KEYINPUT86), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n554), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n548), .A2(new_n308), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n467), .A2(G87), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT87), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n561), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT88), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n548), .A2(G190), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT88), .B1(new_n566), .B2(new_n570), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n511), .A2(G169), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n511), .A2(new_n282), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n506), .B2(new_n516), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n544), .A2(new_n565), .A3(new_n576), .A4(new_n581), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n448), .A2(new_n519), .A3(new_n582), .ZN(G372));
  INV_X1    g0383(.A(new_n352), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n349), .B1(new_n584), .B2(new_n377), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n424), .A2(new_n438), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT81), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n424), .A2(KEYINPUT81), .A3(new_n438), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n442), .B1(new_n590), .B2(KEYINPUT17), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n424), .A2(new_n433), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n593), .B(KEYINPUT18), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n592), .A2(new_n595), .B1(new_n314), .B2(new_n315), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n596), .A2(new_n305), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n571), .A2(new_n574), .B1(new_n550), .B2(new_n564), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n491), .A2(new_n495), .A3(new_n518), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n537), .A2(new_n540), .ZN(new_n600));
  XOR2_X1   g0400(.A(new_n600), .B(KEYINPUT89), .Z(new_n601));
  AOI21_X1  g0401(.A(new_n599), .B1(new_n601), .B2(new_n581), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n492), .A2(new_n493), .B1(new_n461), .B2(new_n468), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n565), .A2(new_n576), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT26), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n550), .A2(new_n564), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n469), .A2(new_n472), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n494), .A3(new_n598), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n605), .B(new_n606), .C1(KEYINPUT26), .C2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n597), .B1(new_n448), .B2(new_n610), .ZN(G369));
  NAND3_X1  g0411(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(G213), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(G343), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n533), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n544), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n601), .B2(new_n618), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G330), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n581), .A2(new_n617), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n506), .A2(new_n516), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n617), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n580), .B1(new_n624), .B2(new_n518), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n617), .B1(new_n537), .B2(new_n540), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n625), .A2(new_n631), .B1(new_n581), .B2(new_n617), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(G399));
  INV_X1    g0434(.A(new_n228), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(G41), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G1), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n233), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT28), .ZN(new_n641));
  INV_X1    g0441(.A(new_n617), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n608), .A2(KEYINPUT26), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n565), .A2(new_n576), .A3(new_n603), .A4(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n645), .A3(new_n606), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n600), .A2(new_n580), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n599), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(KEYINPUT29), .B(new_n642), .C1(new_n646), .C2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n610), .A2(new_n617), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(KEYINPUT29), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n582), .A2(new_n519), .A3(new_n617), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n511), .A2(new_n548), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(new_n527), .A3(KEYINPUT30), .A4(new_n484), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT30), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n484), .A2(new_n511), .A3(new_n548), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n656), .B2(new_n526), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n548), .B1(new_n525), .B2(new_n521), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n511), .A2(G179), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n487), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n654), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n617), .A3(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n661), .A2(new_n617), .ZN(new_n665));
  OAI211_X1 g0465(.A(KEYINPUT91), .B(new_n664), .C1(new_n665), .C2(KEYINPUT31), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT91), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n661), .A2(new_n617), .A3(new_n663), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT31), .B1(new_n661), .B2(new_n617), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(G330), .B1(new_n652), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT92), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(KEYINPUT92), .B(G330), .C1(new_n652), .C2(new_n671), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n651), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n641), .B1(new_n678), .B2(G1), .ZN(G364));
  INV_X1    g0479(.A(G13), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G20), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n208), .B1(new_n681), .B2(G45), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n636), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n235), .B1(G20), .B2(new_n328), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT95), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT95), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(G13), .A2(G33), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT94), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G20), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT96), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n228), .A2(G355), .A3(new_n266), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(G116), .B2(new_n228), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n228), .A2(new_n263), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT93), .Z(new_n699));
  AOI22_X1  g0499(.A1(new_n255), .A2(G45), .B1(new_n234), .B2(new_n273), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n684), .B1(new_n695), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n209), .A2(G179), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n542), .A3(G200), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT97), .Z(new_n705));
  NOR2_X1   g0505(.A1(G190), .A2(G200), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n705), .A2(G283), .B1(G329), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT98), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n209), .A2(new_n282), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G200), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n542), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G326), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n542), .A2(G179), .A3(G200), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n209), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n703), .A2(G190), .A3(G200), .ZN(new_n717));
  OAI221_X1 g0517(.A(new_n714), .B1(new_n509), .B2(new_n716), .C1(new_n523), .C2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n712), .A2(G190), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT33), .B(G317), .Z(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(KEYINPUT99), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(KEYINPUT99), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n711), .A2(new_n706), .ZN(new_n723));
  INV_X1    g0523(.A(G311), .ZN(new_n724));
  INV_X1    g0524(.A(G322), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n711), .A2(G190), .A3(new_n308), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n263), .B1(new_n723), .B2(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  NOR4_X1   g0527(.A1(new_n710), .A2(new_n718), .A3(new_n722), .A4(new_n727), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(KEYINPUT100), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(KEYINPUT100), .ZN(new_n730));
  INV_X1    g0530(.A(new_n719), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n731), .A2(new_n213), .B1(new_n717), .B2(new_n215), .ZN(new_n732));
  INV_X1    g0532(.A(new_n713), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n708), .A2(G159), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n733), .A2(new_n202), .B1(new_n734), .B2(KEYINPUT32), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n705), .A2(G107), .ZN(new_n737));
  INV_X1    g0537(.A(new_n297), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n266), .B1(new_n723), .B2(new_n219), .C1(new_n738), .C2(new_n726), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n716), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n734), .A2(KEYINPUT32), .B1(new_n741), .B2(G97), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n736), .A2(new_n737), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n729), .A2(new_n730), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n702), .B1(new_n744), .B2(new_n688), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n620), .B2(new_n693), .ZN(new_n746));
  INV_X1    g0546(.A(new_n684), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n621), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n620), .A2(G330), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT101), .ZN(G396));
  NOR2_X1   g0551(.A1(new_n377), .A2(new_n617), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n375), .B1(new_n361), .B2(new_n642), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n752), .B1(new_n753), .B2(new_n377), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n650), .B(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n684), .B1(new_n755), .B2(new_n677), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n677), .B2(new_n755), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n688), .A2(new_n690), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n747), .B1(new_n758), .B2(new_n219), .ZN(new_n759));
  INV_X1    g0559(.A(new_n705), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n215), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G97), .A2(new_n741), .B1(new_n719), .B2(G283), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(new_n523), .B2(new_n733), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n263), .B1(new_n717), .B2(new_n221), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT102), .ZN(new_n765));
  INV_X1    g0565(.A(new_n726), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n766), .A2(G294), .B1(new_n708), .B2(G311), .ZN(new_n767));
  INV_X1    g0567(.A(G116), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n768), .B2(new_n723), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n761), .A2(new_n763), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT103), .ZN(new_n772));
  INV_X1    g0572(.A(new_n723), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n766), .A2(G143), .B1(new_n773), .B2(G159), .ZN(new_n774));
  INV_X1    g0574(.A(G137), .ZN(new_n775));
  INV_X1    g0575(.A(G150), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n774), .B1(new_n733), .B2(new_n775), .C1(new_n776), .C2(new_n731), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT34), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n705), .A2(G68), .ZN(new_n781));
  INV_X1    g0581(.A(G132), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n266), .B1(new_n707), .B2(new_n782), .C1(new_n716), .C2(new_n738), .ZN(new_n783));
  INV_X1    g0583(.A(new_n717), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(G50), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n771), .A2(KEYINPUT103), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n772), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n759), .B1(new_n689), .B2(new_n788), .C1(new_n754), .C2(new_n691), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n757), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G384));
  NOR2_X1   g0591(.A1(new_n681), .A2(new_n208), .ZN(new_n792));
  INV_X1    g0592(.A(G330), .ZN(new_n793));
  INV_X1    g0593(.A(new_n615), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n418), .A2(new_n288), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n388), .B1(new_n402), .B2(G68), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT104), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT16), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n794), .B1(new_n800), .B2(new_n381), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n800), .A2(new_n381), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n801), .B1(new_n803), .B2(new_n433), .ZN(new_n804));
  OAI21_X1  g0604(.A(KEYINPUT37), .B1(new_n590), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n421), .B(new_n426), .C1(new_n434), .C2(new_n794), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT37), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n806), .A2(new_n807), .A3(new_n588), .A4(new_n589), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n446), .A2(new_n802), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(KEYINPUT105), .B1(new_n809), .B2(KEYINPUT38), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT38), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n422), .A2(new_n423), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n425), .B1(new_n812), .B2(new_n382), .ZN(new_n813));
  AOI211_X1 g0613(.A(KEYINPUT80), .B(new_n381), .C1(new_n422), .C2(new_n423), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n444), .B1(new_n815), .B2(new_n434), .ZN(new_n816));
  INV_X1    g0616(.A(new_n445), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n801), .B1(new_n818), .B2(new_n591), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n805), .A2(new_n808), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n811), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n810), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(KEYINPUT105), .B(new_n811), .C1(new_n819), .C2(new_n820), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n349), .B(new_n352), .C1(new_n347), .C2(new_n642), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n348), .B(new_n617), .C1(new_n332), .C2(new_n584), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n754), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n665), .A2(KEYINPUT31), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n663), .B2(new_n665), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n652), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n822), .A2(new_n823), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT40), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT106), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n832), .A2(KEYINPUT106), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n809), .A2(KEYINPUT38), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n421), .A2(new_n426), .A3(new_n794), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n591), .B2(new_n594), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n590), .A2(KEYINPUT37), .ZN(new_n841));
  INV_X1    g0641(.A(new_n593), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n839), .A2(new_n586), .A3(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n841), .A2(new_n806), .B1(new_n843), .B2(KEYINPUT37), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n811), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT107), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n838), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n838), .B2(new_n845), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n831), .A2(KEYINPUT40), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n836), .A2(new_n837), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT108), .Z(new_n853));
  NOR2_X1   g0653(.A1(new_n448), .A2(new_n830), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n793), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n853), .B2(new_n854), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n595), .A2(new_n615), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n642), .B(new_n754), .C1(new_n602), .C2(new_n609), .ZN(new_n858));
  INV_X1    g0658(.A(new_n752), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n826), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n822), .A2(new_n823), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n857), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n838), .A2(new_n845), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT39), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(KEYINPUT39), .B2(new_n862), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n332), .A2(new_n348), .A3(new_n642), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n863), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n597), .B1(new_n651), .B2(new_n448), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n871), .B(new_n872), .Z(new_n873));
  AOI21_X1  g0673(.A(new_n792), .B1(new_n856), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n873), .B2(new_n856), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(G116), .A3(new_n236), .A4(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT36), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n234), .A2(G77), .A3(new_n411), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(G50), .B2(new_n213), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G1), .A3(new_n680), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n875), .A2(new_n879), .A3(new_n882), .ZN(G367));
  NAND2_X1  g0683(.A1(new_n607), .A2(new_n617), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n495), .A3(new_n491), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n607), .A2(new_n494), .A3(new_n617), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n629), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n580), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n617), .B1(new_n891), .B2(new_n495), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n626), .A2(new_n887), .A3(new_n630), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT109), .Z(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n894), .B2(KEYINPUT42), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(KEYINPUT42), .B2(new_n894), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n570), .A2(new_n617), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n598), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n606), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT43), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n899), .A2(KEYINPUT43), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n896), .A2(KEYINPUT43), .A3(new_n899), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n890), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OR3_X1    g0705(.A1(new_n903), .A2(new_n890), .A3(new_n904), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n636), .B(KEYINPUT41), .Z(new_n907));
  NOR2_X1   g0707(.A1(new_n633), .A2(new_n887), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT44), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT110), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n633), .A2(new_n910), .A3(new_n887), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT110), .B1(new_n888), .B2(new_n632), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT45), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT45), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(new_n628), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n626), .B(new_n631), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n621), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n678), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n907), .B1(new_n922), .B2(new_n678), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n905), .B(new_n906), .C1(new_n923), .C2(new_n683), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n228), .A2(new_n355), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n695), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n699), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(new_n243), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n747), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AOI22_X1  g0729(.A1(G50), .A2(new_n773), .B1(new_n708), .B2(G137), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n266), .C1(new_n776), .C2(new_n726), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n713), .A2(G143), .B1(new_n784), .B2(new_n297), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n219), .B2(new_n704), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n731), .A2(new_n384), .B1(new_n213), .B2(new_n716), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT111), .Z(new_n936));
  OAI22_X1  g0736(.A1(new_n731), .A2(new_n509), .B1(new_n451), .B2(new_n704), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n733), .A2(new_n724), .B1(new_n221), .B2(new_n716), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G317), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n263), .B1(new_n707), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(G283), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n726), .A2(new_n523), .B1(new_n723), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT46), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n784), .A2(G116), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n941), .B(new_n943), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n939), .B(new_n946), .C1(new_n944), .C2(new_n945), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n936), .A2(KEYINPUT47), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n688), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT47), .B1(new_n936), .B2(new_n947), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n929), .B1(new_n949), .B2(new_n950), .C1(new_n693), .C2(new_n899), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n924), .A2(new_n951), .ZN(G387));
  AOI22_X1  g0752(.A1(new_n766), .A2(G317), .B1(new_n773), .B2(G303), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n733), .B2(new_n725), .C1(new_n724), .C2(new_n731), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT48), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n741), .A2(G283), .B1(new_n784), .B2(G294), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n960), .A2(KEYINPUT49), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(KEYINPUT49), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n704), .A2(new_n768), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n266), .B(new_n963), .C1(G326), .C2(new_n708), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n299), .A2(new_n731), .B1(new_n213), .B2(new_n723), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT113), .Z(new_n967));
  OR2_X1    g0767(.A1(new_n563), .A2(new_n716), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n266), .B1(new_n726), .B2(new_n202), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G150), .B2(new_n708), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n717), .A2(new_n219), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G159), .B2(new_n713), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n968), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n967), .B(new_n973), .C1(new_n451), .C2(new_n760), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n689), .B1(new_n965), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n247), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n699), .B1(new_n976), .B2(new_n273), .ZN(new_n977));
  INV_X1    g0777(.A(new_n638), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n228), .A3(new_n266), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n356), .A2(KEYINPUT50), .A3(G50), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT50), .B1(new_n356), .B2(G50), .ZN(new_n982));
  AOI21_X1  g0782(.A(G45), .B1(G68), .B2(G77), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n981), .A2(new_n638), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n980), .A2(new_n984), .B1(new_n221), .B2(new_n635), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n684), .B1(new_n985), .B2(new_n695), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT112), .Z(new_n987));
  AOI211_X1 g0787(.A(new_n975), .B(new_n987), .C1(new_n627), .C2(new_n692), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT114), .Z(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n920), .B2(new_n683), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n921), .A2(new_n636), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n678), .A2(new_n920), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(G393));
  NAND2_X1  g0793(.A1(new_n918), .A2(new_n921), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n922), .A2(new_n636), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT115), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n682), .B1(new_n918), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n996), .B2(new_n918), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n927), .A2(new_n251), .B1(new_n451), .B2(new_n228), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n684), .B1(new_n999), .B2(new_n695), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n263), .B1(new_n707), .B2(new_n725), .C1(new_n942), .C2(new_n717), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n705), .B2(G107), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT117), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n741), .A2(G116), .B1(new_n773), .B2(G294), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n523), .B2(new_n731), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n733), .A2(new_n940), .B1(new_n724), .B2(new_n726), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n716), .A2(new_n219), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G68), .B2(new_n784), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n202), .B2(new_n731), .ZN(new_n1012));
  INV_X1    g0812(.A(G143), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n266), .B1(new_n707), .B2(new_n1013), .C1(new_n356), .C2(new_n723), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n761), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G150), .A2(new_n713), .B1(new_n766), .B2(G159), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT51), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n1003), .A2(new_n1009), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1000), .B1(new_n1018), .B2(new_n688), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n887), .B2(new_n693), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n995), .A2(new_n998), .A3(new_n1020), .ZN(G390));
  NAND2_X1  g0821(.A1(new_n753), .A2(new_n377), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n642), .B(new_n1022), .C1(new_n646), .C2(new_n648), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n859), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(KEYINPUT118), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT118), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1026), .A3(new_n859), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n826), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n849), .A2(new_n869), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n676), .A2(new_n754), .A3(new_n826), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n861), .A2(new_n869), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1029), .B(new_n1030), .C1(new_n868), .C2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n864), .A2(KEYINPUT107), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n838), .A2(new_n845), .A3(new_n846), .ZN(new_n1035));
  AND4_X1   g0835(.A1(new_n869), .A2(new_n1028), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n862), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n866), .B1(new_n1037), .B2(new_n865), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1036), .B1(new_n1038), .B2(new_n1031), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n830), .A2(new_n793), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n827), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1033), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n826), .B1(new_n676), .B2(new_n754), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1042), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n860), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1040), .A2(new_n754), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n826), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1030), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n379), .A2(new_n447), .A3(new_n1040), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n597), .B(new_n1053), .C1(new_n651), .C2(new_n448), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n637), .B1(new_n1043), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1033), .B(new_n1058), .C1(new_n1039), .C2(new_n1042), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT54), .B(G143), .ZN(new_n1061));
  INV_X1    g0861(.A(G125), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n723), .A2(new_n1061), .B1(new_n707), .B2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n263), .B(new_n1063), .C1(G132), .C2(new_n766), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n717), .A2(new_n776), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT53), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G159), .A2(new_n741), .B1(new_n719), .B2(G137), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n704), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n713), .A2(G128), .B1(new_n1068), .B2(G50), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n263), .B1(new_n717), .B2(new_n215), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT119), .Z(new_n1072));
  OAI22_X1  g0872(.A1(new_n726), .A2(new_n768), .B1(new_n723), .B2(new_n451), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G294), .B2(new_n708), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n719), .A2(G107), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1010), .B1(G283), .B2(new_n713), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n781), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1070), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n688), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n747), .B1(new_n758), .B2(new_n299), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n868), .C2(new_n691), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1043), .B2(new_n682), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1060), .A2(new_n1082), .ZN(G378));
  INV_X1    g0883(.A(KEYINPUT123), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n871), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n303), .A2(new_n794), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT55), .Z(new_n1087));
  AND2_X1   g0887(.A1(new_n316), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n316), .A2(new_n1087), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OR3_X1    g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n836), .A2(new_n837), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n793), .B1(new_n849), .B2(new_n851), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n832), .A2(KEYINPUT106), .A3(new_n833), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT106), .B1(new_n832), .B2(new_n833), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1096), .B(new_n1094), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1085), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1094), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n871), .A3(new_n1100), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n682), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1094), .A2(new_n691), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n747), .B1(new_n758), .B2(new_n202), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT121), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n266), .A2(G41), .ZN(new_n1111));
  AOI211_X1 g0911(.A(G50), .B(new_n1111), .C1(new_n259), .C2(new_n274), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1111), .B1(new_n942), .B2(new_n707), .C1(new_n221), .C2(new_n726), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n971), .B(new_n1113), .C1(G68), .C2(new_n741), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n713), .A2(G116), .B1(new_n1068), .B2(new_n297), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n451), .B2(new_n731), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1114), .B(new_n1117), .C1(new_n563), .C2(new_n723), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT58), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1112), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT120), .B(G124), .ZN(new_n1121));
  AOI211_X1 g0921(.A(G33), .B(G41), .C1(new_n708), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(G128), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n726), .A2(new_n1123), .B1(new_n723), .B2(new_n775), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1061), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n719), .A2(G132), .B1(new_n784), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1062), .B2(new_n733), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1124), .B(new_n1127), .C1(G150), .C2(new_n741), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT59), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1122), .B1(new_n384), .B2(new_n704), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1128), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1120), .B1(new_n1119), .B2(new_n1118), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1110), .B1(new_n1133), .B2(new_n688), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1108), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1084), .B1(new_n1107), .B2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1105), .A2(new_n871), .A3(new_n1100), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n871), .B1(new_n1105), .B2(new_n1100), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n683), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(KEYINPUT123), .A3(new_n1135), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1059), .A2(new_n1055), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1143), .B(KEYINPUT57), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n636), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1142), .A2(new_n1148), .ZN(G375));
  NAND2_X1  g0949(.A1(new_n1049), .A2(new_n690), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT124), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n688), .A2(G68), .A3(new_n690), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n731), .A2(new_n768), .B1(new_n733), .B2(new_n509), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G97), .B2(new_n784), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n705), .A2(G77), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n726), .A2(new_n942), .B1(new_n707), .B2(new_n523), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n266), .B(new_n1156), .C1(G107), .C2(new_n773), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n968), .A3(new_n1155), .A4(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n719), .A2(new_n1125), .B1(new_n784), .B2(G159), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n202), .B2(new_n716), .C1(new_n738), .C2(new_n704), .ZN(new_n1160));
  OR3_X1    g0960(.A1(new_n733), .A2(KEYINPUT125), .A3(new_n782), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n766), .A2(G137), .B1(new_n773), .B2(G150), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT125), .B1(new_n733), .B2(new_n782), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n263), .B1(new_n708), .B2(G128), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1158), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n747), .B(new_n1152), .C1(new_n1166), .C2(new_n688), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1052), .A2(new_n683), .B1(new_n1151), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1052), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1054), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1058), .A2(new_n907), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1168), .B1(new_n1171), .B2(new_n1172), .ZN(G381));
  NOR2_X1   g0973(.A1(new_n1060), .A2(new_n1082), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1142), .A2(new_n1148), .A3(new_n1174), .ZN(new_n1175));
  OR4_X1    g0975(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1176));
  OR4_X1    g0976(.A1(G387), .A2(new_n1175), .A3(G381), .A4(new_n1176), .ZN(G407));
  NAND2_X1  g0977(.A1(new_n616), .A2(G213), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT126), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(G407), .B(G213), .C1(new_n1175), .C2(new_n1180), .ZN(G409));
  NAND3_X1  g0981(.A1(new_n1142), .A2(new_n1148), .A3(G378), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1140), .B(new_n1135), .C1(new_n1144), .C2(new_n907), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1174), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT60), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1170), .B1(new_n1186), .B2(new_n1058), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1169), .A2(KEYINPUT60), .A3(new_n1054), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n636), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1168), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n790), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(G384), .A3(new_n1168), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1185), .A2(new_n1178), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT63), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1185), .A2(new_n1178), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n616), .A2(G213), .A3(G2897), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1191), .A2(new_n1192), .A3(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1191), .A2(new_n1192), .B1(G2897), .B2(new_n1179), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1197), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1179), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(KEYINPUT63), .A3(new_n1193), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(G387), .A2(new_n995), .A3(new_n1020), .A4(new_n998), .ZN(new_n1206));
  XOR2_X1   g1006(.A(G393), .B(G396), .Z(new_n1207));
  NAND3_X1  g1007(.A1(new_n924), .A2(new_n951), .A3(G390), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1209), .A2(new_n1210), .A3(KEYINPUT61), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1196), .A2(new_n1203), .A3(new_n1205), .A4(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT61), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1204), .B2(new_n1201), .ZN(new_n1214));
  XOR2_X1   g1014(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1215));
  NAND2_X1  g1015(.A1(new_n1194), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1204), .A2(KEYINPUT62), .A3(new_n1193), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1212), .B1(new_n1218), .B2(new_n1219), .ZN(G405));
  NAND2_X1  g1020(.A1(G375), .A2(new_n1174), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1182), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1193), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1222), .A2(new_n1193), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1224), .A2(new_n1225), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1225), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n1223), .A3(new_n1219), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(G402));
endmodule


