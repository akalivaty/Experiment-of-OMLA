//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G68), .A2(G238), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G50), .A2(G226), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G116), .A2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n214), .B(new_n220), .C1(G97), .C2(G257), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G1), .B2(G20), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  INV_X1    g0023(.A(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n206), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n207), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n210), .B(new_n223), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT72), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n247));
  INV_X1    g0047(.A(G274), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n225), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AND3_X1   g0052(.A1(new_n252), .A2(G226), .A3(new_n247), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G222), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT64), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G77), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT64), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n254), .A2(new_n264), .A3(G222), .A4(new_n255), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n254), .A2(G223), .A3(G1698), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n258), .A2(new_n263), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n252), .ZN(new_n268));
  AOI211_X1 g0068(.A(new_n249), .B(new_n253), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n246), .B1(new_n269), .B2(G190), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n268), .ZN(new_n271));
  INV_X1    g0071(.A(new_n249), .ZN(new_n272));
  INV_X1    g0072(.A(new_n253), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G200), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n226), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n206), .A2(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G50), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n224), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G58), .A2(G68), .ZN(new_n286));
  INV_X1    g0086(.A(G50), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n207), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(KEYINPUT8), .A2(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT8), .A2(G58), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT66), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT66), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(new_n297), .A3(new_n294), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n207), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI211_X1 g0101(.A(new_n288), .B(new_n292), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n281), .B(new_n285), .C1(new_n302), .C2(new_n279), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n303), .A2(KEYINPUT9), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(KEYINPUT9), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n270), .B(new_n275), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT12), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n283), .B2(G68), .ZN(new_n309));
  INV_X1    g0109(.A(G68), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n282), .A2(KEYINPUT12), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n279), .A2(new_n280), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n309), .B(new_n311), .C1(new_n312), .C2(new_n310), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n290), .A2(new_n287), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n300), .A2(new_n216), .B1(new_n207), .B2(G68), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n278), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g0119(.A(new_n319), .B(KEYINPUT11), .Z(new_n320));
  NOR2_X1   g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  INV_X1    g0122(.A(G232), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G1698), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(G226), .B2(G1698), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n322), .B1(new_n325), .B2(new_n262), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n249), .B1(new_n326), .B2(new_n268), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n252), .A2(new_n247), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G238), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n327), .B2(new_n329), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G190), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n321), .B(new_n335), .C1(new_n334), .C2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT67), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n274), .A2(new_n338), .A3(G179), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT67), .B1(new_n269), .B2(new_n340), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n303), .B1(G169), .B2(new_n269), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n307), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT70), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n254), .A2(G238), .A3(G1698), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n345), .B1(new_n203), .B2(new_n254), .C1(new_n256), .C2(new_n323), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n268), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n328), .A2(G244), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n272), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT68), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n347), .A2(KEYINPUT68), .A3(new_n272), .A4(new_n348), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G200), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT15), .B(G87), .Z(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n301), .B1(G20), .B2(G77), .ZN(new_n356));
  INV_X1    g0156(.A(new_n295), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n289), .A2(KEYINPUT69), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n289), .A2(KEYINPUT69), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n279), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n312), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(G77), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n282), .A2(new_n216), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n344), .B1(new_n354), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n351), .A2(new_n352), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G190), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n353), .A2(KEYINPUT70), .A3(new_n364), .A4(new_n363), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n367), .A2(new_n340), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n351), .A2(new_n372), .A3(new_n352), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n373), .A3(new_n365), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT71), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n370), .A2(KEYINPUT71), .A3(new_n374), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n343), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n260), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n250), .A2(KEYINPUT75), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G33), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n380), .B1(new_n384), .B2(KEYINPUT3), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT7), .B1(new_n385), .B2(G20), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT76), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT75), .B(G33), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n260), .B1(new_n389), .B2(new_n259), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n207), .ZN(new_n394));
  OAI211_X1 g0194(.A(G68), .B(new_n386), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n381), .A2(new_n383), .A3(new_n259), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n399), .B2(new_n261), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n400), .A2(new_n393), .B1(new_n254), .B2(new_n394), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n397), .B1(new_n401), .B2(new_n310), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n398), .A2(new_n404), .A3(new_n278), .ZN(new_n405));
  INV_X1    g0205(.A(new_n299), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n283), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n362), .B2(new_n406), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n250), .A2(new_n218), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n385), .B1(G223), .B2(G1698), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n255), .A2(G226), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n249), .B1(new_n414), .B2(new_n268), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n328), .A2(G232), .ZN(new_n416));
  AOI21_X1  g0216(.A(G169), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G223), .A2(G1698), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n390), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n268), .B1(new_n419), .B2(new_n410), .ZN(new_n420));
  AND4_X1   g0220(.A1(new_n340), .A2(new_n420), .A3(new_n416), .A4(new_n272), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n417), .A2(KEYINPUT77), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT77), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n415), .A2(new_n340), .A3(new_n416), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(new_n416), .A3(new_n272), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n372), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n423), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n409), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT77), .B1(new_n417), .B2(new_n421), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n424), .A2(new_n423), .A3(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(KEYINPUT18), .A3(new_n409), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n415), .A2(G190), .A3(new_n416), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n425), .A2(G200), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n405), .A2(new_n408), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n438), .A2(new_n439), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT78), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n438), .A2(new_n439), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT78), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n438), .A2(new_n439), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n435), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n334), .A2(KEYINPUT74), .A3(new_n372), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT14), .ZN(new_n451));
  INV_X1    g0251(.A(new_n334), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(new_n340), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n450), .B1(new_n453), .B2(new_n449), .C1(new_n316), .C2(new_n320), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n379), .A2(new_n448), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n379), .A2(KEYINPUT79), .A3(new_n448), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n207), .A2(G87), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n260), .C1(new_n389), .C2(new_n259), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n262), .B2(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT87), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT82), .B(G116), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n384), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n207), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n207), .A2(G107), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT23), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT24), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(KEYINPUT88), .A3(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n466), .A2(new_n468), .B1(new_n207), .B2(new_n471), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n476), .A2(KEYINPUT88), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(KEYINPUT88), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n478), .A2(new_n474), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n477), .A2(new_n278), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n250), .A2(G1), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n278), .A2(new_n282), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G107), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n282), .A2(new_n203), .ZN(new_n486));
  XOR2_X1   g0286(.A(new_n486), .B(KEYINPUT25), .Z(new_n487));
  NAND3_X1  g0287(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n219), .A2(G1698), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n260), .B(new_n489), .C1(new_n389), .C2(new_n259), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT89), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n389), .A2(G294), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n382), .A2(G33), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n250), .A2(KEYINPUT75), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT3), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT89), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(new_n260), .A4(new_n489), .ZN(new_n497));
  AND2_X1   g0297(.A1(G257), .A2(G1698), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n260), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n491), .A2(new_n492), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n268), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT90), .ZN(new_n502));
  XNOR2_X1  g0302(.A(KEYINPUT5), .B(G41), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n206), .A3(G45), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n504), .A2(new_n252), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G264), .ZN(new_n506));
  INV_X1    g0306(.A(G45), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n507), .A2(new_n248), .A3(G1), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT90), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n500), .A2(new_n511), .A3(new_n268), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n502), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT91), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n502), .A2(KEYINPUT91), .A3(new_n510), .A4(new_n512), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n372), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n510), .A2(new_n501), .A3(G179), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n488), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT92), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(KEYINPUT92), .B(new_n488), .C1(new_n517), .C2(new_n519), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G190), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n515), .A2(new_n525), .A3(new_n516), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n510), .A2(new_n501), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n336), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n484), .A2(new_n355), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT84), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n310), .A2(G20), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n260), .B(new_n535), .C1(new_n389), .C2(new_n259), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n207), .B1(new_n322), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n218), .A2(new_n202), .A3(new_n203), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n537), .B1(new_n300), .B2(new_n202), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT83), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT83), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n543), .B(new_n537), .C1(new_n300), .C2(new_n202), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n536), .A2(new_n540), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n278), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n283), .A2(new_n355), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n534), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI211_X1 g0349(.A(KEYINPUT84), .B(new_n547), .C1(new_n545), .C2(new_n278), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n533), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT85), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(KEYINPUT85), .B(new_n533), .C1(new_n549), .C2(new_n550), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n508), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n252), .B(G250), .C1(G1), .C2(new_n507), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G238), .A2(G1698), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n217), .B2(G1698), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n471), .B1(new_n385), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n556), .B(new_n557), .C1(new_n560), .C2(new_n252), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G169), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n340), .B2(new_n561), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n283), .A2(G97), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT80), .ZN(new_n567));
  XNOR2_X1  g0367(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT6), .B1(new_n204), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G20), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n289), .A2(G77), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n401), .C2(new_n203), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n565), .B1(new_n573), .B2(new_n278), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n484), .A2(G97), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G283), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n254), .B2(G250), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n577), .B(new_n578), .C1(new_n580), .C2(new_n255), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT4), .B1(new_n385), .B2(G244), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n268), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n504), .A2(G257), .A3(new_n252), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n509), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n372), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(new_n260), .C1(new_n389), .C2(new_n259), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n579), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n260), .A2(new_n261), .A3(G250), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT4), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n589), .A2(new_n577), .A3(new_n578), .A4(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n584), .B1(new_n593), .B2(new_n268), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n340), .A3(new_n509), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n576), .A2(new_n587), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n586), .A2(G200), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(G190), .A3(new_n509), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(new_n574), .A4(new_n575), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT81), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n547), .B1(new_n545), .B2(new_n278), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n602), .B(new_n534), .ZN(new_n603));
  INV_X1    g0403(.A(new_n471), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n495), .A2(new_n260), .A3(new_n559), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n252), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n557), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n606), .A2(new_n607), .A3(new_n508), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G190), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n484), .A2(G87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n561), .A2(G200), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n603), .A2(new_n609), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n564), .A2(new_n601), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n470), .A2(G20), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n578), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n278), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT20), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n278), .A2(KEYINPUT20), .A3(new_n615), .A4(new_n616), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n619), .A2(new_n620), .B1(new_n282), .B2(new_n470), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n484), .A2(G116), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n504), .A2(G270), .A3(new_n252), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT86), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n255), .A2(G264), .ZN(new_n628));
  NOR2_X1   g0428(.A1(G257), .A2(G1698), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n390), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(G303), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n254), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n268), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n627), .A2(new_n509), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n624), .B(new_n635), .C1(new_n525), .C2(new_n634), .ZN(new_n636));
  INV_X1    g0436(.A(new_n634), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n623), .A2(new_n637), .A3(G179), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n372), .B1(new_n621), .B2(new_n622), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n639), .A2(new_n640), .A3(new_n634), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n639), .B2(new_n634), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n636), .B(new_n638), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n600), .B1(new_n596), .B2(new_n599), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n614), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n459), .A2(new_n532), .A3(new_n645), .ZN(G372));
  NAND2_X1  g0446(.A1(new_n442), .A2(new_n446), .ZN(new_n647));
  INV_X1    g0447(.A(new_n374), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n337), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n454), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n435), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n307), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n342), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n459), .ZN(new_n655));
  INV_X1    g0455(.A(new_n596), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n564), .A2(new_n613), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT93), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n563), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n562), .B(KEYINPUT93), .C1(new_n340), .C2(new_n561), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n657), .A2(KEYINPUT26), .B1(new_n555), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n555), .A2(new_n661), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n613), .A3(new_n664), .A4(new_n656), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n596), .A2(new_n599), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n612), .B1(new_n555), .B2(new_n661), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n531), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n500), .A2(new_n511), .A3(new_n268), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n511), .B1(new_n500), .B2(new_n268), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT91), .B1(new_n672), .B2(new_n510), .ZN(new_n673));
  INV_X1    g0473(.A(new_n516), .ZN(new_n674));
  OAI21_X1  g0474(.A(G169), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n518), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n669), .B1(new_n676), .B2(new_n488), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n662), .B(new_n665), .C1(new_n668), .C2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n654), .B1(new_n655), .B2(new_n679), .ZN(G369));
  NOR2_X1   g0480(.A1(new_n224), .A2(G20), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n206), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT94), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n532), .B1(new_n530), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n676), .A2(new_n488), .A3(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n669), .A2(new_n623), .A3(new_n689), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n690), .A2(new_n624), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n643), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n669), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n689), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n532), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n676), .A2(new_n488), .A3(new_n690), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n700), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n208), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n539), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n228), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n678), .A2(new_n690), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT98), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n524), .B2(new_n701), .ZN(new_n717));
  AOI211_X1 g0517(.A(KEYINPUT98), .B(new_n669), .C1(new_n522), .C2(new_n523), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n717), .A2(new_n718), .A3(new_n668), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n663), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n664), .B1(new_n667), .B2(new_n656), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n690), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n715), .B1(new_n724), .B2(KEYINPUT29), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n524), .A2(new_n645), .A3(new_n531), .A4(new_n690), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT95), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n594), .A2(new_n509), .A3(new_n633), .A4(new_n627), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n608), .A2(new_n501), .A3(G179), .A4(new_n506), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n727), .B(new_n732), .C1(new_n728), .C2(new_n729), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n527), .A2(new_n586), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT96), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(new_n634), .A3(new_n561), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n340), .B1(new_n734), .B2(new_n735), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n731), .B(new_n733), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT97), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT31), .B1(new_n739), .B2(new_n689), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n739), .A2(new_n689), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n745), .A2(KEYINPUT97), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n726), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G330), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n725), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n713), .B1(new_n751), .B2(G1), .ZN(G364));
  NAND2_X1  g0552(.A1(new_n681), .A2(G45), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n709), .A2(G1), .A3(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n698), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n697), .A2(G330), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(G355), .A2(new_n254), .A3(new_n208), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n392), .A2(new_n707), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G45), .B2(new_n228), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n241), .A2(new_n507), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n758), .B1(G116), .B2(new_n208), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n226), .B1(G20), .B2(new_n372), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n766), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n697), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n207), .A2(new_n340), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n771), .A2(new_n525), .A3(new_n336), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G322), .A2(new_n773), .B1(new_n775), .B2(G311), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n771), .A2(new_n525), .A3(G200), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT33), .B(G317), .Z(new_n778));
  OAI21_X1  g0578(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n772), .A2(new_n336), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n779), .B1(G326), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n336), .A2(G179), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(G20), .A3(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G303), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n525), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT100), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(G179), .A3(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G329), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G179), .A2(G200), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n207), .B1(new_n790), .B2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n262), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n787), .A2(G179), .A3(new_n336), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(new_n794), .B2(G283), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n781), .A2(new_n785), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n773), .ZN(new_n797));
  INV_X1    g0597(.A(G58), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n798), .B1(new_n310), .B2(new_n777), .ZN(new_n799));
  INV_X1    g0599(.A(new_n794), .ZN(new_n800));
  INV_X1    g0600(.A(new_n780), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n203), .B1(new_n287), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n791), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n799), .B(new_n802), .C1(G97), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n784), .A2(G87), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n788), .A2(G159), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT32), .Z(new_n807));
  OR2_X1    g0607(.A1(new_n775), .A2(KEYINPUT99), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n775), .A2(KEYINPUT99), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G77), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n804), .A2(new_n805), .A3(new_n807), .A4(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n796), .B1(new_n813), .B2(new_n262), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n770), .B1(new_n763), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n757), .B1(new_n815), .B2(new_n754), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n816), .B(new_n817), .ZN(G396));
  NOR2_X1   g0618(.A1(new_n374), .A2(new_n689), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n689), .A2(new_n365), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT104), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n370), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n819), .B1(new_n823), .B2(new_n374), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n668), .A2(new_n677), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n564), .A2(new_n656), .A3(new_n613), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n663), .B(new_n665), .C1(new_n826), .C2(new_n664), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n690), .B(new_n824), .C1(new_n825), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT105), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n678), .A2(KEYINPUT105), .A3(new_n690), .A4(new_n824), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n714), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n824), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(new_n749), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n749), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n836), .A3(new_n754), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n800), .A2(new_n218), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G97), .B2(new_n803), .ZN(new_n839));
  INV_X1    g0639(.A(G283), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n801), .A2(new_n631), .B1(new_n840), .B2(new_n777), .ZN(new_n841));
  INV_X1    g0641(.A(new_n470), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n811), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n773), .A2(G294), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n262), .B1(new_n783), .B2(new_n203), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n788), .B2(G311), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n839), .A2(new_n843), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n794), .A2(G68), .B1(G50), .B2(new_n784), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G137), .A2(new_n780), .B1(new_n773), .B2(G143), .ZN(new_n849));
  INV_X1    g0649(.A(G159), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n291), .B2(new_n777), .C1(new_n810), .C2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G58), .B2(new_n803), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n852), .ZN(new_n855));
  INV_X1    g0655(.A(new_n788), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n392), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT103), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n854), .A2(new_n855), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n847), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n763), .A2(new_n764), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n863), .A2(new_n763), .B1(new_n216), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n754), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(new_n824), .C2(new_n765), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n837), .A2(new_n867), .ZN(G384));
  NAND2_X1  g0668(.A1(new_n398), .A2(new_n278), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT16), .B1(new_n395), .B2(new_n397), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n408), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n686), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT106), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n871), .A2(KEYINPUT106), .A3(new_n686), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n447), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n433), .A2(new_n871), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n438), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n409), .A2(new_n686), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n428), .A2(new_n881), .A3(new_n438), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT109), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n428), .A2(new_n438), .A3(new_n882), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(new_n881), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n440), .A2(new_n441), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n882), .B1(new_n435), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n887), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n885), .A2(new_n886), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n886), .B1(new_n885), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n740), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n742), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT108), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n726), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n726), .B2(new_n897), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n337), .B1(new_n321), .B2(new_n690), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n454), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n454), .A2(new_n689), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n824), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n895), .A2(KEYINPUT40), .A3(new_n901), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(KEYINPUT107), .A2(KEYINPUT40), .ZN(new_n909));
  OR2_X1    g0709(.A1(KEYINPUT107), .A2(KEYINPUT40), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n877), .A2(new_n884), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n887), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n885), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n907), .B1(new_n899), .B2(new_n900), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n909), .B(new_n910), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n908), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n901), .A2(new_n459), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n917), .B(new_n918), .Z(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G330), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n885), .A2(new_n892), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n904), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n651), .A2(new_n687), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n819), .B1(new_n830), .B2(new_n831), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n905), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n913), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n928), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n715), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT92), .B1(new_n676), .B2(new_n488), .ZN(new_n936));
  INV_X1    g0736(.A(new_n523), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n701), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT98), .ZN(new_n939));
  INV_X1    g0739(.A(new_n668), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n524), .A2(new_n716), .A3(new_n701), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n689), .B1(new_n942), .B2(new_n722), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT29), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n935), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n653), .B1(new_n945), .B2(new_n459), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n934), .B(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n920), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n206), .B2(new_n681), .ZN(new_n949));
  INV_X1    g0749(.A(G116), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n568), .A2(new_n570), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(KEYINPUT35), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n952), .B(new_n227), .C1(KEYINPUT35), .C2(new_n951), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT36), .ZN(new_n954));
  OAI21_X1  g0754(.A(G77), .B1(new_n798), .B2(new_n310), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n955), .A2(new_n228), .B1(G50), .B2(new_n310), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n224), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n954), .A3(new_n957), .ZN(G367));
  INV_X1    g0758(.A(new_n777), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G150), .A2(new_n773), .B1(new_n959), .B2(G159), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n810), .B2(new_n287), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G77), .A2(new_n794), .B1(new_n788), .B2(G137), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n791), .A2(new_n310), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n262), .B1(new_n784), .B2(G58), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n961), .B(new_n966), .C1(G143), .C2(new_n780), .ZN(new_n967));
  INV_X1    g0767(.A(new_n392), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n773), .A2(G303), .B1(G107), .B2(new_n803), .ZN(new_n969));
  XNOR2_X1  g0769(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n783), .B2(new_n470), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g0772(.A1(KEYINPUT46), .A2(G116), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n788), .A2(G317), .B1(new_n784), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n780), .A2(G311), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n202), .C2(new_n800), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n972), .B(new_n976), .C1(G283), .C2(new_n811), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n959), .A2(G294), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n967), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n754), .B1(new_n980), .B2(new_n763), .ZN(new_n981));
  INV_X1    g0781(.A(new_n355), .ZN(new_n982));
  INV_X1    g0782(.A(new_n759), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n767), .B1(new_n208), .B2(new_n982), .C1(new_n983), .C2(new_n237), .ZN(new_n984));
  INV_X1    g0784(.A(new_n667), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n690), .B1(new_n603), .B2(new_n610), .ZN(new_n986));
  MUX2_X1   g0786(.A(new_n985), .B(new_n663), .S(new_n986), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n766), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n981), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n753), .A2(G1), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n689), .A2(new_n576), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n666), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n596), .B2(new_n690), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n705), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n705), .A2(new_n993), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n699), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n995), .A2(new_n700), .A3(new_n998), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n703), .B1(new_n693), .B2(new_n702), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(new_n698), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n751), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n708), .B(KEYINPUT41), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n990), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n987), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT43), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n703), .A2(new_n992), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT42), .Z(new_n1012));
  OR2_X1    g0812(.A1(new_n524), .A2(new_n992), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n689), .B1(new_n1013), .B2(new_n596), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1009), .B1(new_n1010), .B2(new_n987), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1015), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n699), .A2(new_n993), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n989), .B1(new_n1007), .B2(new_n1019), .ZN(G387));
  AOI21_X1  g0820(.A(new_n709), .B1(new_n1004), .B2(new_n750), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1004), .A2(new_n750), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n773), .A2(G317), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G322), .A2(new_n780), .B1(new_n959), .B2(G311), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n810), .C2(new_n631), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n784), .A2(G294), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n803), .A2(G283), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n788), .A2(G326), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n392), .B1(new_n842), .B2(new_n794), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n856), .A2(new_n291), .B1(new_n406), .B2(new_n777), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G77), .B2(new_n784), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n803), .A2(new_n355), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n794), .A2(G97), .B1(G68), .B2(new_n775), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n797), .A2(new_n287), .B1(new_n801), .B2(new_n850), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n968), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n759), .B1(new_n234), .B2(new_n507), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n710), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n208), .A3(new_n254), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n310), .A2(new_n216), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n357), .A2(new_n287), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1048), .B1(new_n1052), .B2(KEYINPUT50), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n507), .C1(KEYINPUT50), .C2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1050), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(G107), .B2(new_n208), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1046), .A2(new_n763), .B1(new_n767), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n866), .B(new_n1057), .C1(new_n693), .C2(new_n769), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n990), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1023), .B(new_n1058), .C1(new_n1059), .C2(new_n1004), .ZN(G393));
  OR2_X1    g0860(.A1(new_n993), .A2(new_n769), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n767), .B1(new_n202), .B2(new_n208), .C1(new_n983), .C2(new_n244), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G311), .A2(new_n773), .B1(new_n780), .B2(G317), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT52), .Z(new_n1064));
  NAND2_X1  g0864(.A1(new_n784), .A2(G283), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G107), .A2(new_n794), .B1(new_n788), .B2(G322), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n777), .A2(new_n631), .B1(new_n791), .B2(new_n470), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n254), .B(new_n1067), .C1(G294), .C2(new_n775), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G150), .A2(new_n780), .B1(new_n773), .B2(G159), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT51), .Z(new_n1071));
  AOI21_X1  g0871(.A(new_n968), .B1(new_n811), .B2(new_n357), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n838), .B1(G143), .B2(new_n788), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n959), .A2(G50), .B1(new_n803), .B2(G77), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n783), .A2(new_n310), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1069), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n754), .B1(new_n1077), .B2(new_n763), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1061), .A2(new_n1062), .A3(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1002), .B(KEYINPUT113), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n990), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT114), .B1(new_n1002), .B2(new_n1022), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n709), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1002), .A2(new_n1022), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1002), .A2(KEYINPUT114), .A3(new_n1022), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1081), .A2(new_n1086), .ZN(G390));
  NOR3_X1   g0887(.A1(new_n893), .A2(new_n894), .A3(new_n927), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n823), .A2(new_n374), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n819), .B1(new_n943), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n905), .B(KEYINPUT115), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n904), .B1(new_n930), .B2(new_n905), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n925), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n824), .A2(G330), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n748), .A2(new_n932), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n899), .B2(new_n900), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(KEYINPUT116), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1092), .A2(new_n1094), .A3(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n932), .B(new_n1096), .C1(new_n899), .C2(new_n900), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT116), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n990), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n254), .B1(new_n780), .B2(G283), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1108), .B(new_n805), .C1(new_n203), .C2(new_n777), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G68), .B2(new_n794), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n788), .A2(G294), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n773), .A2(G116), .B1(G77), .B2(new_n803), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT119), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n811), .A2(G97), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1110), .A2(new_n1111), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n797), .A2(new_n857), .B1(new_n791), .B2(new_n850), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT54), .B(G143), .Z(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n811), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n959), .A2(G137), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G50), .A2(new_n794), .B1(new_n788), .B2(G125), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n783), .A2(new_n291), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n254), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1122), .B2(new_n1121), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n801), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1115), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1128), .A2(new_n763), .B1(new_n406), .B2(new_n864), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n866), .B(new_n1129), .C1(new_n926), .C2(new_n765), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1107), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT118), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1092), .A2(new_n1094), .A3(new_n1099), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n690), .B(new_n1089), .C1(new_n719), .C2(new_n723), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n819), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1091), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1138), .A2(new_n1088), .B1(new_n925), .B2(new_n1093), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1133), .B1(new_n1139), .B2(new_n1104), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n901), .A2(new_n459), .A3(G330), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n654), .B(new_n1141), .C1(new_n725), .C2(new_n655), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n742), .B1(KEYINPUT97), .B2(new_n740), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n747), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1095), .B1(new_n1146), .B2(new_n726), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT117), .B1(new_n1147), .B2(new_n932), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n748), .A2(new_n1096), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT117), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(new_n905), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n1101), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n931), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1097), .B1(new_n1098), .B2(new_n1091), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1090), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1143), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1132), .B1(new_n1140), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1152), .A2(new_n931), .B1(new_n1154), .B2(new_n1090), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n1142), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1093), .A2(new_n925), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n921), .A2(KEYINPUT109), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n885), .A2(new_n892), .A3(new_n886), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n904), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1103), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1160), .A2(new_n1166), .A3(KEYINPUT118), .A4(new_n1133), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1158), .A2(new_n1167), .B1(new_n1140), .B2(new_n1157), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1131), .B1(new_n1168), .B2(new_n708), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(G378));
  INV_X1    g0970(.A(KEYINPUT122), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n307), .A2(new_n342), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT55), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n303), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n687), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1172), .B(KEYINPUT55), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n303), .A3(new_n686), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1171), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1179), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(KEYINPUT122), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1182), .A2(new_n1187), .A3(new_n764), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n864), .A2(new_n287), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1117), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1190), .A2(new_n783), .B1(new_n291), .B2(new_n791), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G125), .A2(new_n780), .B1(new_n773), .B2(G128), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n857), .B2(new_n777), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(G137), .C2(new_n775), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT59), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G41), .B1(new_n788), .B2(G124), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G33), .B1(new_n794), .B2(G159), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n794), .A2(G58), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n788), .A2(G283), .ZN(new_n1200));
  AND4_X1   g1000(.A1(new_n251), .A2(new_n1199), .A3(new_n1200), .A4(new_n964), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n797), .A2(new_n203), .B1(new_n801), .B2(new_n950), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G77), .B2(new_n784), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n982), .A2(new_n774), .B1(new_n202), .B2(new_n777), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT120), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1201), .A2(new_n968), .A3(new_n1203), .A4(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT58), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G41), .B1(new_n392), .B2(G33), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1198), .B(new_n1207), .C1(G50), .C2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n754), .B1(new_n1209), .B2(new_n763), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1188), .A2(new_n1189), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1213));
  INV_X1    g1013(.A(G330), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n917), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1216), .A2(G330), .A3(new_n916), .A4(new_n908), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT123), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n934), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1218), .B(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1212), .B1(new_n1222), .B2(new_n990), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT118), .B1(new_n1106), .B2(new_n1160), .ZN(new_n1224));
  AND4_X1   g1024(.A1(KEYINPUT118), .A2(new_n1160), .A3(new_n1166), .A4(new_n1133), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1143), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1226), .B2(new_n1222), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1142), .B1(new_n1158), .B2(new_n1167), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n928), .A2(new_n929), .A3(new_n933), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1218), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1215), .A2(new_n1217), .A3(new_n934), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(KEYINPUT57), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n708), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1223), .B1(new_n1227), .B2(new_n1233), .ZN(G375));
  NAND3_X1  g1034(.A1(new_n1156), .A2(KEYINPUT124), .A3(new_n990), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT124), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1159), .B2(new_n1059), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1199), .B1(new_n850), .B2(new_n783), .C1(new_n856), .C2(new_n1126), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G50), .B2(new_n803), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n773), .A2(G137), .B1(new_n959), .B2(new_n1117), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n291), .B2(new_n774), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(new_n968), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1239), .B(new_n1242), .C1(new_n857), .C2(new_n801), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n777), .A2(new_n470), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n797), .A2(new_n840), .B1(new_n801), .B2(new_n792), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n811), .B2(G107), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n794), .A2(G77), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n262), .B1(new_n783), .B2(new_n202), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n788), .B2(G303), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1041), .A4(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1243), .B1(new_n1244), .B2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1251), .A2(new_n763), .B1(new_n310), .B2(new_n864), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n866), .B(new_n1252), .C1(new_n1137), .C2(new_n765), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1235), .A2(new_n1237), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1235), .A2(new_n1237), .A3(KEYINPUT125), .A4(new_n1253), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1159), .A2(new_n1142), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1157), .A2(new_n1006), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(G381));
  NOR2_X1   g1061(.A1(G390), .A2(G387), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1220), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1211), .B1(new_n1267), .B2(new_n1059), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1230), .A2(KEYINPUT57), .A3(new_n1231), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n709), .B1(new_n1226), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT57), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1228), .B2(new_n1267), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1268), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1169), .ZN(new_n1274));
  INV_X1    g1074(.A(G384), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1258), .A2(new_n1275), .A3(new_n1260), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1264), .A2(new_n1274), .A3(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1277), .A2(KEYINPUT126), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(KEYINPUT126), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1278), .A2(new_n1279), .ZN(G407));
  NAND3_X1  g1080(.A1(new_n1273), .A2(new_n688), .A3(new_n1169), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G213), .B(new_n1281), .C1(new_n1278), .C2(new_n1279), .ZN(G409));
  XOR2_X1   g1082(.A(G393), .B(G396), .Z(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G390), .A2(G387), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1286), .B2(new_n1262), .ZN(new_n1287));
  OR2_X1    g1087(.A1(G390), .A2(G387), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n688), .A2(G213), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1226), .A2(new_n1006), .A3(new_n1222), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1230), .A2(new_n990), .A3(new_n1231), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(new_n1169), .A3(new_n1211), .A4(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1292), .B(new_n1295), .C1(new_n1273), .C2(new_n1169), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1259), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n709), .B1(new_n1298), .B2(KEYINPUT60), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1259), .A2(new_n1297), .A3(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1157), .A3(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1258), .A2(new_n1302), .A3(G384), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G384), .B1(new_n1258), .B2(new_n1302), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(KEYINPUT62), .B1(new_n1296), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n688), .A2(G213), .A3(G2897), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1258), .A2(new_n1302), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1275), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1258), .A2(new_n1302), .A3(G384), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n1315), .A3(new_n1310), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1296), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G375), .A2(G378), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1319), .A2(new_n1305), .A3(new_n1292), .A4(new_n1295), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT62), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1291), .B1(new_n1309), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT61), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1296), .A2(new_n1306), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT63), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n1296), .B2(new_n1317), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1323), .B(new_n1325), .C1(new_n1324), .C2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1322), .A2(new_n1328), .ZN(G405));
  NAND2_X1  g1129(.A1(new_n1319), .A2(new_n1274), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1305), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1319), .A2(new_n1274), .A3(new_n1306), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1290), .ZN(G402));
endmodule


