//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT89), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT2), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G113), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT65), .A2(G116), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT65), .A2(G116), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G116), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n194), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT65), .A2(G116), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT65), .A2(G116), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(G119), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n200), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n191), .A2(new_n193), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n201), .A2(new_n202), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(new_n206), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT66), .A3(new_n194), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G104), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G101), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(G101), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n213), .A2(new_n216), .A3(new_n222), .A4(new_n217), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(KEYINPUT4), .A3(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n209), .A2(new_n211), .A3(new_n220), .A4(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT88), .A2(KEYINPUT5), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT88), .A2(KEYINPUT5), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n190), .B1(new_n228), .B2(new_n200), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n210), .B2(new_n228), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n212), .A2(G107), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n215), .A2(G104), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT83), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n223), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n223), .B2(new_n233), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n230), .B(new_n208), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n225), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT6), .ZN(new_n239));
  XNOR2_X1  g053(.A(G110), .B(G122), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n225), .A2(new_n237), .A3(new_n240), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT6), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n240), .B1(new_n225), .B2(new_n237), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n189), .B(new_n242), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n245), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(KEYINPUT89), .A3(KEYINPUT6), .A4(new_n243), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT1), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G128), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(KEYINPUT1), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n250), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT64), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n253), .A2(KEYINPUT64), .A3(new_n256), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n254), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n257), .A2(new_n259), .A3(new_n267), .ZN(new_n268));
  OR2_X1    g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n268), .B1(new_n271), .B2(new_n253), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G125), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G224), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(G953), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n274), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n249), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT90), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n240), .B(KEYINPUT8), .Z(new_n284));
  NAND2_X1  g098(.A1(new_n223), .A2(new_n233), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n230), .B2(new_n208), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(KEYINPUT83), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n223), .A2(new_n233), .A3(new_n234), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT5), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n229), .B1(new_n210), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n208), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT91), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n287), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n290), .A2(KEYINPUT91), .A3(new_n208), .A4(new_n292), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT7), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n274), .B1(new_n298), .B2(new_n276), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n273), .A4(new_n277), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n243), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n283), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n278), .B1(new_n246), .B2(new_n248), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(KEYINPUT90), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n282), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT92), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT92), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n309), .B(new_n306), .C1(new_n282), .C2(new_n304), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n282), .A2(new_n304), .A3(new_n306), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n188), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G217), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT74), .B(G902), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G234), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT76), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n265), .A2(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(G146), .B(new_n320), .C1(new_n323), .C2(new_n318), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G125), .B(G140), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n324), .B1(new_n330), .B2(G146), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n197), .A2(G128), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n255), .A2(KEYINPUT23), .A3(G119), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n197), .A2(G128), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n332), .B(new_n333), .C1(new_n334), .C2(KEYINPUT23), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G110), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT24), .B(G110), .ZN(new_n337));
  OR3_X1    g151(.A1(new_n255), .A2(KEYINPUT77), .A3(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n338), .B(new_n339), .C1(new_n197), .C2(G128), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n336), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n320), .B1(new_n323), .B2(new_n318), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n250), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n343), .A2(new_n324), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n335), .A2(G110), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n340), .B2(new_n337), .ZN(new_n346));
  OAI22_X1  g160(.A1(new_n331), .A2(new_n341), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT22), .B(G137), .ZN(new_n348));
  INV_X1    g162(.A(G953), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(G221), .A3(G234), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n348), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n347), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n315), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n354), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n317), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n316), .A2(G902), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n360), .B(KEYINPUT80), .Z(new_n361));
  OR2_X1    g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n257), .A2(new_n259), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n363), .A2(new_n255), .B1(KEYINPUT1), .B2(new_n251), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT64), .B1(new_n253), .B2(new_n256), .ZN(new_n365));
  AND4_X1   g179(.A1(KEYINPUT64), .A2(new_n256), .A3(new_n257), .A4(new_n259), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT11), .ZN(new_n368));
  INV_X1    g182(.A(G134), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(G137), .ZN(new_n370));
  INV_X1    g184(.A(G137), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT11), .A3(G134), .ZN(new_n372));
  INV_X1    g186(.A(G131), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(G137), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n371), .A2(G134), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n369), .A2(G137), .ZN(new_n377));
  OAI21_X1  g191(.A(G131), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n367), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n370), .A2(new_n374), .A3(new_n372), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G131), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n375), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT67), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n268), .B(new_n386), .C1(new_n271), .C2(new_n253), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n381), .A2(new_n388), .A3(KEYINPUT30), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n262), .A2(new_n263), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n379), .B1(new_n391), .B2(new_n364), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n272), .B1(new_n375), .B2(new_n384), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n209), .A2(new_n211), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n398));
  NOR2_X1   g212(.A1(G237), .A2(G953), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G210), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n398), .B(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT26), .B(G101), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n395), .A2(new_n381), .A3(new_n388), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n397), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT31), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT31), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n397), .A2(new_n408), .A3(new_n404), .A4(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n211), .B(new_n209), .C1(new_n392), .C2(new_n393), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n405), .A3(KEYINPUT69), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT69), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n396), .B(new_n413), .C1(new_n392), .C2(new_n393), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(KEYINPUT28), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT28), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n405), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n404), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT70), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n411), .A2(new_n405), .A3(KEYINPUT69), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT28), .B1(new_n411), .B2(KEYINPUT69), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n417), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n403), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n407), .A4(new_n409), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(G472), .A2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT32), .ZN(new_n429));
  INV_X1    g243(.A(new_n427), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n419), .B2(new_n425), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT32), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n381), .A2(new_n388), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n396), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n395), .A2(new_n381), .A3(new_n388), .A4(KEYINPUT71), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n387), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n258), .A2(G146), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n270), .B(new_n269), .C1(new_n440), .C2(new_n251), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n386), .B1(new_n441), .B2(new_n268), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n392), .B1(new_n443), .B2(new_n385), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT71), .B1(new_n444), .B2(new_n395), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT28), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT72), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT73), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n417), .B(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n405), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n436), .A3(new_n437), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT72), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT28), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n404), .A2(KEYINPUT29), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n447), .A2(new_n449), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n315), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT75), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(KEYINPUT75), .A3(new_n315), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n415), .A2(new_n404), .A3(new_n417), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n397), .A2(new_n405), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT29), .B1(new_n462), .B2(new_n403), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G472), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n362), .B1(new_n434), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G237), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(new_n349), .A3(G214), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n258), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n399), .B(G214), .C1(KEYINPUT93), .C2(G143), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G131), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT17), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n373), .A3(new_n472), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(KEYINPUT17), .A3(G131), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT95), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n373), .B1(new_n471), .B2(new_n472), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT95), .B1(new_n481), .B2(KEYINPUT17), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n344), .B(new_n477), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G113), .B(G122), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(new_n212), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT18), .A2(G131), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n471), .A2(new_n486), .A3(new_n472), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n473), .A2(KEYINPUT18), .A3(G131), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n326), .A2(new_n328), .A3(G146), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n327), .A2(new_n250), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n483), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n474), .A2(new_n476), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n323), .A2(new_n325), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT19), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n323), .A2(KEYINPUT94), .A3(KEYINPUT19), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n327), .B2(new_n496), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n324), .B(new_n493), .C1(new_n501), .C2(G146), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n502), .A2(new_n491), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n492), .B1(new_n503), .B2(new_n485), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT20), .ZN(new_n505));
  NOR2_X1   g319(.A1(G475), .A2(G902), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT96), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n504), .A2(new_n509), .A3(new_n505), .A4(new_n506), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n485), .B1(new_n502), .B2(new_n491), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n490), .B1(new_n329), .B2(new_n250), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n488), .A2(new_n487), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n344), .A2(new_n477), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n478), .B(new_n479), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n511), .B1(new_n517), .B2(new_n485), .ZN(new_n518));
  INV_X1    g332(.A(new_n506), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT20), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n508), .A2(new_n510), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n492), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n485), .B1(new_n483), .B2(new_n491), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n283), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G475), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n203), .A2(G122), .A3(new_n204), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n199), .A2(G122), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n215), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n258), .A2(G128), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n255), .A2(G143), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n533), .A2(new_n534), .A3(G134), .ZN(new_n535));
  AOI21_X1  g349(.A(G134), .B1(new_n533), .B2(new_n534), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n530), .A2(new_n538), .A3(new_n531), .ZN(new_n539));
  OAI21_X1  g353(.A(G107), .B1(new_n530), .B2(new_n538), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n532), .B(new_n537), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n533), .A2(new_n534), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT13), .B1(new_n255), .B2(G143), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n369), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT13), .A4(G134), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n530), .A2(new_n215), .A3(new_n531), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n215), .B1(new_n530), .B2(new_n531), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT9), .B(G234), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n550), .A2(new_n314), .A3(G953), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n541), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n551), .B1(new_n541), .B2(new_n549), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n315), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT97), .B(new_n315), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n529), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n528), .B1(new_n554), .B2(new_n555), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT98), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT98), .B1(new_n558), .B2(new_n559), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G952), .ZN(new_n565));
  AOI211_X1 g379(.A(G953), .B(new_n565), .C1(G234), .C2(G237), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n349), .B(new_n315), .C1(G234), .C2(G237), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n526), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G221), .B1(new_n550), .B2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n385), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n264), .A2(KEYINPUT82), .A3(new_n285), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT82), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n367), .B2(new_n286), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n574), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n367), .B(KEYINPUT10), .C1(new_n235), .C2(new_n236), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n224), .A2(new_n387), .A3(new_n382), .A4(new_n220), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n573), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT82), .B1(new_n264), .B2(new_n285), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n367), .A2(new_n576), .A3(new_n286), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT10), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n580), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n585), .A2(new_n586), .A3(new_n385), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n349), .A2(G227), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT81), .ZN(new_n589));
  XNOR2_X1  g403(.A(G110), .B(G140), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n582), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT85), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n290), .B2(new_n367), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n264), .A2(new_n288), .A3(KEYINPUT85), .A4(new_n289), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n595), .B(new_n596), .C1(new_n575), .C2(new_n577), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT12), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n578), .A2(new_n581), .A3(new_n573), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n597), .A2(new_n602), .A3(new_n598), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n593), .B1(new_n604), .B2(new_n592), .ZN(new_n605));
  OAI21_X1  g419(.A(G469), .B1(new_n605), .B2(G902), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT87), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n587), .B2(new_n592), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n601), .A2(KEYINPUT87), .A3(new_n591), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n600), .A3(new_n603), .A4(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n592), .B1(new_n582), .B2(new_n587), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT86), .B(G469), .Z(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n315), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n572), .B1(new_n606), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n570), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n313), .A2(new_n467), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  NAND3_X1  g432(.A1(new_n249), .A2(KEYINPUT90), .A3(new_n279), .ZN(new_n619));
  INV_X1    g433(.A(new_n302), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n303), .A2(KEYINPUT90), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n307), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n188), .B1(new_n623), .B2(new_n312), .ZN(new_n624));
  INV_X1    g438(.A(new_n569), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n552), .A2(new_n553), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT33), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(G478), .A3(new_n315), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n554), .A2(new_n527), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n526), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n624), .A2(new_n625), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n426), .A2(new_n315), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n431), .B1(new_n635), .B2(G472), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n358), .A2(new_n361), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n636), .A2(new_n637), .A3(new_n615), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n520), .A2(new_n507), .B1(G475), .B2(new_n524), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n556), .A2(new_n557), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n528), .ZN(new_n645));
  INV_X1    g459(.A(new_n559), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n561), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n558), .A2(KEYINPUT98), .A3(new_n559), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n643), .B(new_n625), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT99), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n564), .A2(new_n651), .A3(new_n625), .A4(new_n643), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n621), .A2(new_n307), .A3(new_n622), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n306), .B1(new_n282), .B2(new_n304), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n187), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n642), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n624), .A2(KEYINPUT100), .A3(new_n650), .A4(new_n652), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n638), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NAND2_X1  g476(.A1(new_n635), .A2(G472), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n428), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n347), .B(KEYINPUT101), .Z(new_n665));
  INV_X1    g479(.A(KEYINPUT36), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n351), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n665), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n359), .ZN(new_n669));
  INV_X1    g483(.A(new_n357), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n355), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n669), .B1(new_n671), .B2(new_n317), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n664), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n313), .A2(new_n616), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  NAND2_X1  g491(.A1(new_n434), .A2(new_n466), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n520), .A2(new_n507), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n525), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n563), .B2(new_n562), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n566), .B1(new_n567), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n656), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n678), .A2(new_n686), .A3(new_n615), .A4(new_n672), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  NAND2_X1  g502(.A1(new_n462), .A2(new_n404), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n283), .B1(new_n452), .B2(new_n404), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n434), .A2(KEYINPUT102), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT102), .B1(new_n434), .B2(new_n692), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n623), .A2(new_n309), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n655), .A2(KEYINPUT92), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n312), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT38), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n526), .A2(new_n564), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n673), .A2(new_n187), .A3(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n696), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n683), .B(KEYINPUT39), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n615), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT103), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT40), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n704), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  AOI21_X1  g526(.A(new_n432), .B1(new_n426), .B2(new_n427), .ZN(new_n713));
  AOI211_X1 g527(.A(KEYINPUT32), .B(new_n430), .C1(new_n419), .C2(new_n425), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(G472), .ZN(new_n716));
  INV_X1    g530(.A(new_n464), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n457), .B2(new_n458), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n716), .B1(new_n718), .B2(new_n460), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n615), .B(new_n672), .C1(new_n715), .C2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n526), .A2(new_n630), .A3(new_n684), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n624), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n723), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT104), .B1(new_n725), .B2(new_n656), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n721), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  INV_X1    g542(.A(new_n315), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n610), .B2(new_n611), .ZN(new_n730));
  INV_X1    g544(.A(G469), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n613), .ZN(new_n733));
  AOI211_X1 g547(.A(new_n729), .B(new_n733), .C1(new_n610), .C2(new_n611), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n732), .A2(new_n734), .A3(new_n572), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n467), .A2(new_n634), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  OAI211_X1 g552(.A(new_n637), .B(new_n735), .C1(new_n715), .C2(new_n719), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n659), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  OAI211_X1 g556(.A(new_n614), .B(new_n571), .C1(new_n731), .C2(new_n730), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n656), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n678), .A2(new_n744), .A3(new_n570), .A4(new_n672), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  NAND2_X1  g560(.A1(new_n449), .A2(new_n454), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n453), .B1(new_n452), .B2(KEYINPUT28), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n403), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n410), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n430), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n635), .B2(G472), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n735), .A2(new_n752), .A3(new_n637), .A4(new_n625), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n624), .A2(new_n702), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  AND2_X1   g570(.A1(new_n752), .A2(new_n672), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n744), .A3(new_n723), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G125), .ZN(G27));
  AND2_X1   g573(.A1(new_n312), .A2(new_n187), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n697), .A2(new_n615), .A3(new_n760), .A4(new_n698), .ZN(new_n761));
  NOR2_X1   g575(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n467), .A2(new_n761), .A3(new_n723), .A4(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n637), .B1(new_n715), .B2(new_n719), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n615), .A2(new_n760), .A3(new_n697), .A4(new_n698), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n765), .A2(new_n725), .A3(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n768));
  OAI21_X1  g582(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT106), .B(G131), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G33));
  NOR3_X1   g585(.A1(new_n765), .A2(new_n685), .A3(new_n766), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n369), .ZN(G36));
  INV_X1    g587(.A(new_n526), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n630), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT43), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n777), .A3(new_n630), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n664), .A3(new_n672), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n760), .A2(new_n697), .A3(new_n698), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT107), .Z(new_n784));
  NAND4_X1  g598(.A1(new_n779), .A2(KEYINPUT44), .A3(new_n664), .A4(new_n672), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n731), .A2(new_n283), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n605), .A2(KEYINPUT45), .ZN(new_n789));
  OAI21_X1  g603(.A(G469), .B1(new_n605), .B2(KEYINPUT45), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n734), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n571), .A3(new_n705), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n786), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(new_n371), .ZN(G39));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n571), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT47), .ZN(new_n799));
  OR4_X1    g613(.A1(new_n678), .A2(new_n783), .A3(new_n637), .A4(new_n725), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n319), .ZN(G42));
  NOR2_X1   g616(.A1(G952), .A2(G953), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n467), .A2(new_n761), .A3(new_n723), .ZN(new_n804));
  INV_X1    g618(.A(new_n768), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n772), .B1(new_n806), .B2(new_n764), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n313), .B(new_n616), .C1(new_n467), .C2(new_n674), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n741), .A2(new_n808), .A3(new_n736), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n672), .B1(new_n715), .B2(new_n719), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n735), .A2(new_n624), .A3(new_n570), .ZN(new_n811));
  OAI22_X1  g625(.A1(new_n810), .A2(new_n811), .B1(new_n753), .B2(new_n754), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n521), .B(new_n525), .C1(new_n558), .C2(new_n559), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n569), .B1(new_n631), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n636), .A3(new_n637), .A4(new_n615), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n699), .A2(new_n187), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n752), .A2(new_n672), .A3(new_n723), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n766), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n643), .A2(new_n560), .A3(new_n684), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT109), .Z(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n783), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(new_n721), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n807), .A2(new_n809), .A3(new_n818), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n673), .A2(new_n615), .A3(new_n684), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n754), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n830), .B1(new_n694), .B2(new_n695), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n726), .A2(new_n724), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n687), .B(new_n758), .C1(new_n833), .C2(new_n720), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n828), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n687), .A2(new_n758), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n831), .A3(new_n727), .A4(KEYINPUT52), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n827), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n741), .A2(new_n808), .A3(new_n736), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n313), .A2(new_n638), .A3(new_n814), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n755), .A3(new_n745), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(KEYINPUT110), .A3(new_n807), .A4(new_n824), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n740), .B1(new_n659), .B2(new_n634), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n818), .A2(new_n808), .A3(new_n845), .A4(new_n824), .ZN(new_n846));
  INV_X1    g660(.A(new_n772), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n769), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n844), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n835), .A2(new_n837), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n843), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n852));
  AOI221_X4 g666(.A(KEYINPUT54), .B1(new_n826), .B2(new_n838), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n825), .A2(new_n844), .B1(new_n835), .B2(new_n837), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  INV_X1    g669(.A(new_n852), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n843), .A4(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n843), .A2(new_n849), .A3(new_n850), .A4(new_n856), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT112), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n851), .A2(new_n827), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n853), .B1(KEYINPUT54), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n614), .B1(new_n731), .B2(new_n730), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n863), .A2(new_n571), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n799), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n776), .A2(new_n566), .A3(new_n778), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n752), .A2(new_n637), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n784), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n869), .A2(KEYINPUT51), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n783), .A2(new_n743), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n637), .A2(new_n566), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n526), .A2(new_n630), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n696), .A2(new_n871), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n866), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n757), .A3(new_n871), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT113), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n743), .A2(new_n187), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n701), .A2(new_n868), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n880), .B(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n874), .A2(new_n883), .A3(new_n876), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n878), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n885), .A2(KEYINPUT114), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(KEYINPUT114), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n870), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n868), .A2(new_n744), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n889), .A2(KEYINPUT115), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(KEYINPUT115), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n890), .A2(new_n891), .A3(new_n565), .A4(G953), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n875), .A2(new_n467), .A3(new_n871), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT48), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n696), .A2(new_n632), .A3(new_n871), .A4(new_n872), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n877), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n869), .A2(new_n897), .A3(new_n882), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n888), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n803), .B1(new_n862), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n637), .A2(new_n187), .A3(new_n571), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n775), .B(new_n904), .C1(KEYINPUT49), .C2(new_n863), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n863), .A2(KEYINPUT49), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT108), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n696), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n701), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT116), .B1(new_n903), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT116), .ZN(new_n912));
  INV_X1    g726(.A(new_n910), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n858), .A2(KEYINPUT112), .B1(new_n851), .B2(new_n827), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n857), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n916), .A2(new_n901), .A3(new_n853), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n912), .B(new_n913), .C1(new_n917), .C2(new_n803), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n911), .A2(new_n918), .ZN(G75));
  NAND2_X1  g733(.A1(new_n565), .A2(G953), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT118), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n851), .A2(new_n852), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n826), .A2(new_n838), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n315), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT56), .B1(new_n924), .B2(new_n307), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n249), .A2(new_n279), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n303), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n921), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n925), .A2(new_n928), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT117), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n925), .A2(KEYINPUT117), .A3(new_n928), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G51));
  INV_X1    g748(.A(new_n921), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n922), .A2(new_n923), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n914), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n853), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n787), .B(KEYINPUT57), .Z(new_n939));
  OAI21_X1  g753(.A(new_n612), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n789), .A2(new_n790), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n924), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n935), .B1(new_n940), .B2(new_n942), .ZN(G54));
  NAND3_X1  g757(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(new_n504), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n504), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n935), .B1(new_n945), .B2(new_n946), .ZN(G60));
  XNOR2_X1  g761(.A(new_n627), .B(KEYINPUT119), .ZN(new_n948));
  NAND2_X1  g762(.A1(G478), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT59), .Z(new_n950));
  OR2_X1    g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n921), .B1(new_n938), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n950), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n916), .B2(new_n853), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n948), .B2(new_n954), .ZN(G63));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT120), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n936), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n668), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n921), .B1(new_n960), .B2(new_n352), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n956), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n960), .A2(new_n352), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n965), .A2(KEYINPUT61), .A3(new_n921), .A4(new_n961), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(G66));
  OAI21_X1  g781(.A(G953), .B1(new_n568), .B2(new_n275), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n842), .B2(G953), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n246), .B(new_n248), .C1(G898), .C2(new_n349), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  XNOR2_X1  g785(.A(new_n834), .B(KEYINPUT122), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n711), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n631), .A2(new_n813), .ZN(new_n976));
  AND4_X1   g790(.A1(new_n467), .A2(new_n761), .A3(new_n705), .A4(new_n976), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n801), .A2(new_n796), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n974), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n349), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n501), .B(KEYINPUT121), .Z(new_n981));
  NAND2_X1  g795(.A1(new_n389), .A2(new_n394), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n467), .A2(new_n624), .A3(new_n702), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n795), .B1(new_n786), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n801), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n807), .B(KEYINPUT123), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n972), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(G900), .A2(G953), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n983), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n985), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n983), .B1(new_n979), .B2(new_n349), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n991), .A2(new_n993), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT125), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(G227), .ZN(new_n1001));
  OAI21_X1  g815(.A(G953), .B1(new_n1001), .B2(new_n682), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n983), .B2(KEYINPUT124), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n996), .A2(new_n1003), .A3(new_n999), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  INV_X1    g823(.A(new_n842), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n990), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n462), .A2(new_n404), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n935), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n974), .A2(new_n842), .A3(new_n975), .A4(new_n978), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n1009), .ZN(new_n1015));
  AOI21_X1  g829(.A(KEYINPUT126), .B1(new_n1015), .B2(new_n690), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT126), .ZN(new_n1017));
  AOI211_X1 g831(.A(new_n1017), .B(new_n689), .C1(new_n1014), .C2(new_n1009), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1013), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1012), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1020), .A2(new_n689), .A3(new_n1009), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT127), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1019), .B1(new_n861), .B2(new_n1022), .ZN(G57));
endmodule


