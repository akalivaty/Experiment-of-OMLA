//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  XOR2_X1   g000(.A(KEYINPUT26), .B(G101), .Z(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT29), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT2), .B(G113), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n197), .A2(new_n199), .A3(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n197), .B2(new_n199), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n206), .B2(new_n201), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT0), .A4(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT64), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT0), .A4(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(new_n211), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT0), .B(G128), .Z(new_n218));
  AOI22_X1  g032(.A1(new_n213), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT11), .B1(new_n220), .B2(G137), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT11), .ZN(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G134), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT65), .B(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n220), .A2(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n221), .A2(new_n224), .B1(new_n220), .B2(G137), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n214), .A2(new_n233), .A3(G128), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n209), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT68), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(KEYINPUT67), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n238), .B(new_n209), .C1(new_n240), .C2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n237), .A2(G128), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n235), .B1(new_n244), .B2(new_n217), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n227), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n223), .A2(G134), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n227), .A2(new_n246), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n228), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n207), .B(new_n232), .C1(new_n245), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT72), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n251), .A2(new_n228), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n209), .B1(new_n240), .B2(new_n242), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(KEYINPUT68), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n214), .B1(new_n258), .B2(new_n243), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n255), .B1(new_n259), .B2(new_n235), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n207), .A4(new_n232), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n206), .A2(new_n201), .ZN(new_n263));
  INV_X1    g077(.A(new_n202), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n241), .A2(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n266), .A2(new_n267), .B1(G143), .B2(new_n208), .ZN(new_n268));
  OAI21_X1  g082(.A(G128), .B1(new_n268), .B2(new_n238), .ZN(new_n269));
  INV_X1    g083(.A(new_n243), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n217), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n252), .B1(new_n271), .B2(new_n234), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n219), .A2(new_n231), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n265), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n254), .A2(new_n262), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT28), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(KEYINPUT73), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n253), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT73), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n275), .B2(KEYINPUT28), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n195), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n260), .A2(KEYINPUT28), .A3(new_n207), .A4(new_n232), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n284), .A3(new_n274), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n285), .A2(new_n193), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT30), .B1(new_n272), .B2(new_n273), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n288), .B(new_n232), .C1(new_n245), .C2(new_n252), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n207), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n253), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n286), .B(new_n194), .C1(new_n192), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n282), .A2(new_n283), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G472), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n285), .A2(new_n193), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n253), .A2(new_n192), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n287), .A2(new_n289), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(new_n265), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT31), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n288), .B1(new_n260), .B2(new_n232), .ZN(new_n302));
  INV_X1    g116(.A(new_n289), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n265), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n297), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n299), .A2(KEYINPUT71), .A3(new_n300), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n301), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(G472), .A2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n310), .A2(KEYINPUT32), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT32), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n304), .A2(new_n305), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n315), .A2(KEYINPUT31), .B1(new_n193), .B2(new_n285), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT71), .B1(new_n299), .B2(new_n300), .ZN(new_n317));
  NOR4_X1   g131(.A1(new_n290), .A2(new_n307), .A3(KEYINPUT31), .A4(new_n297), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n314), .B1(new_n319), .B2(new_n311), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n295), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G140), .ZN(new_n322));
  INV_X1    g136(.A(G953), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n323), .A2(G227), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n322), .B(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT84), .ZN(new_n326));
  INV_X1    g140(.A(G104), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT3), .B1(new_n327), .B2(G107), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n329));
  INV_X1    g143(.A(G107), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G104), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(G107), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(G101), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT82), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT82), .A4(G101), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(G101), .ZN(new_n340));
  INV_X1    g154(.A(G101), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n328), .A2(new_n331), .A3(new_n341), .A4(new_n332), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(KEYINPUT4), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n219), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n327), .A2(G107), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n330), .A2(G104), .ZN(new_n347));
  OAI21_X1  g161(.A(G101), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n211), .A2(new_n241), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n256), .B2(new_n217), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n349), .B1(new_n234), .B2(new_n354), .ZN(new_n355));
  OAI22_X1  g169(.A1(new_n245), .A2(new_n352), .B1(new_n355), .B2(KEYINPUT10), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n326), .B(new_n231), .C1(new_n345), .C2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n351), .B1(new_n259), .B2(new_n235), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n234), .ZN(new_n359));
  INV_X1    g173(.A(new_n349), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n350), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n231), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n228), .B(KEYINPUT83), .C1(new_n229), .C2(new_n230), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n358), .A2(new_n344), .A3(new_n362), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT84), .ZN(new_n368));
  INV_X1    g182(.A(new_n231), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT10), .B1(new_n359), .B2(new_n360), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n271), .A2(new_n234), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(new_n351), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n369), .B1(new_n372), .B2(new_n344), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n325), .B(new_n357), .C1(new_n368), .C2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n361), .B1(new_n371), .B2(new_n360), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT12), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n231), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n355), .B1(new_n245), .B2(new_n349), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT12), .B1(new_n378), .B2(new_n369), .ZN(new_n379));
  INV_X1    g193(.A(new_n325), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n377), .A2(new_n379), .A3(new_n367), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G469), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n283), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n283), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n357), .B1(new_n368), .B2(new_n373), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n380), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n379), .A3(new_n367), .ZN(new_n389));
  XOR2_X1   g203(.A(new_n325), .B(KEYINPUT80), .Z(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(G469), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n384), .A2(new_n386), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT9), .B(G234), .ZN(new_n394));
  OAI21_X1  g208(.A(G221), .B1(new_n394), .B2(G902), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G214), .B1(G237), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n198), .A2(G119), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n196), .A2(G116), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT69), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n197), .A2(new_n199), .A3(new_n203), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G113), .B1(new_n197), .B2(KEYINPUT5), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT85), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT5), .B1(new_n204), .B2(new_n205), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n407));
  INV_X1    g221(.A(new_n404), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n202), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT88), .B1(new_n410), .B2(new_n360), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n403), .A2(KEYINPUT85), .A3(new_n404), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n264), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n349), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n349), .A2(new_n202), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n408), .B1(new_n398), .B2(new_n200), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G122), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT8), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT87), .B(G224), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n424), .A2(G953), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT7), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n259), .A2(G125), .A3(new_n235), .ZN(new_n427));
  INV_X1    g241(.A(G125), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n219), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n426), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n429), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n245), .A2(new_n428), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT7), .A4(new_n425), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n417), .B1(new_n412), .B2(new_n413), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n265), .A2(new_n339), .A3(new_n343), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n421), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n430), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n423), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n429), .B1(new_n428), .B2(new_n245), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n425), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n435), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n421), .B(KEYINPUT86), .Z(new_n442));
  AOI22_X1  g256(.A1(new_n436), .A2(KEYINPUT6), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n442), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G210), .B1(G237), .B2(G902), .ZN(new_n446));
  AND4_X1   g260(.A1(new_n283), .A2(new_n438), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(G902), .B1(new_n423), .B2(new_n437), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n448), .B2(new_n445), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n397), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n396), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n323), .A2(G221), .A3(G234), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT78), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G137), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G125), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n428), .A2(G140), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT76), .ZN(new_n460));
  OR3_X1    g274(.A1(new_n457), .A2(KEYINPUT76), .A3(G125), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT16), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT16), .B1(new_n457), .B2(G125), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n208), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT77), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI211_X1 g281(.A(KEYINPUT77), .B(new_n208), .C1(new_n462), .C2(new_n464), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT75), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n196), .B2(G128), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n256), .A2(KEYINPUT75), .A3(G119), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n196), .A2(G128), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT24), .B(G110), .Z(new_n474));
  NAND3_X1  g288(.A1(new_n256), .A2(KEYINPUT23), .A3(G119), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n196), .A2(G128), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n472), .B(new_n475), .C1(new_n476), .C2(KEYINPUT23), .ZN(new_n477));
  OAI22_X1  g291(.A1(new_n473), .A2(new_n474), .B1(new_n477), .B2(G110), .ZN(new_n478));
  XNOR2_X1  g292(.A(G125), .B(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n208), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n467), .A2(new_n468), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n473), .A2(new_n474), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(G110), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n457), .A2(KEYINPUT76), .A3(G125), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n479), .B2(KEYINPUT76), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n463), .B1(new_n487), .B2(KEYINPUT16), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n208), .ZN(new_n489));
  INV_X1    g303(.A(new_n465), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n456), .B1(new_n482), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT77), .B1(new_n488), .B2(new_n208), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n465), .A2(new_n466), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n480), .A4(new_n478), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n462), .A2(new_n464), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G146), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n483), .B(new_n484), .C1(new_n497), .C2(new_n465), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n498), .A3(new_n455), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n492), .A2(new_n283), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n492), .A2(KEYINPUT25), .A3(new_n499), .A4(new_n283), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G234), .ZN(new_n505));
  OAI21_X1  g319(.A(G217), .B1(new_n505), .B2(G902), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT74), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n492), .A2(new_n499), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n505), .B2(G217), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(KEYINPUT79), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT79), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n507), .B1(new_n502), .B2(new_n503), .ZN(new_n515));
  INV_X1    g329(.A(new_n512), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n520));
  INV_X1    g334(.A(G475), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n283), .ZN(new_n522));
  AND2_X1   g336(.A1(KEYINPUT89), .A2(G143), .ZN(new_n523));
  NOR2_X1   g337(.A1(KEYINPUT89), .A2(G143), .ZN(new_n524));
  OAI211_X1 g338(.A(G214), .B(new_n188), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G237), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n323), .A3(G214), .ZN(new_n527));
  NAND2_X1  g341(.A1(KEYINPUT89), .A2(G143), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(KEYINPUT90), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(KEYINPUT18), .A2(G131), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n487), .A2(G146), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n480), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n493), .A2(new_n494), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n525), .A2(new_n226), .A3(new_n529), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n226), .B1(new_n525), .B2(new_n529), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT91), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n525), .A2(new_n529), .ZN(new_n542));
  INV_X1    g356(.A(new_n226), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n525), .A2(new_n226), .A3(new_n529), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n460), .B2(new_n461), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n479), .A2(KEYINPUT19), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n208), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n541), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n537), .B1(new_n538), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(G113), .B(G122), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(new_n327), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n540), .A2(KEYINPUT17), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n539), .A2(new_n540), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n497), .A2(new_n465), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n555), .B(KEYINPUT92), .Z(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n537), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n522), .B1(new_n557), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT20), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n520), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n532), .A2(new_n533), .B1(new_n480), .B2(new_n535), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n561), .B2(new_n562), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n556), .A2(new_n553), .B1(new_n570), .B2(new_n564), .ZN(new_n571));
  OAI211_X1 g385(.A(KEYINPUT93), .B(KEYINPUT20), .C1(new_n571), .C2(new_n522), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n522), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n521), .A2(new_n283), .A3(KEYINPUT94), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n567), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n573), .B1(new_n571), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n557), .A2(new_n565), .ZN(new_n579));
  INV_X1    g393(.A(new_n577), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(KEYINPUT95), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n568), .A2(new_n572), .A3(new_n578), .A4(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n563), .A2(new_n537), .A3(new_n564), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n555), .B1(new_n563), .B2(new_n537), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n283), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT96), .B(G475), .Z(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT15), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G217), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n394), .A2(new_n593), .A3(G953), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n210), .A2(KEYINPUT13), .A3(G128), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n256), .A2(G143), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(KEYINPUT97), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT13), .B1(new_n210), .B2(G128), .ZN(new_n598));
  OAI221_X1 g412(.A(G134), .B1(KEYINPUT97), .B2(new_n595), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(G116), .B(G122), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n330), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n210), .A2(G128), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(new_n596), .A3(new_n220), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n599), .A2(new_n601), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n602), .A2(new_n596), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G134), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n609), .A2(new_n603), .B1(new_n330), .B2(new_n600), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n198), .A2(KEYINPUT14), .A3(G122), .ZN(new_n611));
  INV_X1    g425(.A(new_n600), .ZN(new_n612));
  OAI211_X1 g426(.A(G107), .B(new_n611), .C1(new_n612), .C2(KEYINPUT14), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n594), .B1(new_n607), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n607), .A2(new_n614), .A3(new_n594), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n592), .B1(new_n618), .B2(new_n283), .ZN(new_n619));
  AOI211_X1 g433(.A(G902), .B(new_n591), .C1(new_n616), .C2(new_n617), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n589), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n617), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n615), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n591), .B1(new_n623), .B2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n618), .A2(new_n283), .A3(new_n592), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT99), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n323), .A2(G952), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n505), .B2(new_n526), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n283), .B(new_n323), .C1(G234), .C2(G237), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT21), .B(G898), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n588), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n321), .A2(new_n451), .A3(new_n519), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  NAND2_X1  g451(.A1(new_n319), .A2(new_n311), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n308), .A2(new_n309), .ZN(new_n639));
  AOI21_X1  g453(.A(G902), .B1(new_n639), .B2(new_n316), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n393), .A2(new_n513), .A3(new_n517), .A4(new_n395), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n634), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n397), .B(new_n645), .C1(new_n447), .C2(new_n449), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n618), .A2(new_n590), .A3(new_n283), .ZN(new_n649));
  NAND2_X1  g463(.A1(G478), .A2(G902), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT33), .B1(new_n594), .B2(KEYINPUT100), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n623), .B(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n649), .B(new_n650), .C1(new_n652), .C2(new_n590), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n582), .B2(new_n587), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT101), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n654), .A2(KEYINPUT101), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT34), .B(G104), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  AND3_X1   g475(.A1(new_n587), .A2(new_n621), .A3(new_n626), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n566), .A2(new_n567), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n568), .A2(new_n572), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n648), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT35), .B(G107), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  INV_X1    g482(.A(new_n642), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n495), .A2(new_n498), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n456), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n515), .B1(new_n511), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n669), .A2(new_n451), .A3(new_n635), .A4(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  OAI21_X1  g491(.A(KEYINPUT32), .B1(new_n310), .B2(new_n312), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n319), .A2(new_n314), .A3(new_n311), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n678), .A2(new_n679), .B1(G472), .B2(new_n294), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n680), .A2(new_n396), .A3(new_n673), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n632), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n630), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n662), .A2(new_n664), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n397), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n438), .A2(new_n445), .A3(new_n283), .ZN(new_n687));
  INV_X1    g501(.A(new_n446), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n448), .A2(new_n446), .A3(new_n445), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n686), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n685), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n662), .A2(new_n664), .A3(new_n684), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT102), .B1(new_n450), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n681), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  INV_X1    g512(.A(new_n396), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n684), .B(KEYINPUT39), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n678), .A2(new_n679), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n299), .B1(new_n275), .B2(new_n193), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n704), .B2(G902), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n674), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n689), .A2(new_n690), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT38), .Z(new_n709));
  AOI21_X1  g523(.A(new_n627), .B1(new_n582), .B2(new_n587), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n397), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n702), .A2(new_n707), .A3(new_n709), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n210), .ZN(G45));
  INV_X1    g527(.A(new_n653), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n588), .A2(new_n714), .A3(new_n684), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n321), .A2(new_n716), .A3(new_n451), .A4(new_n674), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  OAI21_X1  g532(.A(new_n647), .B1(new_n656), .B2(new_n657), .ZN(new_n719));
  AOI21_X1  g533(.A(G902), .B1(new_n374), .B2(new_n381), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n720), .A2(new_n383), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n395), .A3(new_n384), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n321), .A2(new_n519), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT103), .B1(new_n719), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n654), .A2(KEYINPUT101), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n646), .B1(new_n726), .B2(new_n655), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n680), .A2(new_n518), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n723), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT104), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n731), .B(new_n733), .ZN(G15));
  NOR2_X1   g548(.A1(new_n646), .A2(new_n665), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n321), .A2(new_n735), .A3(new_n519), .A4(new_n723), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  NOR2_X1   g551(.A1(new_n722), .A2(new_n450), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n321), .A2(new_n738), .A3(new_n635), .A4(new_n674), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  OAI21_X1  g554(.A(G472), .B1(new_n310), .B2(G902), .ZN(new_n741));
  OAI22_X1  g555(.A1(new_n317), .A2(new_n318), .B1(new_n300), .B2(new_n299), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n277), .A2(new_n281), .A3(new_n192), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n311), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n515), .A2(new_n516), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n741), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT105), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n741), .A2(new_n744), .A3(new_n748), .A4(new_n745), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n691), .A2(new_n710), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n634), .A3(new_n722), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n751), .B1(new_n750), .B2(new_n753), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(G122), .Z(G24));
  NAND3_X1  g571(.A1(new_n741), .A2(new_n744), .A3(new_n674), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n716), .A3(new_n738), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  INV_X1    g575(.A(new_n395), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n385), .B1(new_n720), .B2(new_n383), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n391), .A2(KEYINPUT107), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n389), .A2(new_n765), .A3(new_n390), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n764), .A2(new_n388), .A3(G469), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n762), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n689), .A2(new_n397), .A3(new_n690), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n769), .A2(new_n715), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n745), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n680), .A2(KEYINPUT108), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n321), .B2(new_n745), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n771), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT42), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n769), .A2(new_n770), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n715), .A2(KEYINPUT42), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n728), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n229), .ZN(G33));
  NAND3_X1  g596(.A1(new_n728), .A2(new_n685), .A3(new_n778), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND4_X1  g598(.A1(new_n764), .A2(new_n388), .A3(KEYINPUT45), .A4(new_n766), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n388), .A2(new_n391), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n785), .B(G469), .C1(new_n786), .C2(KEYINPUT45), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT46), .B1(new_n787), .B2(new_n386), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n788), .B1(new_n383), .B2(new_n720), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n386), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n791), .A2(new_n395), .A3(new_n700), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n714), .A2(new_n582), .A3(new_n587), .ZN(new_n793));
  AND2_X1   g607(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n794));
  NOR2_X1   g608(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n793), .B2(new_n795), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n642), .A3(new_n674), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n770), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n792), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  AND2_X1   g617(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n804));
  NOR2_X1   g618(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n791), .B(new_n395), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n321), .A2(new_n519), .A3(new_n715), .A4(new_n770), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n762), .B1(new_n789), .B2(new_n790), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n806), .B(new_n807), .C1(new_n808), .C2(new_n805), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NAND2_X1  g624(.A1(new_n797), .A2(new_n631), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n722), .A3(new_n770), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n759), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n703), .A2(new_n705), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n722), .A2(new_n770), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n519), .A4(new_n631), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n582), .A2(new_n587), .A3(new_n653), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n750), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n811), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n709), .A2(KEYINPUT116), .A3(new_n686), .A4(new_n723), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n709), .A2(new_n686), .A3(new_n723), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n818), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n806), .B1(new_n808), .B2(new_n805), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n721), .A2(new_n384), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(new_n395), .B2(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n819), .A2(new_n811), .A3(new_n770), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n829), .A2(KEYINPUT51), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT51), .B1(new_n829), .B2(new_n834), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n820), .A2(new_n738), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n837), .B(new_n629), .C1(new_n658), .C2(new_n816), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n773), .A2(new_n775), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n812), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n812), .A2(new_n841), .A3(KEYINPUT119), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(KEYINPUT48), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT48), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n842), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n838), .A2(new_n839), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n840), .A2(new_n846), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  OR3_X1    g664(.A1(new_n835), .A2(new_n836), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n588), .A2(new_n714), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT112), .B1(new_n852), .B2(new_n646), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n691), .A2(new_n654), .A3(new_n854), .A4(new_n645), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n644), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n636), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT113), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n859), .A3(new_n636), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n858), .B(new_n860), .C1(new_n754), .C2(new_n755), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n619), .A2(new_n620), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n588), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n644), .A2(new_n647), .A3(new_n863), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n675), .A2(new_n864), .A3(new_n736), .A4(new_n739), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n731), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n693), .A2(new_n695), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n321), .A2(new_n699), .A3(new_n674), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n760), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n691), .A2(new_n768), .A3(new_n684), .A4(new_n710), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n706), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n717), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n871), .A2(new_n874), .A3(KEYINPUT115), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n758), .A2(new_n715), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n681), .A2(new_n696), .B1(new_n738), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n673), .B1(new_n703), .B2(new_n295), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n708), .A2(new_n395), .A3(new_n393), .A4(new_n397), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n715), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n706), .A2(new_n872), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n876), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n868), .B1(new_n875), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n664), .A2(new_n587), .A3(new_n862), .A4(new_n684), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n770), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n321), .A2(new_n699), .A3(new_n674), .A4(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n879), .A2(KEYINPUT114), .A3(new_n699), .A4(new_n886), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n889), .A2(new_n890), .B1(new_n877), .B2(new_n778), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n777), .A2(new_n891), .A3(new_n780), .A4(new_n783), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT115), .B1(new_n871), .B2(new_n874), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n882), .A2(new_n697), .A3(new_n876), .A4(new_n760), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(KEYINPUT52), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n867), .A2(new_n884), .A3(new_n892), .A4(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n777), .A2(new_n891), .A3(new_n780), .A4(new_n783), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n899), .A2(new_n861), .A3(new_n866), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT52), .B1(new_n893), .B2(new_n894), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n868), .B1(new_n878), .B2(new_n882), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT53), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT54), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n896), .A2(new_n897), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n900), .A2(new_n903), .A3(KEYINPUT53), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n851), .A2(new_n910), .B1(G952), .B2(G953), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n831), .B(KEYINPUT49), .Z(new_n912));
  NOR4_X1   g726(.A1(new_n793), .A2(new_n772), .A3(new_n762), .A4(new_n686), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n814), .A3(new_n709), .A4(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT111), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n911), .A2(new_n915), .ZN(G75));
  NAND2_X1  g730(.A1(new_n906), .A2(new_n908), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(G210), .A3(G902), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(KEYINPUT56), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n443), .A2(new_n444), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n440), .ZN(new_n922));
  XOR2_X1   g736(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n918), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n918), .B2(new_n920), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n323), .A2(G952), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(G51));
  XNOR2_X1  g742(.A(new_n385), .B(KEYINPUT57), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n382), .B(KEYINPUT122), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n917), .A2(G902), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n935), .A2(new_n787), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n927), .B1(new_n934), .B2(new_n936), .ZN(G54));
  NAND2_X1  g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n571), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n927), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n935), .A2(new_n571), .A3(new_n938), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(G60));
  XNOR2_X1  g757(.A(new_n650), .B(KEYINPUT59), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n652), .B(new_n944), .C1(new_n930), .C2(new_n931), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n940), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n652), .B1(new_n910), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n917), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n510), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n950), .B1(new_n906), .B2(new_n908), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n927), .B1(new_n955), .B2(new_n672), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n955), .B2(new_n672), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n954), .B(new_n956), .C1(new_n958), .C2(KEYINPUT61), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n900), .A2(new_n903), .A3(KEYINPUT53), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n893), .A2(KEYINPUT52), .A3(new_n894), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(new_n901), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT53), .B1(new_n962), .B2(new_n900), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n672), .B(new_n951), .C1(new_n960), .C2(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n964), .B(new_n940), .C1(new_n510), .C2(new_n955), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT61), .B1(new_n964), .B2(KEYINPUT123), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n959), .A2(new_n967), .ZN(G66));
  OAI21_X1  g782(.A(G953), .B1(new_n424), .B2(new_n633), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n867), .B2(G953), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n921), .B1(G898), .B2(new_n323), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT124), .Z(new_n972));
  XNOR2_X1  g786(.A(new_n970), .B(new_n972), .ZN(G69));
  OR2_X1    g787(.A1(new_n549), .A2(new_n550), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n298), .B(new_n974), .Z(new_n975));
  NOR2_X1   g789(.A1(new_n863), .A2(new_n654), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n701), .A2(new_n976), .A3(new_n770), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n728), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n809), .A2(new_n802), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n878), .A2(new_n717), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  OR3_X1    g795(.A1(new_n712), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n712), .B2(new_n980), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n975), .B1(new_n984), .B2(G953), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n323), .A2(G900), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT126), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  INV_X1    g802(.A(new_n752), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n841), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n808), .A2(new_n700), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n792), .A2(KEYINPUT127), .A3(new_n989), .A4(new_n841), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n783), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n781), .A2(new_n995), .A3(new_n980), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n994), .A2(new_n996), .A3(new_n802), .A4(new_n809), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n987), .B1(new_n997), .B2(new_n323), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n985), .B1(new_n998), .B2(new_n975), .ZN(new_n999));
  OAI21_X1  g813(.A(KEYINPUT125), .B1(new_n998), .B2(new_n975), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n323), .B1(G227), .B2(G900), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n999), .B1(new_n1002), .B2(new_n1000), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(G72));
  NOR2_X1   g819(.A1(new_n292), .A2(new_n192), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n984), .A2(new_n867), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n291), .B2(new_n290), .ZN(new_n1011));
  INV_X1    g825(.A(new_n867), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1009), .B1(new_n997), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n193), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1006), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n898), .A2(new_n904), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1009), .B1(new_n1006), .B2(new_n299), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n940), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1015), .A2(new_n1018), .ZN(G57));
endmodule


