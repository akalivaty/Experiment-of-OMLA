//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n452), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n466), .A2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n466), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n476), .A2(KEYINPUT69), .A3(G124), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n479), .A2(new_n481), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n473), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT3), .B(G2104), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .A3(G138), .A4(new_n473), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT70), .A2(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(G2105), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n490), .A2(G126), .A3(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n489), .A2(new_n491), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n503), .A2(KEYINPUT71), .A3(G62), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n509), .B1(G651), .B2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT72), .B(G51), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n524), .B1(new_n507), .B2(new_n525), .C1(new_n526), .C2(new_n505), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n503), .A2(G63), .ZN(new_n529));
  NAND3_X1  g104(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n527), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n505), .A2(new_n534), .B1(new_n507), .B2(new_n535), .ZN(new_n536));
  XOR2_X1   g111(.A(new_n536), .B(KEYINPUT74), .Z(new_n537));
  AOI22_X1  g112(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT73), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n515), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT75), .B(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n505), .A2(new_n546), .B1(new_n507), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  INV_X1    g130(.A(new_n505), .ZN(new_n556));
  NOR2_X1   g131(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n504), .A2(G53), .A3(G543), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n556), .A2(G91), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n560));
  OR3_X1    g135(.A1(new_n558), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n515), .B2(new_n563), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n564), .A2(KEYINPUT77), .A3(G651), .ZN(new_n565));
  AOI21_X1  g140(.A(KEYINPUT77), .B1(new_n564), .B2(G651), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n559), .B(new_n561), .C1(new_n565), .C2(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(new_n537), .A2(new_n540), .ZN(G301));
  INV_X1    g143(.A(G166), .ZN(G303));
  AOI21_X1  g144(.A(G74), .B1(new_n512), .B2(new_n514), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT78), .B1(new_n570), .B2(new_n528), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n504), .A2(G49), .A3(G543), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n503), .A2(new_n504), .A3(G87), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n574), .B(G651), .C1(new_n503), .C2(G74), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n575), .ZN(G288));
  NAND3_X1  g151(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n504), .A2(new_n579), .A3(G48), .A4(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n515), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n578), .A2(new_n580), .B1(new_n583), .B2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n556), .A2(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n556), .A2(G85), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI221_X1 g164(.A(new_n587), .B1(new_n588), .B2(new_n507), .C1(new_n528), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n556), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(G66), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(G66), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n503), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G79), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n511), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n507), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n504), .A2(KEYINPUT81), .A3(G543), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n604), .A2(G54), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n602), .B1(new_n601), .B2(new_n606), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n594), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n591), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n591), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  XNOR2_X1  g189(.A(G299), .B(KEYINPUT84), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT85), .ZN(G148));
  NAND2_X1  g195(.A1(new_n611), .A2(new_n618), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g199(.A1(G123), .A2(new_n476), .B1(new_n480), .B2(G135), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n473), .A2(G111), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT86), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n634), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2430), .ZN(new_n637));
  INV_X1    g212(.A(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2438), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT87), .B(KEYINPUT16), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2451), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2454), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n644), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n648), .B1(new_n645), .B2(new_n649), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n636), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n636), .B(new_n654), .C1(new_n650), .C2(new_n651), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(G14), .ZN(new_n659));
  INV_X1    g234(.A(new_n652), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n659), .B1(new_n660), .B2(new_n653), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n663), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G2100), .Z(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  AOI21_X1  g246(.A(KEYINPUT18), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n682), .A2(new_n675), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT89), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n682), .A2(new_n675), .A3(new_n678), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n680), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT92), .Z(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT91), .B(G1981), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT90), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n689), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  NAND2_X1  g271(.A1(new_n476), .A2(G129), .ZN(new_n697));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT26), .Z(new_n699));
  AOI22_X1  g274(.A1(new_n490), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n697), .B(new_n699), .C1(G2105), .C2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G29), .B2(G32), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT27), .B(G1996), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT102), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT103), .Z(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NOR2_X1   g288(.A1(G171), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G5), .B2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G1961), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G27), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n719), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT104), .B(G2078), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT105), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n717), .A2(new_n718), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n719), .A2(G26), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n476), .A2(G128), .ZN(new_n727));
  OR2_X1    g302(.A1(G104), .A2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT100), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n473), .ZN(new_n732));
  INV_X1    g307(.A(G140), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n480), .A2(KEYINPUT100), .A3(G140), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n730), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n726), .B1(new_n736), .B2(G29), .ZN(new_n737));
  MUX2_X1   g312(.A(new_n726), .B(new_n737), .S(KEYINPUT28), .Z(new_n738));
  INV_X1    g313(.A(G2067), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n712), .A2(new_n725), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n713), .A2(KEYINPUT23), .A3(G20), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n743));
  INV_X1    g318(.A(G20), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G16), .ZN(new_n745));
  INV_X1    g320(.A(G299), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n742), .B(new_n745), .C1(new_n746), .C2(new_n713), .ZN(new_n747));
  INV_X1    g322(.A(G1956), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n719), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n719), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT29), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT106), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n713), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n611), .B2(new_n713), .ZN(new_n758));
  INV_X1    g333(.A(G1348), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(KEYINPUT24), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(KEYINPUT24), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n719), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G160), .B2(new_n719), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n707), .A2(new_n710), .B1(G2084), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n713), .A2(G21), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G168), .B2(new_n713), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G11), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n480), .A2(G139), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n490), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n773), .B(new_n774), .C1(new_n473), .C2(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G33), .B(new_n776), .S(G29), .Z(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G2072), .Z(new_n778));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G28), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(G28), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n780), .A2(new_n781), .A3(new_n719), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n770), .A2(new_n771), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n766), .B(new_n783), .C1(new_n754), .C2(new_n753), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n741), .A2(new_n756), .A3(new_n760), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n713), .A2(G19), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n549), .B2(new_n713), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1341), .Z(new_n789));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n790));
  NOR2_X1   g365(.A1(G95), .A2(G2105), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n480), .A2(G131), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n476), .A2(G119), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT94), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n719), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n803));
  NOR2_X1   g378(.A1(G25), .A2(G29), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n803), .B1(new_n802), .B2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT35), .B(G1991), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G6), .B(G305), .S(G16), .Z(new_n810));
  XOR2_X1   g385(.A(KEYINPUT32), .B(G1981), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n713), .A2(G22), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G166), .B2(new_n713), .ZN(new_n814));
  INV_X1    g389(.A(G1971), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n713), .A2(G23), .ZN(new_n817));
  INV_X1    g392(.A(G288), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n713), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT33), .B(G1976), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT98), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n812), .A2(new_n816), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT34), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(G16), .A2(G24), .ZN(new_n826));
  XNOR2_X1  g401(.A(G290), .B(KEYINPUT96), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(G16), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT97), .B(G1986), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n809), .A2(new_n825), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n809), .A2(new_n833), .A3(new_n825), .A4(new_n830), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n823), .A2(new_n824), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n790), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g413(.A(KEYINPUT36), .B(new_n836), .C1(new_n832), .C2(new_n834), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n786), .B(new_n789), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n765), .A2(G2084), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n629), .A2(new_n719), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(G311));
  NAND2_X1  g419(.A1(new_n835), .A2(new_n837), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT36), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n835), .A2(new_n790), .A3(new_n837), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n785), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n843), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n848), .A2(new_n841), .A3(new_n849), .A4(new_n789), .ZN(G150));
  AOI22_X1  g425(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n528), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n504), .A2(G55), .A3(G543), .ZN(new_n853));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n505), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n549), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n852), .A2(new_n855), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n545), .B2(new_n548), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n611), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n858), .B1(new_n866), .B2(G860), .ZN(G145));
  NAND2_X1  g442(.A1(new_n476), .A2(G130), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n480), .A2(G142), .ZN(new_n869));
  NOR2_X1   g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n501), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n629), .A2(G160), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n629), .A2(G160), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(G162), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(G162), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n799), .B(new_n632), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n705), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n797), .B(new_n632), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(new_n704), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n877), .B(new_n879), .C1(new_n881), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n705), .A2(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n704), .ZN(new_n886));
  INV_X1    g461(.A(new_n877), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n878), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n736), .B(new_n776), .Z(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n884), .B2(new_n888), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n874), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n884), .A2(new_n888), .ZN(new_n894));
  INV_X1    g469(.A(new_n889), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n873), .A3(new_n890), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g475(.A(new_n621), .B(new_n862), .Z(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n610), .A2(G299), .ZN(new_n903));
  INV_X1    g478(.A(new_n609), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n607), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n746), .B1(new_n905), .B2(new_n594), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n902), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n610), .A2(G299), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n746), .A3(new_n594), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT41), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n901), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n903), .A2(new_n906), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n901), .A2(new_n913), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n911), .A2(new_n914), .A3(KEYINPUT42), .ZN(new_n915));
  AND2_X1   g490(.A1(G290), .A2(G166), .ZN(new_n916));
  NOR2_X1   g491(.A1(G290), .A2(G166), .ZN(new_n917));
  OR3_X1    g492(.A1(new_n916), .A2(new_n917), .A3(new_n818), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n818), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(G305), .B(KEYINPUT107), .Z(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n921), .A3(new_n919), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT42), .B1(new_n911), .B2(new_n914), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n915), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n915), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(G868), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(G868), .B2(new_n860), .ZN(G295));
  OAI21_X1  g506(.A(new_n930), .B1(G868), .B2(new_n860), .ZN(G331));
  NAND3_X1  g507(.A1(new_n859), .A2(G286), .A3(new_n861), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G286), .B1(new_n859), .B2(new_n861), .ZN(new_n935));
  OAI21_X1  g510(.A(G301), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n862), .A2(G168), .ZN(new_n937));
  NAND3_X1  g512(.A1(G171), .A2(new_n937), .A3(new_n933), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n907), .A3(new_n910), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT108), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n939), .A2(new_n907), .A3(new_n942), .A4(new_n910), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n912), .A2(new_n938), .A3(new_n936), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n912), .A2(KEYINPUT109), .A3(new_n938), .A4(new_n936), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n941), .A2(new_n943), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n926), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n925), .A2(new_n940), .A3(new_n944), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n951), .A2(new_n898), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n898), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n925), .B1(new_n940), .B2(new_n944), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n949), .A2(KEYINPUT43), .A3(new_n952), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  MUX2_X1   g535(.A(new_n957), .B(new_n960), .S(KEYINPUT44), .Z(G397));
  INV_X1    g536(.A(G1996), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n704), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n501), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n469), .A2(new_n474), .A3(G40), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G1996), .B1(new_n702), .B2(new_n703), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n963), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n730), .A2(new_n739), .A3(new_n734), .A4(new_n735), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n735), .A2(new_n734), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n727), .A2(new_n729), .ZN(new_n975));
  OAI21_X1  g550(.A(G2067), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n977), .B(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT111), .B1(new_n979), .B2(new_n969), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n977), .A2(new_n978), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT110), .B1(new_n973), .B2(new_n976), .ZN(new_n983));
  OAI211_X1 g558(.A(KEYINPUT111), .B(new_n969), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n972), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n808), .B(KEYINPUT112), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n799), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n799), .A2(new_n986), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n969), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(G290), .B(G1986), .Z(new_n990));
  OAI211_X1 g565(.A(new_n985), .B(new_n989), .C1(new_n970), .C2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT113), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT122), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT45), .B1(new_n501), .B2(new_n964), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n996), .A2(new_n997), .A3(new_n968), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(new_n998), .B2(G1966), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n469), .A2(new_n474), .A3(G40), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n501), .A2(new_n1001), .A3(new_n964), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G2084), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT114), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n1006), .B(new_n1001), .C1(new_n501), .C2(new_n964), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1003), .B(new_n1004), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n967), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(KEYINPUT119), .A3(new_n769), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n999), .A2(G168), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT51), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n999), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(G286), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G303), .A2(G8), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT55), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n965), .A2(KEYINPUT50), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1021), .A2(new_n754), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT118), .B(new_n1022), .C1(new_n998), .C2(G1971), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(G8), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1010), .A2(new_n815), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT118), .B1(new_n1025), .B2(new_n1022), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1020), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n584), .A2(new_n1028), .A3(new_n585), .ZN(new_n1029));
  XOR2_X1   g604(.A(KEYINPUT117), .B(G86), .Z(new_n1030));
  NAND2_X1  g605(.A1(new_n556), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n584), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT49), .B(new_n1029), .C1(new_n1032), .C2(new_n1028), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n584), .A2(new_n1028), .A3(new_n585), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1028), .B1(new_n584), .B2(new_n1031), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  INV_X1    g613(.A(new_n965), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(new_n1000), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1033), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n965), .B2(new_n968), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(G288), .B2(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n571), .A2(new_n575), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n573), .A2(new_n572), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1046), .A2(new_n1048), .A3(KEYINPUT115), .A4(G1976), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1042), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n818), .A2(G1976), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1050), .B(KEYINPUT116), .C1(KEYINPUT52), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1045), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1040), .A2(new_n1053), .A3(new_n1051), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1040), .A2(new_n1053), .A3(KEYINPUT116), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1041), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(new_n1019), .B(KEYINPUT55), .Z(new_n1059));
  OAI21_X1  g634(.A(new_n1003), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1025), .B1(new_n1060), .B2(G2090), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1061), .A3(G8), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1027), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G2078), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n967), .A2(new_n1064), .A3(new_n1000), .A4(new_n1009), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n996), .A2(new_n997), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(KEYINPUT53), .A3(new_n1064), .A4(new_n1000), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1021), .A2(new_n1006), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n965), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1067), .B(new_n1069), .C1(new_n1073), .C2(G1961), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G171), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1060), .A2(new_n716), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1076), .A2(G301), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(KEYINPUT54), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1018), .A2(new_n1063), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(KEYINPUT121), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1074), .A2(new_n1081), .A3(G171), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT54), .B1(new_n1083), .B2(new_n1077), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n994), .B1(new_n1079), .B2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(G299), .B(KEYINPUT57), .Z(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1003), .A2(new_n1021), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n748), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n998), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n965), .A2(new_n968), .A3(KEYINPUT120), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT120), .B1(new_n965), .B2(new_n968), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1096), .A2(new_n739), .B1(new_n1060), .B2(new_n759), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1097), .A2(new_n610), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1086), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT58), .B(G1341), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1010), .A2(G1996), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n549), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT59), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1093), .A2(KEYINPUT61), .A3(new_n1099), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1097), .A2(new_n1111), .A3(new_n611), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1104), .A2(new_n1109), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1097), .A2(new_n610), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1111), .B1(new_n1098), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1093), .B(new_n1101), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1116));
  AND4_X1   g691(.A1(new_n1062), .A2(new_n1078), .A3(new_n1058), .A4(new_n1027), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1074), .A2(new_n1081), .A3(G171), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1081), .B1(new_n1074), .B2(G171), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1077), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1117), .A2(new_n1122), .A3(KEYINPUT122), .A4(new_n1018), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1085), .A2(new_n1116), .A3(new_n1123), .ZN(new_n1124));
  OR3_X1    g699(.A1(new_n1041), .A2(G1976), .A3(G288), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1042), .B1(new_n1125), .B2(new_n1029), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1027), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1016), .A2(G8), .A3(G168), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1129), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1061), .A2(G8), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1127), .B1(new_n1132), .B2(new_n1020), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1131), .A2(new_n1133), .A3(new_n1062), .A4(new_n1058), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1126), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1017), .A2(new_n1013), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1015), .B1(new_n1012), .B2(G8), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT62), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1014), .B(new_n1139), .C1(new_n1013), .C2(new_n1017), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1083), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1138), .A2(new_n1063), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1058), .A2(G8), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1135), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n993), .B1(new_n1124), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n969), .B1(new_n979), .B2(new_n704), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n969), .A2(new_n962), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT46), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1149), .A2(KEYINPUT47), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(KEYINPUT47), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n970), .A2(G1986), .A3(G290), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n1154));
  XOR2_X1   g729(.A(new_n1153), .B(new_n1154), .Z(new_n1155));
  NAND3_X1  g730(.A1(new_n985), .A2(new_n989), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n972), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n808), .B1(new_n798), .B2(new_n801), .ZN(new_n1159));
  INV_X1    g734(.A(new_n984), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1158), .B(new_n1159), .C1(new_n980), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n973), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT123), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1164), .A3(new_n973), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1165), .A3(new_n969), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1163), .A2(new_n1165), .A3(KEYINPUT124), .A4(new_n969), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1152), .B(new_n1157), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1145), .A2(KEYINPUT126), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1135), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1085), .A2(new_n1116), .A3(new_n1123), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n992), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1152), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1161), .A2(new_n1164), .A3(new_n973), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1164), .B1(new_n1161), .B2(new_n973), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT124), .B1(new_n1179), .B2(new_n969), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1169), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1176), .B(new_n1156), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1172), .B1(new_n1175), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1171), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g759(.A(G227), .B1(new_n658), .B2(new_n661), .ZN(new_n1186));
  AND2_X1   g760(.A1(new_n899), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g761(.A1(new_n957), .A2(G319), .A3(new_n695), .A4(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g762(.A(new_n1188), .B(KEYINPUT127), .ZN(G308));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1190));
  XNOR2_X1  g764(.A(new_n1188), .B(new_n1190), .ZN(G225));
endmodule


