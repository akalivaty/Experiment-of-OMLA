

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595;

  NOR2_X1 U320 ( .A1(n476), .A2(n475), .ZN(n477) );
  NAND2_X2 U321 ( .A1(n465), .A2(n464), .ZN(n513) );
  XNOR2_X1 U322 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U323 ( .A(KEYINPUT38), .B(n455), .ZN(n511) );
  NOR2_X1 U324 ( .A1(n482), .A2(n481), .ZN(n288) );
  XNOR2_X1 U325 ( .A(n358), .B(KEYINPUT102), .ZN(n359) );
  XNOR2_X1 U326 ( .A(n360), .B(n359), .ZN(n363) );
  XNOR2_X1 U327 ( .A(n478), .B(KEYINPUT117), .ZN(n479) );
  XNOR2_X1 U328 ( .A(n333), .B(n449), .ZN(n334) );
  XNOR2_X1 U329 ( .A(n480), .B(n479), .ZN(n577) );
  XNOR2_X1 U330 ( .A(n335), .B(n334), .ZN(n339) );
  XNOR2_X1 U331 ( .A(n452), .B(n451), .ZN(n461) );
  INV_X1 U332 ( .A(G43GAT), .ZN(n456) );
  XNOR2_X1 U333 ( .A(n490), .B(G169GAT), .ZN(n491) );
  XNOR2_X1 U334 ( .A(n456), .B(KEYINPUT40), .ZN(n457) );
  XNOR2_X1 U335 ( .A(n492), .B(n491), .ZN(G1348GAT) );
  XNOR2_X1 U336 ( .A(n458), .B(n457), .ZN(G1330GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n290) );
  XNOR2_X1 U338 ( .A(G71GAT), .B(G64GAT), .ZN(n289) );
  XNOR2_X1 U339 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U340 ( .A(KEYINPUT13), .B(G57GAT), .Z(n446) );
  XOR2_X1 U341 ( .A(n291), .B(n446), .Z(n295) );
  XOR2_X1 U342 ( .A(G1GAT), .B(KEYINPUT71), .Z(n293) );
  XNOR2_X1 U343 ( .A(G15GAT), .B(G8GAT), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n424) );
  XOR2_X1 U345 ( .A(G22GAT), .B(G155GAT), .Z(n351) );
  XNOR2_X1 U346 ( .A(n424), .B(n351), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U348 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n297) );
  NAND2_X1 U349 ( .A1(G231GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U351 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U352 ( .A(G211GAT), .B(G78GAT), .Z(n301) );
  XNOR2_X1 U353 ( .A(G183GAT), .B(G127GAT), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n302), .B(KEYINPUT12), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n470) );
  INV_X1 U357 ( .A(n470), .ZN(n589) );
  XOR2_X1 U358 ( .A(KEYINPUT18), .B(KEYINPUT86), .Z(n306) );
  XNOR2_X1 U359 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n308) );
  INV_X1 U361 ( .A(KEYINPUT87), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n310) );
  XNOR2_X1 U363 ( .A(G169GAT), .B(G183GAT), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n329) );
  XOR2_X1 U365 ( .A(G120GAT), .B(G71GAT), .Z(n450) );
  XOR2_X1 U366 ( .A(G127GAT), .B(KEYINPUT0), .Z(n312) );
  XNOR2_X1 U367 ( .A(G113GAT), .B(G134GAT), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n380) );
  XNOR2_X1 U369 ( .A(n450), .B(n380), .ZN(n314) );
  XOR2_X1 U370 ( .A(G43GAT), .B(G99GAT), .Z(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U372 ( .A(KEYINPUT65), .B(KEYINPUT85), .Z(n316) );
  NAND2_X1 U373 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XOR2_X1 U374 ( .A(n316), .B(n315), .Z(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U376 ( .A(KEYINPUT88), .B(G176GAT), .Z(n320) );
  XNOR2_X1 U377 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(n321), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n329), .B(n324), .ZN(n325) );
  INV_X1 U382 ( .A(n325), .ZN(n541) );
  XOR2_X1 U383 ( .A(G92GAT), .B(G204GAT), .Z(n327) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(G218GAT), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n335) );
  XOR2_X1 U387 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n331) );
  NAND2_X1 U388 ( .A1(G226GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n332), .B(KEYINPUT99), .Z(n333) );
  XNOR2_X1 U391 ( .A(G176GAT), .B(G64GAT), .ZN(n449) );
  XOR2_X1 U392 ( .A(G211GAT), .B(KEYINPUT21), .Z(n337) );
  XNOR2_X1 U393 ( .A(G197GAT), .B(KEYINPUT90), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n348) );
  XOR2_X1 U395 ( .A(G36GAT), .B(G190GAT), .Z(n403) );
  XNOR2_X1 U396 ( .A(n348), .B(n403), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n459) );
  NOR2_X1 U398 ( .A1(n541), .A2(n459), .ZN(n357) );
  XOR2_X1 U399 ( .A(G162GAT), .B(KEYINPUT74), .Z(n341) );
  XNOR2_X1 U400 ( .A(G50GAT), .B(G218GAT), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n399) );
  XOR2_X1 U402 ( .A(G78GAT), .B(G204GAT), .Z(n342) );
  XOR2_X1 U403 ( .A(G148GAT), .B(n342), .Z(n442) );
  XOR2_X1 U404 ( .A(n399), .B(n442), .Z(n356) );
  XOR2_X1 U405 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n344) );
  NAND2_X1 U406 ( .A1(G228GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U408 ( .A(n345), .B(KEYINPUT24), .Z(n350) );
  XOR2_X1 U409 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n347) );
  XNOR2_X1 U410 ( .A(G141GAT), .B(KEYINPUT91), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n379) );
  XNOR2_X1 U412 ( .A(n348), .B(n379), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n352) );
  XOR2_X1 U414 ( .A(n352), .B(n351), .Z(n354) );
  XNOR2_X1 U415 ( .A(G106GAT), .B(KEYINPUT22), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n482) );
  NOR2_X1 U418 ( .A1(n357), .A2(n482), .ZN(n360) );
  INV_X1 U419 ( .A(KEYINPUT25), .ZN(n358) );
  NAND2_X1 U420 ( .A1(n482), .A2(n541), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n361), .B(KEYINPUT26), .ZN(n579) );
  XNOR2_X1 U422 ( .A(n459), .B(KEYINPUT27), .ZN(n388) );
  NOR2_X1 U423 ( .A1(n579), .A2(n388), .ZN(n362) );
  NOR2_X1 U424 ( .A1(n363), .A2(n362), .ZN(n364) );
  XNOR2_X1 U425 ( .A(KEYINPUT103), .B(n364), .ZN(n387) );
  NAND2_X1 U426 ( .A1(G225GAT), .A2(G233GAT), .ZN(n370) );
  XOR2_X1 U427 ( .A(G155GAT), .B(G148GAT), .Z(n366) );
  XNOR2_X1 U428 ( .A(G120GAT), .B(G162GAT), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U430 ( .A(G29GAT), .B(G85GAT), .Z(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n386) );
  XOR2_X1 U433 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n372) );
  XNOR2_X1 U434 ( .A(KEYINPUT1), .B(KEYINPUT93), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n384) );
  XOR2_X1 U436 ( .A(KEYINPUT97), .B(KEYINPUT92), .Z(n374) );
  XNOR2_X1 U437 ( .A(G1GAT), .B(G57GAT), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U439 ( .A(KEYINPUT96), .B(KEYINPUT4), .Z(n376) );
  XNOR2_X1 U440 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U442 ( .A(n378), .B(n377), .Z(n382) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U445 ( .A(n384), .B(n383), .Z(n385) );
  XNOR2_X1 U446 ( .A(n386), .B(n385), .ZN(n576) );
  NAND2_X1 U447 ( .A1(n387), .A2(n576), .ZN(n392) );
  NOR2_X1 U448 ( .A1(n576), .A2(n388), .ZN(n536) );
  XOR2_X1 U449 ( .A(KEYINPUT28), .B(n482), .Z(n539) );
  NAND2_X1 U450 ( .A1(n536), .A2(n539), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n389), .B(KEYINPUT101), .ZN(n390) );
  NAND2_X1 U452 ( .A1(n390), .A2(n541), .ZN(n391) );
  NAND2_X1 U453 ( .A1(n392), .A2(n391), .ZN(n393) );
  XOR2_X1 U454 ( .A(n393), .B(KEYINPUT104), .Z(n497) );
  NOR2_X1 U455 ( .A1(n589), .A2(n497), .ZN(n394) );
  XNOR2_X1 U456 ( .A(n394), .B(KEYINPUT107), .ZN(n420) );
  INV_X1 U457 ( .A(KEYINPUT80), .ZN(n419) );
  XOR2_X1 U458 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n396) );
  XNOR2_X1 U459 ( .A(KEYINPUT67), .B(KEYINPUT11), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n418) );
  XOR2_X1 U461 ( .A(G85GAT), .B(G92GAT), .Z(n398) );
  XNOR2_X1 U462 ( .A(G99GAT), .B(G106GAT), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n441) );
  XNOR2_X1 U464 ( .A(n399), .B(n441), .ZN(n416) );
  XOR2_X1 U465 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n401) );
  XNOR2_X1 U466 ( .A(G134GAT), .B(KEYINPUT76), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n404) );
  INV_X1 U468 ( .A(n404), .ZN(n402) );
  NAND2_X1 U469 ( .A1(n403), .A2(n402), .ZN(n407) );
  INV_X1 U470 ( .A(n403), .ZN(n405) );
  NAND2_X1 U471 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X1 U472 ( .A1(n407), .A2(n406), .ZN(n409) );
  NAND2_X1 U473 ( .A1(G232GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n410), .B(KEYINPUT75), .ZN(n414) );
  XOR2_X1 U476 ( .A(G29GAT), .B(G43GAT), .Z(n412) );
  XNOR2_X1 U477 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n412), .B(n411), .ZN(n435) );
  XOR2_X1 U479 ( .A(n435), .B(KEYINPUT78), .Z(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n561) );
  XNOR2_X1 U483 ( .A(n419), .B(n561), .ZN(n549) );
  XNOR2_X1 U484 ( .A(KEYINPUT36), .B(n549), .ZN(n592) );
  NOR2_X1 U485 ( .A1(n420), .A2(n592), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n421), .B(KEYINPUT37), .ZN(n526) );
  XOR2_X1 U487 ( .A(G36GAT), .B(G50GAT), .Z(n423) );
  NAND2_X1 U488 ( .A1(G229GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U489 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U490 ( .A(n425), .B(n424), .Z(n433) );
  XOR2_X1 U491 ( .A(G141GAT), .B(G197GAT), .Z(n427) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(G22GAT), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U494 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n429) );
  XNOR2_X1 U495 ( .A(G113GAT), .B(KEYINPUT70), .ZN(n428) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U499 ( .A(n434), .B(KEYINPUT29), .Z(n437) );
  XNOR2_X1 U500 ( .A(n435), .B(KEYINPUT30), .ZN(n436) );
  XNOR2_X1 U501 ( .A(n437), .B(n436), .ZN(n580) );
  XOR2_X1 U502 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n439) );
  NAND2_X1 U503 ( .A1(G230GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U504 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U505 ( .A(n440), .B(KEYINPUT73), .Z(n444) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U507 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U508 ( .A(n445), .B(KEYINPUT72), .Z(n448) );
  XNOR2_X1 U509 ( .A(n446), .B(KEYINPUT33), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n452) );
  NAND2_X1 U511 ( .A1(n580), .A2(n461), .ZN(n499) );
  NOR2_X1 U512 ( .A1(n526), .A2(n499), .ZN(n454) );
  INV_X1 U513 ( .A(KEYINPUT108), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  NOR2_X1 U515 ( .A1(n511), .A2(n541), .ZN(n458) );
  XNOR2_X1 U516 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n461), .A2(n460), .ZN(n465) );
  INV_X1 U518 ( .A(n460), .ZN(n463) );
  INV_X1 U519 ( .A(n461), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U521 ( .A1(n580), .A2(n513), .ZN(n466) );
  XOR2_X1 U522 ( .A(KEYINPUT46), .B(n466), .Z(n467) );
  NOR2_X1 U523 ( .A1(n561), .A2(n467), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n470), .A2(n468), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT47), .ZN(n476) );
  NOR2_X1 U526 ( .A1(n592), .A2(n470), .ZN(n472) );
  XNOR2_X1 U527 ( .A(KEYINPUT45), .B(KEYINPUT66), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n473), .A2(n461), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n474), .A2(n580), .ZN(n475) );
  XNOR2_X1 U531 ( .A(KEYINPUT48), .B(n477), .ZN(n535) );
  NOR2_X1 U532 ( .A1(n459), .A2(n535), .ZN(n480) );
  INV_X1 U533 ( .A(KEYINPUT54), .ZN(n478) );
  INV_X1 U534 ( .A(n576), .ZN(n481) );
  AND2_X1 U535 ( .A1(n577), .A2(n288), .ZN(n483) );
  XNOR2_X1 U536 ( .A(n483), .B(KEYINPUT55), .ZN(n485) );
  NOR2_X1 U537 ( .A1(n541), .A2(n485), .ZN(n484) );
  NAND2_X1 U538 ( .A1(KEYINPUT118), .A2(n484), .ZN(n489) );
  INV_X1 U539 ( .A(KEYINPUT118), .ZN(n487) );
  OR2_X1 U540 ( .A1(n541), .A2(n485), .ZN(n486) );
  NAND2_X1 U541 ( .A1(n487), .A2(n486), .ZN(n488) );
  NAND2_X1 U542 ( .A1(n489), .A2(n488), .ZN(n571) );
  NAND2_X1 U543 ( .A1(n580), .A2(n571), .ZN(n492) );
  XOR2_X1 U544 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n490) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n494) );
  NAND2_X1 U546 ( .A1(n589), .A2(n549), .ZN(n493) );
  XNOR2_X1 U547 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U548 ( .A(n495), .B(KEYINPUT83), .ZN(n496) );
  NOR2_X1 U549 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U550 ( .A(KEYINPUT105), .B(n498), .ZN(n515) );
  OR2_X1 U551 ( .A1(n499), .A2(n515), .ZN(n506) );
  NOR2_X1 U552 ( .A1(n576), .A2(n506), .ZN(n501) );
  XNOR2_X1 U553 ( .A(KEYINPUT34), .B(KEYINPUT106), .ZN(n500) );
  XNOR2_X1 U554 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U555 ( .A(G1GAT), .B(n502), .Z(G1324GAT) );
  NOR2_X1 U556 ( .A1(n459), .A2(n506), .ZN(n503) );
  XOR2_X1 U557 ( .A(G8GAT), .B(n503), .Z(G1325GAT) );
  NOR2_X1 U558 ( .A1(n541), .A2(n506), .ZN(n505) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n504) );
  XNOR2_X1 U560 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NOR2_X1 U561 ( .A1(n539), .A2(n506), .ZN(n507) );
  XOR2_X1 U562 ( .A(G22GAT), .B(n507), .Z(G1327GAT) );
  NOR2_X1 U563 ( .A1(n511), .A2(n576), .ZN(n509) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n508) );
  XNOR2_X1 U565 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  NOR2_X1 U566 ( .A1(n511), .A2(n459), .ZN(n510) );
  XOR2_X1 U567 ( .A(G36GAT), .B(n510), .Z(G1329GAT) );
  NOR2_X1 U568 ( .A1(n539), .A2(n511), .ZN(n512) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  INV_X1 U570 ( .A(n580), .ZN(n514) );
  NAND2_X1 U571 ( .A1(n514), .A2(n513), .ZN(n525) );
  OR2_X1 U572 ( .A1(n525), .A2(n515), .ZN(n522) );
  NOR2_X1 U573 ( .A1(n576), .A2(n522), .ZN(n517) );
  XNOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n516) );
  XNOR2_X1 U575 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n518), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n459), .A2(n522), .ZN(n519) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n519), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n541), .A2(n522), .ZN(n520) );
  XOR2_X1 U580 ( .A(KEYINPUT110), .B(n520), .Z(n521) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(n521), .ZN(G1334GAT) );
  NOR2_X1 U582 ( .A1(n539), .A2(n522), .ZN(n524) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n523) );
  XNOR2_X1 U584 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  OR2_X1 U585 ( .A1(n526), .A2(n525), .ZN(n531) );
  NOR2_X1 U586 ( .A1(n576), .A2(n531), .ZN(n528) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n527) );
  XNOR2_X1 U588 ( .A(n528), .B(n527), .ZN(G1336GAT) );
  NOR2_X1 U589 ( .A1(n459), .A2(n531), .ZN(n529) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n529), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n541), .A2(n531), .ZN(n530) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n539), .A2(n531), .ZN(n533) );
  XNOR2_X1 U594 ( .A(KEYINPUT112), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U596 ( .A(G106GAT), .B(n534), .Z(G1339GAT) );
  XOR2_X1 U597 ( .A(G113GAT), .B(KEYINPUT115), .Z(n544) );
  INV_X1 U598 ( .A(n535), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U600 ( .A(KEYINPUT113), .B(n538), .ZN(n553) );
  NAND2_X1 U601 ( .A1(n553), .A2(n539), .ZN(n540) );
  NOR2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT114), .B(n542), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n580), .A2(n550), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n544), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U607 ( .A1(n550), .A2(n513), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U609 ( .A1(n550), .A2(n589), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  INV_X1 U613 ( .A(n549), .ZN(n570) );
  NAND2_X1 U614 ( .A1(n570), .A2(n550), .ZN(n551) );
  XNOR2_X1 U615 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  INV_X1 U616 ( .A(n579), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT116), .B(n555), .Z(n562) );
  NAND2_X1 U619 ( .A1(n562), .A2(n580), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n556), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n558) );
  NAND2_X1 U622 ( .A1(n562), .A2(n513), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n562), .A2(n589), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U630 ( .A1(n571), .A2(n513), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT56), .Z(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n571), .A2(n589), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT122), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G183GAT), .B(n569), .ZN(G1350GAT) );
  AND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n575) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT123), .ZN(n573) );
  XNOR2_X1 U640 ( .A(KEYINPUT58), .B(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1351GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n588) );
  NAND2_X1 U645 ( .A1(n588), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  INV_X1 U648 ( .A(n588), .ZN(n591) );
  NOR2_X1 U649 ( .A1(n591), .A2(n461), .ZN(n587) );
  XOR2_X1 U650 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n585) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n594) );
  XNOR2_X1 U657 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

