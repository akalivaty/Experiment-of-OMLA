//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND3_X1   g035(.A1(new_n460), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(KEYINPUT66), .B1(new_n460), .B2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G101), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G137), .A3(new_n460), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n460), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n460), .B1(new_n473), .B2(new_n474), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n481), .B(new_n482), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n477), .B(new_n480), .C1(new_n483), .C2(G124), .ZN(G162));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n486), .B1(new_n467), .B2(new_n468), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT68), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n464), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n487), .A2(KEYINPUT68), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(G126), .B2(new_n481), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n491), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n505), .A2(G651), .B1(G50), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n502), .A2(new_n501), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT69), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n507), .A2(new_n508), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  XOR2_X1   g093(.A(KEYINPUT70), .B(G88), .Z(new_n519));
  NAND3_X1  g094(.A1(new_n514), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n510), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT71), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n510), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n509), .A2(G51), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n528));
  AND3_X1   g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n526), .B(new_n527), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n514), .A2(new_n518), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(G89), .B2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n514), .A2(G90), .A3(new_n518), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n509), .A2(G52), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n538), .A2(KEYINPUT73), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT73), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n533), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n503), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G651), .B1(G43), .B2(new_n509), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  OAI211_X1 g130(.A(G53), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n515), .A2(new_n558), .A3(G53), .A4(G543), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT74), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT74), .B1(new_n557), .B2(new_n559), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n514), .A2(G91), .A3(new_n518), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n503), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT75), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n558), .B1(new_n509), .B2(G53), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n575), .A2(new_n576), .A3(new_n567), .A4(new_n563), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n569), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  INV_X1    g155(.A(new_n524), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n523), .B1(new_n510), .B2(new_n520), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n522), .A2(KEYINPUT76), .A3(new_n524), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G303));
  NAND2_X1  g160(.A1(new_n533), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n509), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(G288));
  NAND3_X1  g166(.A1(new_n514), .A2(G86), .A3(new_n518), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n509), .A2(G48), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  OAI21_X1  g169(.A(G61), .B1(new_n501), .B2(new_n502), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n594), .B1(new_n597), .B2(G651), .ZN(new_n598));
  AOI211_X1 g173(.A(KEYINPUT78), .B(new_n536), .C1(new_n595), .C2(new_n596), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n592), .B(new_n593), .C1(new_n598), .C2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n509), .A2(G47), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n514), .A2(new_n518), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI221_X1 g179(.A(new_n601), .B1(new_n536), .B2(new_n602), .C1(new_n603), .C2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(new_n536), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n509), .A2(G54), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n603), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n610), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G284));
  OAI21_X1  g191(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  MUX2_X1   g193(.A(G286), .B(G299), .S(new_n618), .Z(G280));
  XOR2_X1   g194(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g195(.A(new_n615), .ZN(new_n621));
  INV_X1    g196(.A(G860), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(G559), .B2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT80), .Z(G148));
  NAND2_X1  g199(.A1(new_n549), .A2(new_n618), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n621), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n475), .A2(G135), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n460), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n481), .B(KEYINPUT67), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n629), .B1(new_n630), .B2(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT82), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n461), .A2(new_n462), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(new_n464), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(G2100), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n637), .A2(new_n638), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT17), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n668), .B2(new_n666), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(new_n666), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT18), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n668), .A2(new_n671), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n677), .B1(new_n667), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT87), .B(G2096), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n688), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n693), .B(new_n695), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT20), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT89), .ZN(new_n700));
  XOR2_X1   g275(.A(G1981), .B(G1986), .Z(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n700), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NOR2_X1   g283(.A1(G166), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n708), .B2(G22), .ZN(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G16), .A2(G23), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT92), .Z(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G288), .B2(new_n708), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT33), .B(G1976), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n708), .A2(G6), .ZN(new_n719));
  INV_X1    g294(.A(G305), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n708), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT32), .B(G1981), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT91), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n710), .B2(new_n711), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G24), .B(G290), .S(G16), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n483), .A2(G119), .ZN(new_n733));
  NOR2_X1   g308(.A1(G95), .A2(G2105), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT90), .Z(new_n735));
  INV_X1    g310(.A(G2104), .ZN(new_n736));
  INV_X1    g311(.A(G107), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n735), .A2(new_n738), .B1(G131), .B2(new_n475), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n732), .B1(new_n741), .B2(new_n731), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n742), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n730), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n728), .A2(KEYINPUT36), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n726), .B(KEYINPUT34), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(new_n746), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n635), .A2(G29), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT98), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(G28), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n731), .B1(new_n755), .B2(G28), .ZN(new_n757));
  AND2_X1   g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  NOR2_X1   g333(.A1(KEYINPUT31), .A2(G11), .ZN(new_n759));
  OAI22_X1  g334(.A1(new_n756), .A2(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n731), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT28), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n475), .A2(G140), .ZN(new_n763));
  NOR2_X1   g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(new_n460), .B2(G116), .ZN(new_n766));
  INV_X1    g341(.A(G128), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n763), .B1(new_n765), .B2(new_n766), .C1(new_n632), .C2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n760), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  INV_X1    g347(.A(G1341), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n708), .A2(G19), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT93), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n549), .B2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n772), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n731), .A2(G33), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(new_n460), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n475), .A2(G139), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT25), .Z(new_n783));
  NAND3_X1  g358(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT95), .Z(new_n785));
  OAI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(new_n731), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G2072), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n754), .A2(new_n771), .A3(new_n777), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n731), .A2(G35), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G162), .B2(new_n731), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT29), .ZN(new_n791));
  INV_X1    g366(.A(G2090), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(KEYINPUT29), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n731), .A2(G32), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n483), .A2(G129), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n640), .A2(G105), .ZN(new_n797));
  NAND3_X1  g372(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT26), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n475), .A2(G141), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n796), .A2(new_n797), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT27), .B(G1996), .ZN(new_n803));
  NOR2_X1   g378(.A1(G27), .A2(G29), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G164), .B2(G29), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n802), .A2(new_n803), .B1(G2078), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n776), .ZN(new_n807));
  INV_X1    g382(.A(new_n805), .ZN(new_n808));
  INV_X1    g383(.A(G2078), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n807), .A2(G1341), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n794), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n788), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n753), .A2(KEYINPUT98), .ZN(new_n813));
  INV_X1    g388(.A(G34), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT24), .ZN(new_n815));
  AOI21_X1  g390(.A(G29), .B1(new_n814), .B2(KEYINPUT24), .ZN(new_n816));
  AOI22_X1  g391(.A1(G160), .A2(G29), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G2084), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT96), .Z(new_n819));
  OAI211_X1 g394(.A(new_n813), .B(new_n819), .C1(G2072), .C2(new_n786), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n708), .A2(G5), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G171), .B2(new_n708), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n820), .B1(G1961), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(G168), .A2(G16), .ZN(new_n824));
  NOR2_X1   g399(.A1(G16), .A2(G21), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(KEYINPUT97), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(KEYINPUT97), .B2(new_n824), .ZN(new_n827));
  INV_X1    g402(.A(G1966), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n792), .B1(new_n791), .B2(new_n793), .ZN(new_n830));
  NOR2_X1   g405(.A1(G4), .A2(G16), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n615), .B2(G16), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(G1348), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(G1348), .ZN(new_n834));
  NOR4_X1   g409(.A1(new_n829), .A2(new_n830), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n812), .A2(new_n823), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n817), .A2(G2084), .ZN(new_n837));
  OAI221_X1 g412(.A(new_n837), .B1(new_n802), .B2(new_n803), .C1(new_n822), .C2(G1961), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT99), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n708), .A2(G20), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT23), .Z(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G299), .B2(G16), .ZN(new_n842));
  INV_X1    g417(.A(G1956), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n836), .A2(new_n839), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT100), .B1(new_n752), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g421(.A(KEYINPUT100), .B(new_n845), .C1(new_n748), .C2(new_n751), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(G311));
  NAND2_X1  g424(.A1(new_n752), .A2(new_n845), .ZN(G150));
  NAND2_X1  g425(.A1(new_n615), .A2(G559), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT38), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n509), .A2(G55), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G93), .ZN(new_n855));
  OAI221_X1 g430(.A(new_n853), .B1(new_n536), .B2(new_n854), .C1(new_n603), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n549), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n852), .B(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n622), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n853), .B1(new_n854), .B2(new_n536), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n533), .B2(G93), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n622), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(new_n768), .B(new_n498), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n475), .A2(G142), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n460), .A2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  INV_X1    g445(.A(G130), .ZN(new_n871));
  OAI221_X1 g446(.A(new_n868), .B1(new_n869), .B2(new_n870), .C1(new_n632), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n785), .B(new_n801), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n740), .B(KEYINPUT101), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(new_n642), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n876), .A2(new_n642), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n877), .ZN(new_n880));
  INV_X1    g455(.A(new_n801), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n785), .B(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n874), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n882), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n873), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G160), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n635), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G162), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n887), .A3(new_n884), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(new_n856), .A2(new_n618), .ZN(new_n898));
  XOR2_X1   g473(.A(G166), .B(G290), .Z(new_n899));
  XNOR2_X1  g474(.A(G288), .B(new_n720), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT42), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(KEYINPUT104), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n569), .A2(new_n615), .A3(new_n577), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n615), .B1(new_n569), .B2(new_n577), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT41), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(G299), .A2(new_n621), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n906), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n912), .A3(KEYINPUT103), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n626), .B(new_n857), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n906), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT41), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n914), .A2(new_n915), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n920), .B(KEYINPUT102), .Z(new_n921));
  OAI21_X1  g496(.A(new_n905), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n919), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(KEYINPUT104), .B2(new_n904), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n922), .A2(new_n924), .B1(KEYINPUT104), .B2(new_n904), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n898), .B1(new_n925), .B2(new_n618), .ZN(G295));
  OAI21_X1  g501(.A(new_n898), .B1(new_n925), .B2(new_n618), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n909), .A2(new_n912), .ZN(new_n929));
  NAND2_X1  g504(.A1(G301), .A2(G286), .ZN(new_n930));
  OAI211_X1 g505(.A(G168), .B(new_n537), .C1(new_n540), .C2(new_n541), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n857), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n549), .B(new_n863), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(new_n930), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n933), .B2(new_n935), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n932), .A2(new_n857), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(KEYINPUT105), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n937), .B1(new_n942), .B2(new_n915), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n943), .B2(new_n903), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n917), .B(new_n913), .C1(new_n939), .C2(new_n941), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n901), .A2(new_n902), .ZN(new_n946));
  INV_X1    g521(.A(new_n915), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n933), .A2(new_n947), .A3(new_n935), .A4(KEYINPUT106), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n936), .B2(new_n915), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n945), .A2(new_n946), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n945), .A2(new_n948), .A3(new_n950), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n956), .B2(new_n903), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n928), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n903), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n895), .A3(new_n951), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n961), .A2(KEYINPUT43), .B1(new_n955), .B2(new_n944), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n928), .B2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n481), .A2(G126), .ZN(new_n966));
  INV_X1    g541(.A(new_n496), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n493), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n471), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(G40), .A3(new_n463), .A4(new_n465), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n768), .B(G2067), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n975), .B2(new_n801), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT125), .Z(new_n977));
  NOR3_X1   g552(.A1(new_n971), .A2(G1996), .A3(new_n973), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT46), .Z(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n801), .B(G1996), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n982), .A2(new_n975), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n740), .B(new_n744), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n974), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n974), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT48), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n987), .A2(KEYINPUT48), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n741), .A2(new_n743), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n983), .A2(new_n991), .B1(G2067), .B2(new_n768), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n974), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n981), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1976), .ZN(new_n995));
  OR2_X1    g570(.A1(G288), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G40), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n466), .A2(new_n997), .A3(new_n471), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n998), .A2(new_n498), .A3(new_n964), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT110), .B(G8), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT52), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n995), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n996), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G305), .B2(G1981), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n592), .A2(new_n593), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT78), .B1(new_n1013), .B2(new_n536), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n597), .A2(new_n594), .A3(G651), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1011), .A2(KEYINPUT111), .A3(new_n1012), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G305), .A2(G1981), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT112), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1010), .A2(new_n1017), .B1(G1981), .B2(G305), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1002), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1008), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n971), .A2(new_n998), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n711), .ZN(new_n1033));
  NOR2_X1   g608(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n973), .B1(new_n498), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT108), .B(G2090), .Z(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1030), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(G303), .B2(G8), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1040), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1030), .B(new_n1042), .C1(new_n583), .C2(new_n584), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT49), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1024), .B1(new_n1023), .B2(KEYINPUT49), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1027), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G288), .A2(G1976), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1047), .A2(new_n1048), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1029), .A2(new_n1044), .B1(new_n1049), .B2(new_n1002), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1042), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1038), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n973), .B1(new_n969), .B2(new_n970), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1971), .B1(new_n1054), .B2(new_n1031), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1001), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(G303), .A2(G8), .A3(new_n1040), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1047), .A2(new_n1058), .A3(new_n1044), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT124), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(G2084), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1966), .B1(new_n1054), .B2(new_n1031), .ZN(new_n1065));
  OAI211_X1 g640(.A(G286), .B(new_n1001), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1032), .A2(new_n828), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1034), .B1(new_n965), .B2(new_n968), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n998), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n498), .B2(new_n964), .ZN(new_n1071));
  OR3_X1    g646(.A1(new_n1069), .A2(new_n1071), .A3(G2084), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1030), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G168), .A2(new_n1000), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1066), .B(KEYINPUT51), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1001), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1078), .A3(KEYINPUT62), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1961), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1032), .A2(G2078), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(KEYINPUT53), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1032), .B2(G2078), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1079), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT62), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1050), .B1(new_n1062), .B2(new_n1090), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  NOR4_X1   g668(.A1(new_n1092), .A2(new_n1093), .A3(G286), .A4(new_n1076), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(new_n1044), .A3(new_n1028), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1076), .A2(G286), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1028), .A2(new_n1058), .A3(new_n1044), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1093), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1060), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT113), .B1(new_n1100), .B2(new_n1096), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1095), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1091), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1082), .A2(G301), .A3(new_n1084), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1086), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT54), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1086), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1100), .A2(new_n1061), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1060), .A2(KEYINPUT124), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n843), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n971), .A2(new_n998), .A3(new_n1031), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n568), .A2(KEYINPUT114), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n557), .A2(new_n559), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n563), .A2(new_n1122), .A3(new_n567), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n563), .A2(KEYINPUT57), .A3(new_n567), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT115), .B1(new_n562), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n563), .A2(KEYINPUT57), .A3(new_n567), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n575), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1119), .A2(new_n1124), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT116), .B1(new_n1118), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1124), .A2(new_n1119), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT116), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1118), .A2(new_n1130), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1118), .A2(new_n1130), .A3(KEYINPUT120), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1114), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n615), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n968), .ZN(new_n1149));
  AOI21_X1  g724(.A(G1384), .B1(new_n1149), .B2(new_n491), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n998), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n999), .A2(KEYINPUT117), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n770), .ZN(new_n1155));
  AOI21_X1  g730(.A(G1348), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT118), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(G2067), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT118), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n1156), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1148), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n615), .A2(new_n1147), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g739(.A(new_n1148), .B1(new_n1147), .B2(new_n615), .C1(new_n1158), .C2(new_n1161), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1161), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1160), .B1(new_n1159), .B2(new_n1156), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(new_n1167), .A3(new_n1146), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1164), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT58), .B(G1341), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1154), .A2(new_n1170), .B1(new_n1032), .B2(G1996), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1171), .A2(KEYINPUT119), .A3(new_n550), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1171), .A2(KEYINPUT119), .A3(new_n1174), .A4(new_n550), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1134), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1114), .B1(new_n1118), .B2(new_n1130), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1173), .A2(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g753(.A(KEYINPUT121), .B(new_n1114), .C1(new_n1137), .C2(new_n1142), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1145), .A2(new_n1169), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1166), .A2(new_n615), .A3(new_n1167), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1181), .A2(new_n1138), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n1182), .A2(new_n1137), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1113), .B1(new_n1184), .B2(KEYINPUT123), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1180), .A2(new_n1186), .A3(new_n1183), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1103), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  AND2_X1   g763(.A1(G290), .A2(G1986), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT107), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1189), .A2(new_n986), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(G290), .A2(new_n1190), .A3(G1986), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n974), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n985), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n994), .B1(new_n1188), .B2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g770(.A1(new_n684), .A2(new_n706), .A3(new_n664), .A4(G319), .ZN(new_n1197));
  INV_X1    g771(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n896), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g773(.A(KEYINPUT126), .B1(new_n962), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g774(.A(G37), .B1(new_n888), .B2(new_n891), .ZN(new_n1201));
  AOI21_X1  g775(.A(new_n1197), .B1(new_n1201), .B2(new_n894), .ZN(new_n1202));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n1203));
  AND2_X1   g777(.A1(new_n955), .A2(new_n944), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n954), .B1(new_n957), .B2(new_n951), .ZN(new_n1205));
  OAI211_X1 g779(.A(new_n1202), .B(new_n1203), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  AND2_X1   g780(.A1(new_n1200), .A2(new_n1206), .ZN(G308));
  OAI21_X1  g781(.A(new_n1202), .B1(new_n1204), .B2(new_n1205), .ZN(G225));
endmodule


