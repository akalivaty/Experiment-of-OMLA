//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G22gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT22), .ZN(new_n211));
  INV_X1    g010(.A(G211gat), .ZN(new_n212));
  INV_X1    g011(.A(G218gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT29), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G211gat), .A2(G218gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n213), .ZN(new_n220));
  AND2_X1   g019(.A1(G197gat), .A2(G204gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G197gat), .A2(G204gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n219), .B(new_n220), .C1(new_n223), .C2(new_n211), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(new_n214), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT78), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT3), .B1(new_n218), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G141gat), .B(G148gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n232), .B1(G155gat), .B2(G162gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G141gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G148gat), .ZN(new_n236));
  INV_X1    g035(.A(G148gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G141gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G155gat), .B(G162gat), .ZN(new_n240));
  INV_X1    g039(.A(G155gat), .ZN(new_n241));
  INV_X1    g040(.A(G162gat), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT2), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n234), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT79), .B1(new_n227), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT78), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(new_n217), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT79), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n244), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n244), .A3(new_n247), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n216), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n224), .A2(new_n225), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n246), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G228gat), .A2(G233gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT80), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n261), .A3(new_n258), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n254), .B2(new_n255), .ZN(new_n264));
  INV_X1    g063(.A(new_n255), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT3), .B1(new_n265), .B2(new_n216), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n266), .B2(new_n245), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n207), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n206), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n257), .A2(new_n261), .A3(new_n258), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n261), .B1(new_n257), .B2(new_n258), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n267), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(new_n269), .A3(G22gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n207), .B(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT82), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n263), .A2(new_n277), .A3(new_n207), .A4(new_n267), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n270), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n275), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n205), .B1(new_n268), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G15gat), .B(G43gat), .Z(new_n283));
  XNOR2_X1  g082(.A(G71gat), .B(G99gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT64), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT26), .ZN(new_n294));
  AOI211_X1 g093(.A(new_n290), .B(new_n294), .C1(KEYINPUT26), .C2(new_n293), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G183gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT69), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT27), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT69), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n296), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306));
  AOI21_X1  g105(.A(G190gat), .B1(new_n298), .B2(KEYINPUT69), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT27), .B(G183gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n307), .B(KEYINPUT70), .C1(KEYINPUT69), .C2(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n308), .A2(KEYINPUT28), .A3(new_n300), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n295), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313));
  AND2_X1   g112(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n289), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n293), .B1(KEYINPUT23), .B2(new_n291), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(new_n293), .B2(KEYINPUT23), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n289), .A2(KEYINPUT65), .A3(new_n316), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n319), .B1(new_n327), .B2(new_n315), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G169gat), .ZN(new_n330));
  OR2_X1    g129(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(KEYINPUT67), .A3(new_n330), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT25), .B1(new_n328), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n323), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI211_X1 g142(.A(KEYINPUT68), .B(KEYINPUT25), .C1(new_n328), .C2(new_n340), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n312), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G134gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G127gat), .ZN(new_n347));
  INV_X1    g146(.A(G127gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G134gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G113gat), .B(G120gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(KEYINPUT1), .ZN(new_n352));
  INV_X1    g151(.A(G120gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G113gat), .ZN(new_n354));
  INV_X1    g153(.A(G113gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G120gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n352), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n326), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT65), .B1(new_n289), .B2(new_n316), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n315), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT67), .B1(new_n338), .B2(new_n330), .ZN(new_n366));
  AND4_X1   g165(.A1(KEYINPUT67), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n365), .B(new_n320), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n321), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT68), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n341), .A2(new_n342), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(new_n323), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n352), .A2(new_n360), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n312), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n288), .B1(new_n362), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n285), .B1(new_n375), .B2(KEYINPUT33), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n374), .ZN(new_n380));
  AOI221_X4 g179(.A(new_n377), .B1(KEYINPUT33), .B2(new_n285), .C1(new_n380), .C2(new_n287), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT34), .ZN(new_n382));
  INV_X1    g181(.A(new_n286), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n383), .B1(new_n380), .B2(KEYINPUT71), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT71), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n362), .A2(new_n385), .A3(new_n374), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n380), .A2(KEYINPUT34), .A3(new_n287), .ZN(new_n388));
  OAI22_X1  g187(.A1(new_n379), .A2(new_n381), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT72), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n345), .A2(new_n361), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n373), .B1(new_n372), .B2(new_n312), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n287), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT32), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n396), .A3(new_n285), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT71), .B1(new_n391), .B2(new_n392), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(new_n286), .A3(new_n386), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT34), .ZN(new_n400));
  INV_X1    g199(.A(new_n285), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n393), .B(KEYINPUT32), .C1(new_n395), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n388), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n397), .A2(new_n400), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n390), .A3(new_n404), .ZN(new_n405));
  OAI221_X1 g204(.A(KEYINPUT72), .B1(new_n387), .B2(new_n388), .C1(new_n379), .C2(new_n381), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n280), .A2(new_n282), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(new_n253), .A3(new_n361), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n234), .A2(new_n352), .A3(new_n244), .A4(new_n360), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT75), .B1(new_n413), .B2(KEYINPUT4), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(KEYINPUT75), .A3(KEYINPUT4), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n245), .A2(new_n373), .A3(KEYINPUT76), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT76), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT4), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n412), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n251), .A2(new_n361), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n418), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n410), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n418), .A2(new_n420), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n430), .B1(new_n431), .B2(KEYINPUT4), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n411), .A2(KEYINPUT5), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n422), .A2(new_n427), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g233(.A(G1gat), .B(G29gat), .Z(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G57gat), .B(G85gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT6), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n433), .A2(new_n432), .ZN(new_n443));
  INV_X1    g242(.A(new_n416), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n414), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT76), .B1(new_n245), .B2(new_n373), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n413), .A2(new_n419), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n428), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n411), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n425), .A2(new_n426), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n443), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n439), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n442), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n441), .B1(new_n440), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(G226gat), .A2(G233gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n345), .A2(KEYINPUT74), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT74), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n372), .B2(new_n312), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n461), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n461), .A2(KEYINPUT29), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n345), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n255), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n345), .A2(KEYINPUT74), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n372), .A2(new_n463), .A3(new_n312), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n466), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n372), .A2(new_n461), .A3(new_n312), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n471), .A2(new_n255), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n460), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n255), .A3(new_n472), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n469), .A2(new_n470), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n476), .A2(new_n461), .B1(new_n345), .B2(new_n466), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n475), .B(new_n459), .C1(new_n477), .C2(new_n255), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n474), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n468), .A2(new_n473), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT30), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n459), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n456), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n202), .B1(new_n407), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n479), .A2(new_n482), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n389), .A2(new_n404), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT6), .B1(new_n434), .B2(new_n439), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n453), .B1(new_n434), .B2(KEYINPUT83), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n452), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g290(.A(KEYINPUT85), .B(new_n488), .C1(new_n489), .C2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n492), .A2(new_n441), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n488), .B1(new_n489), .B2(new_n491), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT35), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n282), .B1(new_n270), .B2(new_n279), .ZN(new_n498));
  AND4_X1   g297(.A1(new_n485), .A2(new_n487), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n405), .B2(new_n406), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT73), .B1(new_n486), .B2(new_n500), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT73), .ZN(new_n503));
  AOI211_X1 g302(.A(new_n503), .B(KEYINPUT36), .C1(new_n389), .C2(new_n404), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n496), .A2(new_n441), .A3(new_n478), .A4(new_n492), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n471), .A2(new_n265), .A3(new_n472), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n507), .B(KEYINPUT37), .C1(new_n477), .C2(new_n265), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n475), .B1(new_n477), .B2(new_n255), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n508), .B(new_n460), .C1(new_n509), .C2(KEYINPUT37), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT38), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n460), .A2(KEYINPUT37), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n474), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n511), .B1(new_n509), .B2(KEYINPUT37), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n506), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n418), .A2(new_n420), .A3(new_n410), .A4(new_n424), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n518), .A2(KEYINPUT39), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n428), .B1(new_n418), .B2(new_n420), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n408), .A2(new_n253), .A3(new_n361), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n520), .A2(new_n521), .A3(new_n430), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n519), .B1(new_n522), .B2(new_n410), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT4), .B1(new_n446), .B2(new_n447), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n409), .A3(new_n429), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT39), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n526), .A3(new_n426), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n523), .A2(KEYINPUT40), .A3(new_n439), .A4(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n410), .B1(new_n432), .B2(new_n409), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n453), .B1(new_n531), .B2(new_n526), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(KEYINPUT84), .A3(KEYINPUT40), .A4(new_n523), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n439), .B1(new_n452), .B2(new_n490), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n434), .A2(KEYINPUT83), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n523), .A2(new_n439), .A3(new_n527), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT40), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n479), .A2(new_n540), .A3(new_n482), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n498), .ZN(new_n542));
  OAI22_X1  g341(.A1(new_n517), .A2(new_n542), .B1(new_n483), .B2(new_n498), .ZN(new_n543));
  OAI22_X1  g342(.A1(new_n484), .A2(new_n499), .B1(new_n505), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT89), .ZN(new_n545));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n547));
  NAND2_X1  g346(.A1(G29gat), .A2(G36gat), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  NOR3_X1   g348(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n553));
  INV_X1    g352(.A(G29gat), .ZN(new_n554));
  INV_X1    g353(.A(G36gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(KEYINPUT87), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n548), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G43gat), .B(G50gat), .Z(new_n559));
  XOR2_X1   g358(.A(KEYINPUT88), .B(KEYINPUT15), .Z(new_n560));
  AOI22_X1  g359(.A1(new_n559), .A2(new_n560), .B1(new_n556), .B2(new_n549), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n546), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n547), .A2(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n545), .B1(new_n563), .B2(KEYINPUT17), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n547), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(KEYINPUT89), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT90), .ZN(new_n571));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572));
  INV_X1    g371(.A(G1gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT16), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(G1gat), .B2(new_n572), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G8gat), .ZN(new_n577));
  INV_X1    g376(.A(G8gat), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n575), .B(new_n578), .C1(G1gat), .C2(new_n572), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(new_n563), .B2(KEYINPUT17), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n570), .A2(new_n571), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n580), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(new_n563), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n563), .A2(new_n545), .A3(KEYINPUT17), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT89), .B1(new_n567), .B2(new_n568), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n581), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT90), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(G229gat), .B2(G233gat), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n586), .A2(new_n587), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n591), .A2(new_n585), .A3(new_n582), .A4(new_n593), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT91), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(new_n585), .A3(new_n582), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n592), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT93), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n567), .B(new_n580), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n598), .B(KEYINPUT13), .Z(new_n604));
  AND2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G169gat), .B(G197gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT12), .Z(new_n611));
  NOR2_X1   g410(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n599), .A2(KEYINPUT93), .A3(new_n592), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n597), .A2(new_n602), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n605), .B1(new_n599), .B2(new_n592), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n597), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n617), .B2(new_n611), .ZN(new_n618));
  INV_X1    g417(.A(new_n611), .ZN(new_n619));
  AOI211_X1 g418(.A(KEYINPUT92), .B(new_n619), .C1(new_n597), .C2(new_n616), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n614), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n544), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n623));
  INV_X1    g422(.A(G85gat), .ZN(new_n624));
  INV_X1    g423(.A(G92gat), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(KEYINPUT7), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT7), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n623), .B(new_n629), .C1(new_n624), .C2(new_n625), .ZN(new_n630));
  OR2_X1    g429(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(new_n624), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G99gat), .A2(G106gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT8), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n628), .A2(new_n630), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G99gat), .B(G106gat), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n633), .A2(new_n635), .ZN(new_n639));
  INV_X1    g438(.A(new_n637), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n639), .A2(new_n640), .A3(new_n628), .A4(new_n630), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n641), .A3(KEYINPUT99), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n636), .A2(KEYINPUT99), .A3(new_n637), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(KEYINPUT17), .B2(new_n563), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n570), .ZN(new_n646));
  XNOR2_X1  g445(.A(G190gat), .B(G218gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT100), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n649));
  NAND2_X1  g448(.A1(G232gat), .A2(G233gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n644), .B2(new_n567), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n647), .A2(KEYINPUT100), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n653), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G134gat), .B(G162gat), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n649), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(G71gat), .A2(G78gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(G71gat), .A2(G78gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT94), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT9), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(G64gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(G57gat), .ZN(new_n671));
  INV_X1    g470(.A(G57gat), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(G64gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n669), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n673), .A2(KEYINPUT95), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(KEYINPUT95), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n675), .B(new_n676), .C1(G57gat), .C2(new_n670), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n665), .B1(new_n664), .B2(new_n668), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n667), .A2(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT21), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n583), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT96), .Z(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n241), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(G231gat), .ZN(new_n689));
  INV_X1    g488(.A(G233gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n679), .A2(KEYINPUT21), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n679), .B2(KEYINPUT21), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n348), .ZN(new_n696));
  XOR2_X1   g495(.A(G183gat), .B(G211gat), .Z(new_n697));
  NOR2_X1   g496(.A1(new_n694), .A2(G127gat), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n696), .B2(new_n698), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n688), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n699), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n703), .A2(new_n700), .A3(new_n687), .A4(new_n686), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n679), .A2(new_n641), .A3(new_n638), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n644), .B2(new_n679), .ZN(new_n707));
  NAND2_X1  g506(.A1(G230gat), .A2(G233gat), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT101), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT10), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n713), .B(new_n706), .C1(new_n644), .C2(new_n679), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n644), .A2(KEYINPUT10), .A3(new_n679), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n709), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(G120gat), .B(G148gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(G176gat), .B(G204gat), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n719), .B(new_n720), .Z(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n712), .A2(new_n721), .A3(new_n717), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n663), .A2(new_n705), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT102), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n622), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n455), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n573), .ZN(G1324gat));
  INV_X1    g530(.A(new_n485), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n622), .A2(new_n732), .A3(new_n728), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT16), .B(G8gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT103), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(KEYINPUT42), .A3(new_n736), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n735), .B(KEYINPUT104), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n733), .B1(KEYINPUT42), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(G8gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(G1325gat));
  NAND2_X1  g543(.A1(new_n405), .A2(new_n406), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT36), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n486), .A2(KEYINPUT73), .A3(new_n500), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n486), .A2(new_n500), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n503), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G15gat), .B1(new_n729), .B2(new_n750), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n727), .A2(G15gat), .A3(new_n486), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n622), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1326gat));
  NOR2_X1   g553(.A1(new_n729), .A2(new_n498), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT43), .B(G22gat), .Z(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1327gat));
  INV_X1    g556(.A(new_n663), .ZN(new_n758));
  INV_X1    g557(.A(new_n705), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(new_n759), .A3(new_n725), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n622), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(G29gat), .A3(new_n455), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT45), .Z(new_n763));
  NOR2_X1   g562(.A1(new_n758), .A2(KEYINPUT44), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT107), .B1(new_n505), .B2(new_n543), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n483), .A2(new_n498), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n541), .A2(new_n498), .ZN(new_n768));
  AND4_X1   g567(.A1(new_n441), .A2(new_n496), .A3(new_n478), .A4(new_n492), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT38), .B1(new_n514), .B2(new_n508), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT37), .B1(new_n468), .B2(new_n473), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT38), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n460), .B1(new_n509), .B2(KEYINPUT37), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n769), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n767), .B1(new_n768), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n750), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n766), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n745), .A2(new_n483), .A3(new_n498), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n499), .B1(KEYINPUT35), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n765), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n544), .B2(new_n663), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n725), .B(KEYINPUT106), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n621), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n788), .A2(new_n789), .A3(new_n759), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G29gat), .B1(new_n791), .B2(new_n455), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n763), .A2(new_n792), .ZN(G1328gat));
  NOR3_X1   g592(.A1(new_n761), .A2(G36gat), .A3(new_n485), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT46), .ZN(new_n795));
  OAI21_X1  g594(.A(G36gat), .B1(new_n791), .B2(new_n485), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1329gat));
  NOR2_X1   g596(.A1(new_n486), .A2(G43gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n622), .A2(new_n760), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT108), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n505), .B(new_n790), .C1(new_n783), .C2(new_n785), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G43gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT47), .B1(new_n802), .B2(KEYINPUT109), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n800), .B(new_n802), .C1(KEYINPUT109), .C2(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1330gat));
  INV_X1    g606(.A(new_n498), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n808), .B(new_n790), .C1(new_n783), .C2(new_n785), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G50gat), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n761), .A2(G50gat), .A3(new_n498), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n813));
  XNOR2_X1  g612(.A(new_n812), .B(new_n813), .ZN(G1331gat));
  AOI21_X1  g613(.A(new_n781), .B1(new_n766), .B2(new_n778), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n788), .A2(new_n789), .A3(new_n759), .A4(new_n758), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n456), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G57gat), .ZN(G1332gat));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n485), .B(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n815), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n823));
  AND2_X1   g622(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n822), .B2(new_n823), .ZN(G1333gat));
  XNOR2_X1  g625(.A(new_n486), .B(KEYINPUT112), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n817), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(G71gat), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n505), .A2(G71gat), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n829), .A2(new_n830), .B1(new_n817), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n808), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g634(.A1(new_n723), .A2(new_n724), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n621), .A2(new_n759), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n786), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G85gat), .B1(new_n838), .B2(new_n455), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n779), .A2(new_n782), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n789), .A2(new_n705), .A3(new_n663), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(KEYINPUT51), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n815), .B2(new_n841), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n456), .A2(new_n725), .A3(new_n624), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT113), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n839), .B1(new_n846), .B2(new_n848), .ZN(G1336gat));
  NAND2_X1  g648(.A1(new_n843), .A2(new_n845), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n821), .A2(G92gat), .A3(new_n787), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n821), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(new_n837), .C1(new_n783), .C2(new_n785), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n631), .A2(new_n632), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n852), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n786), .A2(new_n732), .A3(new_n837), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n860), .A2(new_n856), .B1(new_n850), .B2(new_n851), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n859), .B1(new_n861), .B2(new_n858), .ZN(G1337gat));
  OAI21_X1  g661(.A(G99gat), .B1(new_n838), .B2(new_n750), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n486), .A2(G99gat), .A3(new_n836), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n846), .B2(new_n864), .ZN(G1338gat));
  OAI211_X1 g664(.A(new_n808), .B(new_n837), .C1(new_n783), .C2(new_n785), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G106gat), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n787), .A2(G106gat), .A3(new_n498), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT114), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n843), .B2(new_n845), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(KEYINPUT115), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(KEYINPUT115), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT53), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n850), .B2(new_n868), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n867), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1339gat));
  NAND2_X1  g675(.A1(new_n789), .A2(new_n726), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n714), .A2(new_n709), .A3(new_n715), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n717), .A2(KEYINPUT54), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n721), .B1(new_n716), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(KEYINPUT55), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n724), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT55), .B1(new_n880), .B2(new_n882), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n598), .B1(new_n586), .B2(new_n591), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n603), .A2(new_n604), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n610), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n663), .A2(new_n886), .A3(new_n614), .A4(new_n889), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n725), .A2(new_n614), .A3(new_n889), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n621), .B2(new_n886), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n892), .B2(new_n663), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n878), .B1(new_n893), .B2(new_n705), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n455), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT117), .B1(new_n895), .B2(new_n407), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n897));
  INV_X1    g696(.A(new_n407), .ZN(new_n898));
  NOR4_X1   g697(.A1(new_n894), .A2(new_n897), .A3(new_n455), .A4(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n621), .B(new_n821), .C1(new_n896), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n893), .A2(new_n705), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n877), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n853), .A2(new_n455), .A3(new_n486), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n498), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT116), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n902), .A2(new_n906), .A3(new_n498), .A4(new_n903), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n789), .A2(new_n355), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n355), .A2(new_n900), .B1(new_n908), .B2(new_n909), .ZN(G1340gat));
  OAI211_X1 g709(.A(new_n725), .B(new_n821), .C1(new_n896), .C2(new_n899), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n787), .A2(new_n353), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n353), .A2(new_n911), .B1(new_n908), .B2(new_n912), .ZN(G1341gat));
  OAI211_X1 g712(.A(new_n759), .B(new_n821), .C1(new_n896), .C2(new_n899), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(G127gat), .B1(new_n915), .B2(KEYINPUT118), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n705), .A2(new_n348), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n916), .A2(new_n918), .B1(new_n908), .B2(new_n919), .ZN(G1342gat));
  NOR2_X1   g719(.A1(new_n732), .A2(new_n758), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n346), .B(new_n921), .C1(new_n896), .C2(new_n899), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(KEYINPUT56), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT56), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n905), .A2(new_n663), .A3(new_n907), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT119), .A3(G134gat), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT119), .B1(new_n928), .B2(G134gat), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n926), .B(new_n927), .C1(new_n929), .C2(new_n930), .ZN(G1343gat));
  NAND3_X1  g730(.A1(new_n750), .A2(new_n456), .A3(new_n821), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n808), .A2(KEYINPUT57), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n934), .B1(new_n884), .B2(new_n885), .ZN(new_n935));
  INV_X1    g734(.A(new_n885), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n936), .A2(KEYINPUT122), .A3(new_n724), .A4(new_n883), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n891), .B1(new_n938), .B2(new_n621), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n890), .B1(new_n939), .B2(new_n663), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n705), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n933), .B1(new_n941), .B2(new_n877), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n894), .B2(new_n498), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n944), .B2(KEYINPUT121), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n902), .A2(new_n808), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(new_n943), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n932), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n235), .B1(new_n949), .B2(new_n621), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n895), .A2(new_n808), .A3(new_n750), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n853), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n235), .A3(new_n621), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT58), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT58), .ZN(new_n956));
  AOI211_X1 g755(.A(new_n789), .B(new_n932), .C1(new_n945), .C2(new_n948), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n956), .B(new_n953), .C1(new_n957), .C2(new_n235), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n955), .A2(new_n958), .ZN(G1344gat));
  NAND3_X1  g758(.A1(new_n952), .A2(new_n237), .A3(new_n725), .ZN(new_n960));
  AOI211_X1 g759(.A(KEYINPUT59), .B(new_n237), .C1(new_n949), .C2(new_n725), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT59), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n946), .A2(KEYINPUT57), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n941), .B1(new_n621), .B2(new_n727), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n943), .A3(new_n808), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n932), .A2(new_n836), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n962), .B1(new_n968), .B2(G148gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n960), .B1(new_n961), .B2(new_n969), .ZN(G1345gat));
  AOI21_X1  g769(.A(G155gat), .B1(new_n952), .B2(new_n759), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n759), .A2(G155gat), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT123), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n949), .B2(new_n973), .ZN(G1346gat));
  AND2_X1   g773(.A1(new_n949), .A2(new_n663), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n921), .A2(new_n242), .ZN(new_n976));
  OAI22_X1  g775(.A1(new_n975), .A2(new_n242), .B1(new_n951), .B2(new_n976), .ZN(G1347gat));
  NOR4_X1   g776(.A1(new_n894), .A2(new_n456), .A3(new_n898), .A4(new_n821), .ZN(new_n978));
  AOI21_X1  g777(.A(G169gat), .B1(new_n978), .B2(new_n621), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n902), .A2(new_n498), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n485), .A2(new_n456), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n828), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n621), .A2(G169gat), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(G1348gat));
  AOI21_X1  g784(.A(G176gat), .B1(new_n978), .B2(new_n725), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n787), .A2(new_n338), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n983), .B2(new_n987), .ZN(G1349gat));
  NAND3_X1  g787(.A1(new_n978), .A2(new_n308), .A3(new_n759), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n980), .A2(new_n705), .A3(new_n982), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n991));
  OAI21_X1  g790(.A(G183gat), .B1(new_n990), .B2(KEYINPUT124), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(KEYINPUT60), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT60), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n995), .B(new_n989), .C1(new_n991), .C2(new_n992), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1350gat));
  NAND3_X1  g796(.A1(new_n978), .A2(new_n300), .A3(new_n663), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n999));
  INV_X1    g798(.A(new_n982), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n902), .A2(new_n498), .A3(new_n663), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n1002));
  AND4_X1   g801(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .A4(G190gat), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n300), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n1004));
  AOI22_X1  g803(.A1(new_n1001), .A2(new_n1004), .B1(new_n999), .B2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n998), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g805(.A(new_n1006), .B(KEYINPUT126), .ZN(G1351gat));
  AND2_X1   g806(.A1(new_n750), .A2(new_n981), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n966), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(G197gat), .ZN(new_n1010));
  NOR3_X1   g809(.A1(new_n1009), .A2(new_n1010), .A3(new_n789), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n750), .A2(new_n853), .A3(new_n808), .ZN(new_n1012));
  AOI211_X1 g811(.A(new_n456), .B(new_n1012), .C1(new_n901), .C2(new_n877), .ZN(new_n1013));
  AOI21_X1  g812(.A(G197gat), .B1(new_n1013), .B2(new_n621), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n1011), .A2(new_n1014), .ZN(G1352gat));
  NOR2_X1   g814(.A1(new_n836), .A2(G204gat), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  OR2_X1    g816(.A1(new_n1017), .A2(KEYINPUT127), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1017), .A2(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g821(.A(G204gat), .B1(new_n1009), .B2(new_n787), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1018), .A2(KEYINPUT62), .A3(new_n1019), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(G1353gat));
  NAND3_X1  g824(.A1(new_n1013), .A2(new_n212), .A3(new_n759), .ZN(new_n1026));
  NAND4_X1  g825(.A1(new_n963), .A2(new_n965), .A3(new_n759), .A4(new_n1008), .ZN(new_n1027));
  AND3_X1   g826(.A1(new_n1027), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1028));
  AOI21_X1  g827(.A(KEYINPUT63), .B1(new_n1027), .B2(G211gat), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(G1354gat));
  OAI21_X1  g829(.A(G218gat), .B1(new_n1009), .B2(new_n758), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1013), .A2(new_n213), .A3(new_n663), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1031), .A2(new_n1032), .ZN(G1355gat));
endmodule


