//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n201), .A2(G77), .A3(new_n204), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G116), .A2(G270), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G87), .A2(G250), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G50), .B2(G226), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n203), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n210), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT66), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT65), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n229), .A2(G1), .A3(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n204), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n213), .B(new_n226), .C1(new_n234), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  AND2_X1   g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT70), .B1(new_n255), .B2(new_n227), .ZN(new_n256));
  AND2_X1   g0056(.A1(G1), .A2(G13), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT70), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n262), .B1(new_n265), .B2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT69), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n261), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n227), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n273));
  OAI211_X1 g0073(.A(G232), .B(new_n268), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT79), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n265), .B1(new_n256), .B2(new_n260), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT79), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(G232), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n271), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT78), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G223), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G1698), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n286), .A2(new_n288), .B1(G33), .B2(G87), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n255), .B1(new_n228), .B2(new_n230), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n280), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n288), .B1(G223), .B2(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G87), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(KEYINPUT78), .A3(new_n290), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n279), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT80), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT16), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT7), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n284), .A2(new_n285), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(G20), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n293), .A2(new_n294), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT7), .A3(new_n233), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n203), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G58), .A2(G68), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n204), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G20), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n233), .A2(new_n283), .A3(KEYINPUT71), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT71), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(G20), .B2(G33), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G159), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n303), .B1(new_n309), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT7), .B1(new_n307), .B2(new_n233), .ZN(new_n320));
  NOR4_X1   g0120(.A1(new_n293), .A2(new_n294), .A3(new_n304), .A4(G20), .ZN(new_n321));
  OAI21_X1  g0121(.A(G68), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT77), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n312), .B(new_n323), .C1(new_n316), .C2(new_n317), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n317), .B1(new_n313), .B2(new_n315), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n233), .B1(new_n204), .B2(new_n310), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT77), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT16), .A4(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n228), .A2(new_n230), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n319), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  XOR2_X1   g0131(.A(KEYINPUT8), .B(G58), .Z(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n233), .A2(G1), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G13), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n330), .A2(new_n334), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n333), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n256), .A2(new_n260), .B1(new_n269), .B2(new_n268), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n266), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n297), .A2(new_n290), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n274), .A2(KEYINPUT79), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n277), .B1(new_n276), .B2(G232), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT80), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n279), .A2(new_n299), .A3(new_n348), .A4(new_n300), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n302), .A2(new_n339), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n350), .B(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n331), .A2(new_n338), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n345), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n279), .A2(new_n299), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT17), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n353), .A2(new_n358), .A3(KEYINPUT17), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G1698), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n305), .A2(G232), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n305), .A2(G238), .A3(G1698), .ZN(new_n366));
  AND2_X1   g0166(.A1(KEYINPUT72), .A2(G107), .ZN(new_n367));
  NOR2_X1   g0167(.A1(KEYINPUT72), .A2(G107), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n365), .B(new_n366), .C1(new_n305), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n290), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n276), .A2(G244), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n341), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n346), .ZN(new_n375));
  NAND2_X1  g0175(.A1(KEYINPUT15), .A2(G87), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT15), .A2(G87), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n233), .A2(G33), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n379), .A2(new_n381), .B1(G20), .B2(G77), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n316), .B2(new_n333), .ZN(new_n383));
  INV_X1    g0183(.A(G77), .ZN(new_n384));
  INV_X1    g0184(.A(new_n335), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n383), .A2(new_n330), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n330), .A2(new_n384), .A3(new_n334), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT73), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n375), .B(new_n389), .C1(G179), .C2(new_n374), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n352), .A2(new_n363), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n305), .B1(G232), .B2(new_n364), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G226), .A2(G1698), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(new_n283), .B2(new_n206), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n271), .B1(new_n290), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n276), .A2(G238), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n290), .ZN(new_n399));
  AND4_X1   g0199(.A1(new_n392), .A2(new_n399), .A3(new_n397), .A4(new_n341), .ZN(new_n400));
  OAI21_X1  g0200(.A(G169), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n402));
  INV_X1    g0202(.A(new_n400), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n396), .A2(new_n397), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT13), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n405), .A3(G179), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(G169), .C1(new_n398), .C2(new_n400), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n402), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G50), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n316), .A2(new_n410), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n380), .A2(new_n384), .B1(new_n233), .B2(G68), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n330), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT11), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n385), .A2(new_n203), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT12), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(KEYINPUT12), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n416), .A2(new_n417), .B1(new_n337), .B2(G68), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n409), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n403), .A2(new_n405), .A3(G190), .ZN(new_n421));
  OAI21_X1  g0221(.A(G200), .B1(new_n398), .B2(new_n400), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n418), .A4(new_n414), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n276), .A2(G226), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n307), .A2(new_n384), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n364), .A2(G223), .ZN(new_n427));
  NOR2_X1   g0227(.A1(G222), .A2(G1698), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n427), .A2(new_n428), .B1(new_n293), .B2(new_n294), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n426), .A2(new_n290), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n341), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G200), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n335), .A2(G50), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n330), .A2(new_n410), .A3(new_n334), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n332), .A2(new_n381), .ZN(new_n435));
  OAI21_X1  g0235(.A(G20), .B1(new_n201), .B2(new_n204), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n313), .A2(new_n315), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G150), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI211_X1 g0239(.A(new_n433), .B(new_n434), .C1(new_n439), .C2(new_n330), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n432), .B1(new_n440), .B2(KEYINPUT9), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n290), .A2(new_n429), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n426), .B1(new_n340), .B2(new_n266), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n443), .A2(KEYINPUT74), .A3(G190), .A4(new_n425), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n341), .A2(new_n425), .A3(new_n430), .A4(G190), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT74), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n441), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT75), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n439), .A2(new_n330), .ZN(new_n451));
  INV_X1    g0251(.A(new_n434), .ZN(new_n452));
  INV_X1    g0252(.A(new_n433), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT9), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT10), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n450), .A2(KEYINPUT10), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n450), .A2(KEYINPUT10), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n454), .A2(new_n455), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n461), .A2(new_n447), .A3(new_n444), .A4(new_n432), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n459), .B(new_n460), .C1(new_n462), .C2(new_n456), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n443), .A2(new_n300), .A3(new_n425), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n431), .A2(new_n346), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(new_n454), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n458), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n389), .B1(G200), .B2(new_n374), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n374), .A2(new_n356), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR4_X1   g0271(.A1(new_n391), .A2(new_n424), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n222), .A2(new_n364), .ZN(new_n474));
  INV_X1    g0274(.A(G244), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G1698), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n474), .B(new_n476), .C1(new_n293), .C2(new_n294), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n290), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n267), .A2(G45), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n261), .A2(G250), .A3(new_n481), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n481), .A2(new_n258), .A3(new_n262), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G200), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G87), .A2(G97), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n367), .B2(new_n368), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n233), .B1(new_n283), .B2(new_n206), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(KEYINPUT19), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n233), .B(G68), .C1(new_n293), .C2(new_n294), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT19), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n380), .B2(new_n206), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n379), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n494), .A2(new_n330), .B1(new_n385), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n483), .B1(new_n479), .B2(new_n290), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G190), .A3(new_n482), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n228), .A2(new_n230), .A3(new_n329), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n267), .A2(G33), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n499), .A2(new_n335), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G87), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n486), .A2(new_n496), .A3(new_n498), .A4(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n488), .A2(KEYINPUT19), .A3(new_n489), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n491), .A2(new_n493), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n330), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n378), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT83), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(new_n376), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT83), .B1(new_n377), .B2(new_n378), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n511), .A2(new_n499), .A3(new_n335), .A4(new_n500), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n495), .A2(new_n385), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n506), .A2(KEYINPUT84), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n497), .A2(G179), .A3(new_n482), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n346), .B1(new_n497), .B2(new_n482), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT84), .B1(new_n496), .B2(new_n512), .ZN(new_n518));
  OAI211_X1 g0318(.A(KEYINPUT85), .B(new_n503), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n485), .A2(G169), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n497), .A2(G179), .A3(new_n482), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n506), .A2(new_n513), .A3(new_n512), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT84), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n526), .A3(new_n514), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT85), .B1(new_n527), .B2(new_n503), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n307), .A2(G303), .ZN(new_n530));
  OAI211_X1 g0330(.A(G257), .B(new_n364), .C1(new_n293), .C2(new_n294), .ZN(new_n531));
  OAI211_X1 g0331(.A(G264), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n290), .ZN(new_n534));
  XNOR2_X1  g0334(.A(KEYINPUT5), .B(G41), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n483), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n481), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n256), .A2(new_n260), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G270), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n534), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G116), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G20), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n543), .B(new_n233), .C1(G33), .C2(new_n206), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n330), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT20), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n499), .A2(G116), .A3(new_n335), .A4(new_n500), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT20), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n330), .A2(new_n548), .A3(new_n542), .A4(new_n544), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n385), .A2(new_n541), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n546), .A2(new_n547), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n540), .A2(new_n551), .A3(G169), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT21), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT21), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n540), .A2(new_n551), .A3(new_n554), .A4(G169), .ZN(new_n555));
  INV_X1    g0355(.A(new_n540), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n551), .A2(G179), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n553), .A2(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n540), .A2(G200), .ZN(new_n559));
  INV_X1    g0359(.A(new_n551), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n356), .C2(new_n540), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G244), .B(new_n364), .C1(new_n293), .C2(new_n294), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT4), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n305), .A2(KEYINPUT4), .A3(G244), .A4(new_n364), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n305), .A2(G250), .A3(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n543), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n290), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n538), .A2(G257), .B1(new_n535), .B2(new_n483), .ZN(new_n571));
  AOI21_X1  g0371(.A(G169), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n369), .B1(new_n320), .B2(new_n321), .ZN(new_n573));
  XNOR2_X1  g0373(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G97), .A2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n208), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT6), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n577), .A2(KEYINPUT81), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(KEYINPUT81), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n578), .A2(new_n579), .B1(new_n206), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n576), .A2(new_n580), .A3(G20), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n437), .A2(G77), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n573), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n330), .B1(G97), .B2(new_n501), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n335), .A2(G97), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n585), .B(KEYINPUT82), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n572), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n570), .A2(new_n300), .A3(new_n571), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n570), .A2(new_n571), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G200), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n570), .A2(G190), .A3(new_n571), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n591), .A2(new_n584), .A3(new_n586), .A4(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n501), .A2(G107), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n233), .A2(KEYINPUT23), .A3(G107), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n478), .A2(G20), .ZN(new_n597));
  OAI21_X1  g0397(.A(G20), .B1(new_n367), .B2(new_n368), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(KEYINPUT23), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n233), .B(G87), .C1(new_n293), .C2(new_n294), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT22), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT22), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n305), .A2(new_n602), .A3(new_n233), .A4(G87), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT24), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n599), .B2(new_n604), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n330), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n335), .A2(G107), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT25), .ZN(new_n610));
  OAI211_X1 g0410(.A(G257), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n611));
  OAI211_X1 g0411(.A(G250), .B(new_n364), .C1(new_n293), .C2(new_n294), .ZN(new_n612));
  INV_X1    g0412(.A(G294), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n611), .B(new_n612), .C1(new_n283), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n290), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n538), .A2(G264), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n536), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n595), .A2(new_n608), .A3(new_n610), .A4(new_n618), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n617), .A2(new_n356), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(G169), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n300), .B2(new_n617), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n608), .A2(new_n595), .A3(new_n610), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n619), .A2(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n529), .A2(new_n563), .A3(new_n594), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n473), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g0426(.A(new_n626), .B(KEYINPUT86), .Z(G372));
  NAND2_X1  g0427(.A1(new_n458), .A2(new_n463), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n420), .A2(new_n390), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(new_n423), .A3(new_n363), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(new_n352), .ZN(new_n631));
  INV_X1    g0431(.A(new_n466), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n503), .B1(new_n517), .B2(new_n518), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT85), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n583), .A2(new_n330), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n501), .A2(G97), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n586), .ZN(new_n639));
  INV_X1    g0439(.A(new_n572), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n639), .A2(new_n640), .A3(new_n588), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n636), .A2(new_n519), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n523), .A2(new_n524), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n587), .A2(new_n503), .A3(new_n588), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(new_n644), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n623), .A2(new_n622), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n557), .A2(new_n556), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n533), .A2(new_n290), .B1(new_n538), .B2(G270), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n346), .B1(new_n651), .B2(new_n536), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n554), .B1(new_n652), .B2(new_n551), .ZN(new_n653));
  INV_X1    g0453(.A(new_n555), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT87), .B1(new_n649), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n623), .A2(new_n622), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT87), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n558), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n644), .A2(new_n503), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n595), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n601), .A2(new_n603), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n597), .B1(new_n598), .B2(KEYINPUT23), .ZN(new_n665));
  INV_X1    g0465(.A(new_n596), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT24), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n663), .B1(new_n670), .B2(new_n330), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(new_n610), .A3(new_n620), .A4(new_n618), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n662), .A2(new_n672), .A3(new_n589), .A4(new_n593), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n643), .B(new_n648), .C1(new_n660), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n472), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n633), .A2(new_n675), .ZN(G369));
  INV_X1    g0476(.A(G13), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G20), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n267), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n623), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n672), .A2(new_n657), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT88), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n672), .A2(new_n657), .A3(new_n685), .A4(KEYINPUT88), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT89), .ZN(new_n690));
  INV_X1    g0490(.A(new_n684), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n657), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n649), .A2(KEYINPUT89), .A3(new_n684), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n688), .A2(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n691), .A2(new_n560), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n655), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n562), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n657), .A2(new_n684), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n688), .A2(new_n689), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n693), .A2(new_n692), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n655), .A2(new_n691), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n700), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n211), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G1), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n370), .A2(new_n541), .A3(new_n487), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n713), .B1(new_n235), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n617), .A2(new_n522), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n570), .A2(new_n651), .A3(new_n571), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n590), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n617), .A2(new_n522), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT30), .A4(new_n651), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n570), .A2(new_n571), .B1(new_n482), .B2(new_n497), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n300), .A3(new_n540), .A4(new_n617), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n684), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n728), .B(new_n729), .C1(new_n625), .C2(new_n684), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT26), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n636), .A2(new_n732), .A3(new_n519), .A4(new_n641), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n647), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n649), .A2(new_n655), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n733), .B(new_n734), .C1(new_n673), .C2(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n736), .A2(KEYINPUT90), .A3(new_n691), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT90), .B1(new_n736), .B2(new_n691), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT29), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n674), .A2(new_n691), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n731), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n715), .B1(new_n743), .B2(G1), .ZN(G364));
  AOI21_X1  g0544(.A(new_n712), .B1(G45), .B2(new_n678), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n232), .B1(G20), .B2(new_n346), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT91), .Z(new_n751));
  NAND2_X1  g0551(.A1(new_n236), .A2(new_n264), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n709), .A2(new_n305), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n752), .B(new_n753), .C1(new_n250), .C2(new_n264), .ZN(new_n754));
  NAND3_X1  g0554(.A1(G355), .A2(new_n305), .A3(new_n211), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(G116), .C2(new_n211), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n233), .A2(new_n300), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(new_n356), .A3(G200), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n759), .A2(new_n203), .B1(new_n760), .B2(new_n410), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(KEYINPUT92), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT92), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n233), .B2(new_n300), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G77), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n356), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n300), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n233), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n765), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT32), .B1(new_n773), .B2(new_n317), .ZN(new_n774));
  OR3_X1    g0574(.A1(new_n773), .A2(KEYINPUT32), .A3(new_n317), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n767), .A2(new_n771), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  AND3_X1   g0576(.A1(new_n762), .A2(new_n768), .A3(new_n764), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n761), .B(new_n776), .C1(G58), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n307), .B1(new_n780), .B2(G87), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n772), .A2(new_n356), .A3(G200), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n778), .B(new_n781), .C1(new_n207), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  INV_X1    g0584(.A(new_n766), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n759), .ZN(new_n788));
  INV_X1    g0588(.A(G317), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT33), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(KEYINPUT33), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n777), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT94), .ZN(new_n796));
  INV_X1    g0596(.A(new_n773), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n770), .A2(G294), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n307), .C1(new_n799), .C2(new_n782), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n780), .A2(G303), .ZN(new_n802));
  INV_X1    g0602(.A(new_n760), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G326), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n784), .B1(new_n787), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT95), .Z(new_n807));
  INV_X1    g0607(.A(new_n746), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n745), .B(new_n757), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n749), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n697), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n697), .A2(G330), .ZN(new_n812));
  INV_X1    g0612(.A(new_n745), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n698), .A2(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n809), .A2(new_n811), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT96), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n389), .A2(new_n684), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n470), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n390), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n390), .A2(new_n684), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n740), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n674), .A2(new_n691), .A3(new_n823), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(new_n731), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n813), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n746), .A2(new_n747), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n384), .ZN(new_n831));
  INV_X1    g0631(.A(G87), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n771), .B1(new_n832), .B2(new_n782), .C1(new_n785), .C2(new_n541), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n307), .B1(new_n793), .B2(new_n613), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n803), .A2(G303), .B1(new_n797), .B2(G311), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n207), .B2(new_n779), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n759), .A2(new_n799), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n833), .A2(new_n834), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G143), .A2(new_n777), .B1(new_n766), .B2(G159), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n803), .A2(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G150), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n759), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT34), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n770), .A2(G58), .B1(new_n797), .B2(G132), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n843), .A2(new_n305), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n782), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(G68), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n410), .B2(new_n779), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT97), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n838), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n745), .B(new_n831), .C1(new_n850), .C2(new_n808), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT98), .Z(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n748), .B2(new_n823), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n829), .A2(new_n853), .ZN(G384));
  AND4_X1   g0654(.A1(new_n636), .A2(new_n519), .A3(new_n589), .A4(new_n593), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n855), .A2(new_n563), .A3(new_n624), .A4(new_n691), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT102), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n726), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n725), .A2(KEYINPUT102), .A3(new_n684), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n727), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n856), .A2(new_n860), .A3(new_n729), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n472), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT103), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n322), .A2(new_n327), .A3(new_n324), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n303), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n328), .A2(new_n330), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n338), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n682), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n350), .B(KEYINPUT18), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n361), .A2(new_n362), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n353), .A2(new_n358), .B1(new_n867), .B2(new_n868), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n867), .A2(new_n302), .A3(new_n347), .A4(new_n349), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n339), .A2(new_n868), .ZN(new_n878));
  AND4_X1   g0678(.A1(new_n874), .A2(new_n350), .A3(new_n359), .A4(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT100), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n359), .A3(new_n869), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT100), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n350), .A2(new_n359), .A3(new_n874), .A4(new_n878), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n873), .A2(new_n880), .A3(KEYINPUT38), .A4(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n878), .B1(new_n352), .B2(new_n363), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n350), .A2(new_n359), .A3(new_n878), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(new_n874), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n691), .B1(new_n414), .B2(new_n418), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT99), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n420), .A2(new_n423), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n409), .A2(new_n419), .A3(new_n684), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n861), .A2(new_n899), .A3(new_n823), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT40), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  AND4_X1   g0702(.A1(new_n902), .A2(new_n861), .A3(new_n899), .A4(new_n823), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n873), .A2(new_n880), .A3(new_n885), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n887), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n886), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n863), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(G330), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n420), .A2(new_n684), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n905), .B2(new_n886), .ZN(new_n913));
  XOR2_X1   g0713(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n914));
  AND3_X1   g0714(.A1(new_n886), .A2(new_n891), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n911), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n899), .ZN(new_n917));
  INV_X1    g0717(.A(new_n822), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n826), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(new_n906), .B1(new_n871), .B2(new_n682), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n739), .A2(new_n472), .A3(new_n742), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n633), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n921), .B(new_n923), .Z(new_n924));
  XNOR2_X1  g0724(.A(new_n910), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n267), .B2(new_n678), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n576), .A2(new_n580), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT35), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n233), .B(new_n232), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(G116), .C1(new_n928), .C2(new_n927), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT36), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n236), .A2(G77), .A3(new_n310), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n201), .A2(new_n203), .ZN(new_n933));
  OAI211_X1 g0733(.A(G1), .B(new_n677), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n926), .A2(new_n931), .A3(new_n934), .ZN(G367));
  INV_X1    g0735(.A(new_n753), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n750), .B1(new_n211), .B2(new_n495), .C1(new_n246), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n770), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(new_n203), .ZN(new_n939));
  INV_X1    g0739(.A(new_n201), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n785), .A2(new_n940), .B1(new_n384), .B2(new_n782), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n939), .B(new_n941), .C1(G150), .C2(new_n777), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n788), .A2(G159), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n307), .B1(new_n803), .B2(G143), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n780), .A2(G58), .B1(new_n797), .B2(G137), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n788), .A2(G294), .B1(new_n797), .B2(G317), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n206), .B2(new_n782), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n305), .B(new_n948), .C1(G303), .C2(new_n777), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n766), .A2(G283), .B1(new_n369), .B2(new_n770), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT111), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n780), .A2(G116), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT46), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n952), .A2(new_n953), .B1(new_n803), .B2(G311), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n949), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n952), .A2(new_n953), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n946), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT47), .Z(new_n958));
  OAI211_X1 g0758(.A(new_n745), .B(new_n937), .C1(new_n958), .C2(new_n808), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n691), .B1(new_n496), .B2(new_n502), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n661), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n647), .A2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n810), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n639), .A2(new_n684), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n704), .A2(new_n594), .A3(new_n706), .A4(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n589), .A2(new_n593), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n641), .A2(new_n684), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT104), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT104), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n971), .A2(new_n975), .A3(new_n972), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n649), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n589), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT105), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(KEYINPUT105), .A3(new_n589), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(new_n691), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n970), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n963), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n983), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n974), .A2(new_n976), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n700), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n970), .A2(new_n985), .A3(new_n984), .A4(new_n982), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n991), .B1(new_n988), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n710), .B(KEYINPUT41), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT108), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n698), .A2(new_n705), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n694), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n743), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n730), .A2(G330), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n736), .A2(new_n691), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT90), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n736), .A2(KEYINPUT90), .A3(new_n691), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n741), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT29), .B1(new_n674), .B2(new_n691), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1002), .B(new_n1000), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT108), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT107), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT44), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n707), .B2(new_n973), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1011), .A2(KEYINPUT44), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n701), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n694), .B2(new_n705), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n973), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1012), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1013), .A2(new_n1015), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n704), .A2(new_n706), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1022), .A2(KEYINPUT45), .A3(new_n1016), .A4(new_n973), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1016), .B(new_n973), .C1(new_n694), .C2(new_n705), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT45), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1023), .A2(new_n1026), .B1(KEYINPUT109), .B2(new_n699), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n699), .A2(KEYINPUT109), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n1021), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1029), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1001), .B(new_n1010), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n997), .B1(new_n1032), .B2(new_n743), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n267), .B1(new_n678), .B2(G45), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(KEYINPUT110), .B(new_n995), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n743), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1019), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n1014), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n699), .A2(KEYINPUT109), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1028), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1021), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1009), .A2(KEYINPUT108), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n998), .B1(new_n743), .B2(new_n1000), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1038), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1034), .B1(new_n1052), .B2(new_n997), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT110), .B1(new_n1053), .B2(new_n995), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n966), .B1(new_n1037), .B2(new_n1054), .ZN(G387));
  INV_X1    g0855(.A(new_n1051), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n710), .C1(new_n743), .C2(new_n1000), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n745), .B1(new_n704), .B2(new_n810), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n511), .A2(new_n770), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G50), .B2(new_n777), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT113), .Z(new_n1061));
  OAI22_X1  g0861(.A1(new_n782), .A2(new_n206), .B1(new_n773), .B2(new_n841), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n305), .B1(new_n333), .B2(new_n759), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n780), .A2(G77), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n203), .B2(new_n785), .C1(new_n317), .C2(new_n760), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G303), .A2(new_n766), .B1(new_n777), .B2(G317), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n786), .B2(new_n759), .C1(new_n794), .C2(new_n760), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT48), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n799), .B2(new_n938), .C1(new_n613), .C2(new_n779), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT49), .Z(new_n1072));
  AOI21_X1  g0872(.A(new_n305), .B1(new_n797), .B2(G326), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n541), .B2(new_n782), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1067), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT114), .Z(new_n1076));
  AOI21_X1  g0876(.A(new_n1058), .B1(new_n1076), .B2(new_n746), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n333), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n713), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(G68), .A2(G77), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT50), .B1(new_n333), .B2(G50), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1079), .A2(new_n264), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n753), .B(new_n1082), .C1(new_n243), .C2(new_n264), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n713), .A2(new_n211), .A3(new_n305), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(G107), .C2(new_n211), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT112), .Z(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n751), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1077), .A2(new_n1087), .B1(new_n1035), .B2(new_n1000), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1057), .A2(new_n1088), .ZN(G393));
  OR2_X1    g0889(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n710), .A3(new_n1032), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n813), .B1(new_n990), .B2(new_n749), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n777), .A2(G159), .B1(G150), .B2(new_n803), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT51), .Z(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n305), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n940), .A2(new_n759), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n785), .A2(new_n333), .ZN(new_n1097));
  INV_X1    g0897(.A(G143), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n782), .A2(new_n832), .B1(new_n773), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n770), .A2(G77), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(new_n203), .C2(new_n779), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n777), .A2(G311), .B1(G317), .B2(new_n803), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT52), .Z(new_n1105));
  AOI22_X1  g0905(.A1(new_n766), .A2(G294), .B1(G116), .B2(new_n770), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n782), .A2(new_n207), .B1(new_n773), .B2(new_n794), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n305), .B(new_n1107), .C1(G303), .C2(new_n788), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G283), .B2(new_n780), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n746), .B1(new_n1103), .B2(new_n1110), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n750), .B1(new_n206), .B2(new_n211), .C1(new_n253), .C2(new_n936), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1092), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1048), .B2(new_n1035), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1091), .A2(new_n1114), .ZN(G390));
  NOR2_X1   g0915(.A1(new_n913), .A2(new_n915), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n826), .A2(new_n918), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n899), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n911), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1005), .A2(new_n1006), .A3(new_n918), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(new_n820), .A3(new_n899), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n886), .A2(new_n891), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1119), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1116), .A2(new_n1120), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n861), .A2(new_n899), .A3(G330), .A4(new_n823), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT115), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n731), .A2(new_n823), .A3(new_n899), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT115), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1127), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n911), .B1(new_n1117), .B2(new_n899), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1133), .A2(new_n913), .A3(new_n915), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n737), .A2(new_n738), .A3(new_n822), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n821), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1124), .B1(new_n1136), .B2(new_n899), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1131), .B(new_n1132), .C1(new_n1134), .C2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1128), .A2(new_n1035), .A3(new_n1130), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1116), .A2(new_n747), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n307), .B(new_n847), .C1(new_n793), .C2(new_n541), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n766), .A2(G97), .B1(G87), .B2(new_n780), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1142), .A2(new_n1101), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n799), .B2(new_n760), .C1(new_n613), .C2(new_n773), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1141), .B(new_n1144), .C1(new_n369), .C2(new_n788), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT117), .Z(new_n1146));
  NAND2_X1  g0946(.A1(new_n780), .A2(G150), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n938), .A2(new_n317), .B1(new_n782), .B2(new_n940), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1148), .A2(new_n307), .A3(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n777), .A2(G132), .B1(G128), .B2(new_n803), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT116), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n788), .A2(G137), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n797), .A2(G125), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT54), .B(G143), .Z(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n766), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n746), .B1(new_n1146), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n830), .A2(new_n333), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1140), .A2(new_n745), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1139), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n472), .A2(G330), .A3(new_n861), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n922), .A2(new_n1162), .A3(new_n633), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n899), .B1(new_n731), .B2(new_n823), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1117), .B1(new_n1164), .B2(new_n1132), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n861), .A2(G330), .A3(new_n823), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n917), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1129), .B(new_n1167), .C1(new_n821), .C2(new_n1135), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1163), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1128), .A2(new_n1130), .A3(new_n1138), .A4(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1170), .A2(new_n710), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1128), .A2(new_n1130), .A3(new_n1138), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1163), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1161), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(G378));
  NAND2_X1  g0978(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT119), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n467), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n440), .A2(new_n682), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n458), .A2(new_n463), .A3(KEYINPUT119), .A4(new_n466), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1182), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n1185), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1181), .A3(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n908), .B2(G330), .ZN(new_n1197));
  INV_X1    g0997(.A(G330), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1198), .B(new_n1195), .C1(new_n901), .C2(new_n907), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n921), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n861), .A2(new_n823), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1123), .A3(new_n899), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1202), .A2(KEYINPUT40), .B1(new_n906), .B2(new_n903), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1195), .B1(new_n1203), .B2(new_n1198), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n908), .A2(G330), .A3(new_n1196), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n916), .A4(new_n920), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1180), .B1(new_n1200), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1179), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT120), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n921), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1204), .A2(new_n1205), .A3(new_n1209), .A4(new_n921), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1174), .B2(new_n1170), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1208), .B(new_n710), .C1(new_n1214), .C2(KEYINPUT57), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1195), .A2(new_n747), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n766), .A2(new_n511), .B1(G97), .B2(new_n788), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT118), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1218), .B(new_n1065), .C1(new_n202), .C2(new_n782), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n939), .B(new_n1219), .C1(G116), .C2(new_n803), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G41), .B(new_n305), .C1(new_n797), .C2(G283), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n207), .C2(new_n793), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT58), .Z(new_n1223));
  OAI21_X1  g1023(.A(new_n410), .B1(new_n293), .B2(G41), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n777), .A2(G128), .B1(new_n780), .B2(new_n1156), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n766), .A2(G137), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n788), .A2(G132), .B1(new_n770), .B2(G150), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G125), .B2(new_n803), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G41), .B1(new_n1230), .B2(KEYINPUT59), .ZN(new_n1231));
  AOI21_X1  g1031(.A(G33), .B1(new_n797), .B2(G124), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(new_n317), .C2(new_n782), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1224), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n746), .B1(new_n1223), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n830), .A2(new_n940), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1216), .A2(new_n745), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1213), .B2(new_n1034), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1215), .A2(new_n1240), .ZN(G375));
  NAND2_X1  g1041(.A1(new_n917), .A2(new_n747), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n785), .A2(new_n841), .B1(new_n202), .B2(new_n782), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G50), .B2(new_n770), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n803), .A2(G132), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n307), .B1(new_n777), .B2(G137), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n788), .A2(new_n1156), .B1(new_n797), .B2(G128), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n780), .A2(G159), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n759), .A2(new_n541), .B1(new_n782), .B2(new_n384), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n305), .B(new_n1251), .C1(G303), .C2(new_n797), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1059), .B1(G97), .B2(new_n780), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n777), .A2(G283), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n803), .A2(G294), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n785), .A2(new_n370), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1250), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n746), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n830), .A2(new_n203), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1242), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1173), .A2(new_n1035), .B1(new_n745), .B2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1165), .A2(new_n1168), .A3(new_n1163), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n996), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1264), .B2(new_n1169), .ZN(G381));
  NOR3_X1   g1065(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1266));
  XOR2_X1   g1066(.A(new_n1266), .B(KEYINPUT121), .Z(new_n1267));
  INV_X1    g1067(.A(KEYINPUT110), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1032), .A2(new_n743), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1035), .B1(new_n1269), .B2(new_n996), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n995), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1268), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n965), .B1(new_n1272), .B2(new_n1036), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(G390), .A2(G381), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1267), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT122), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1179), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1180), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n711), .B1(new_n1179), .B2(new_n1207), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1239), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1177), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT122), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1267), .A2(new_n1284), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1276), .A2(new_n1283), .A3(new_n1285), .ZN(G407));
  OAI211_X1 g1086(.A(G407), .B(G213), .C1(G343), .C2(new_n1282), .ZN(G409));
  AOI21_X1  g1087(.A(new_n1177), .B1(new_n1215), .B2(new_n1240), .ZN(new_n1288));
  INV_X1    g1088(.A(G213), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1289), .A2(G343), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1179), .A2(new_n1277), .A3(new_n996), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1200), .A2(new_n1206), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1035), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1139), .A2(new_n1160), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1170), .A2(new_n710), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1296), .B(new_n1238), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1291), .B1(new_n1295), .B2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1288), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT60), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1263), .A2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1165), .A2(new_n1168), .A3(new_n1163), .A4(KEYINPUT60), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1303), .A2(new_n1175), .A3(new_n710), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1262), .ZN(new_n1306));
  INV_X1    g1106(.A(G384), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT123), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT123), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1305), .A2(new_n1309), .A3(G384), .A4(new_n1262), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT124), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1306), .A2(new_n1312), .A3(new_n1307), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1311), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT63), .B1(new_n1301), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NOR4_X1   g1119(.A1(new_n1288), .A2(new_n1300), .A3(new_n1316), .A4(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(G393), .B(new_n816), .ZN(new_n1322));
  OAI21_X1  g1122(.A(KEYINPUT127), .B1(new_n1273), .B2(G390), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT127), .ZN(new_n1324));
  INV_X1    g1124(.A(G390), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(G387), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n966), .B(G390), .C1(new_n1037), .C2(new_n1054), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(KEYINPUT126), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1272), .A2(new_n1036), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1330), .A2(new_n1331), .A3(new_n966), .A4(G390), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1322), .B1(new_n1327), .B2(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1273), .A2(G390), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1328), .ZN(new_n1336));
  NOR3_X1   g1136(.A1(new_n1335), .A2(new_n1336), .A3(new_n1322), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1334), .A2(new_n1338), .ZN(new_n1339));
  OR2_X1    g1139(.A1(new_n1291), .A2(KEYINPUT125), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1311), .B(new_n1340), .C1(new_n1313), .C2(new_n1315), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1290), .A2(G2897), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1341), .B(new_n1342), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1177), .A2(new_n1238), .A3(new_n1292), .A4(new_n1294), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1344), .B(new_n1291), .C1(new_n1281), .C2(new_n1177), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT61), .B1(new_n1343), .B2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1321), .A2(new_n1339), .A3(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(KEYINPUT62), .B1(new_n1345), .B2(new_n1316), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1341), .A2(G2897), .A3(new_n1290), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1313), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1314), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1351), .A2(new_n1342), .A3(new_n1340), .A4(new_n1311), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1345), .A2(new_n1349), .A3(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1300), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G375), .A2(G378), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT62), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1354), .A2(new_n1355), .A3(new_n1356), .A4(new_n1317), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT61), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1348), .A2(new_n1353), .A3(new_n1357), .A4(new_n1358), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1323), .A2(new_n1329), .A3(new_n1326), .A4(new_n1332), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1337), .B1(new_n1322), .B2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1359), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1347), .A2(new_n1362), .ZN(G405));
  NAND3_X1  g1163(.A1(new_n1355), .A2(new_n1282), .A3(new_n1316), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1317), .B1(new_n1283), .B2(new_n1288), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1361), .A2(new_n1364), .A3(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1364), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1339), .A2(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1366), .A2(new_n1368), .ZN(G402));
endmodule


