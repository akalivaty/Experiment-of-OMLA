

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600;

  INV_X1 U329 ( .A(KEYINPUT64), .ZN(n483) );
  XNOR2_X1 U330 ( .A(KEYINPUT100), .B(KEYINPUT25), .ZN(n425) );
  XNOR2_X1 U331 ( .A(n426), .B(n425), .ZN(n427) );
  INV_X1 U332 ( .A(G99GAT), .ZN(n387) );
  XNOR2_X1 U333 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U334 ( .A(n406), .B(n311), .ZN(n312) );
  XNOR2_X1 U335 ( .A(n411), .B(n389), .ZN(n390) );
  XNOR2_X1 U336 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U337 ( .A(n486), .B(KEYINPUT55), .ZN(n487) );
  XNOR2_X1 U338 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U339 ( .A(n488), .B(n487), .ZN(n492) );
  XNOR2_X1 U340 ( .A(n399), .B(n398), .ZN(n403) );
  XNOR2_X1 U341 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U342 ( .A(G50GAT), .B(KEYINPUT108), .ZN(n463) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n461) );
  XNOR2_X1 U344 ( .A(n496), .B(n495), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n464), .B(n463), .ZN(G1331GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n298) );
  XNOR2_X1 U347 ( .A(G71GAT), .B(G57GAT), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n333) );
  XNOR2_X1 U349 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n300) );
  AND2_X1 U350 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n301), .B(KEYINPUT32), .ZN(n310) );
  XNOR2_X1 U353 ( .A(G106GAT), .B(G78GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n302), .B(G148GAT), .ZN(n369) );
  XNOR2_X1 U355 ( .A(G99GAT), .B(G85GAT), .ZN(n308) );
  INV_X1 U356 ( .A(G92GAT), .ZN(n303) );
  NAND2_X1 U357 ( .A1(n303), .A2(KEYINPUT71), .ZN(n306) );
  INV_X1 U358 ( .A(KEYINPUT71), .ZN(n304) );
  NAND2_X1 U359 ( .A1(n304), .A2(G92GAT), .ZN(n305) );
  NAND2_X1 U360 ( .A1(n306), .A2(n305), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n353) );
  XNOR2_X1 U362 ( .A(n369), .B(n353), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n313) );
  XOR2_X1 U364 ( .A(G176GAT), .B(G64GAT), .Z(n406) );
  XNOR2_X1 U365 ( .A(G120GAT), .B(G204GAT), .ZN(n311) );
  XOR2_X1 U366 ( .A(n333), .B(n314), .Z(n465) );
  XOR2_X1 U367 ( .A(G169GAT), .B(G8GAT), .Z(n408) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G1GAT), .Z(n330) );
  XNOR2_X1 U369 ( .A(n408), .B(n330), .ZN(n329) );
  XOR2_X1 U370 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n316) );
  NAND2_X1 U371 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U373 ( .A(G141GAT), .B(G22GAT), .Z(n372) );
  XOR2_X1 U374 ( .A(n317), .B(n372), .Z(n327) );
  XOR2_X1 U375 ( .A(G43GAT), .B(G29GAT), .Z(n319) );
  XNOR2_X1 U376 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U378 ( .A(n320), .B(KEYINPUT68), .Z(n322) );
  XNOR2_X1 U379 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n361) );
  XOR2_X1 U381 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n324) );
  XNOR2_X1 U382 ( .A(G197GAT), .B(G113GAT), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n361), .B(n325), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n589) );
  XOR2_X1 U387 ( .A(n589), .B(KEYINPUT69), .Z(n553) );
  INV_X1 U388 ( .A(n553), .ZN(n579) );
  NOR2_X1 U389 ( .A1(n465), .A2(n579), .ZN(n501) );
  XOR2_X1 U390 ( .A(G183GAT), .B(G211GAT), .Z(n405) );
  XOR2_X1 U391 ( .A(n405), .B(G78GAT), .Z(n332) );
  XNOR2_X1 U392 ( .A(n330), .B(G22GAT), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U394 ( .A(G127GAT), .B(G155GAT), .Z(n431) );
  XOR2_X1 U395 ( .A(n333), .B(n431), .Z(n335) );
  NAND2_X1 U396 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U398 ( .A(n337), .B(n336), .Z(n339) );
  XNOR2_X1 U399 ( .A(G8GAT), .B(G64GAT), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n347) );
  XOR2_X1 U401 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n341) );
  XNOR2_X1 U402 ( .A(KEYINPUT14), .B(KEYINPUT79), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U404 ( .A(KEYINPUT81), .B(KEYINPUT77), .Z(n343) );
  XNOR2_X1 U405 ( .A(KEYINPUT80), .B(KEYINPUT78), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U407 ( .A(n345), .B(n344), .Z(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n594) );
  INV_X1 U409 ( .A(n594), .ZN(n497) );
  XOR2_X1 U410 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n349) );
  XNOR2_X1 U411 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U413 ( .A(G190GAT), .B(KEYINPUT75), .Z(n407) );
  XOR2_X1 U414 ( .A(n350), .B(n407), .Z(n352) );
  XNOR2_X1 U415 ( .A(G134GAT), .B(G218GAT), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n357) );
  XOR2_X1 U417 ( .A(KEYINPUT72), .B(G162GAT), .Z(n371) );
  XOR2_X1 U418 ( .A(n371), .B(n353), .Z(n355) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U421 ( .A(n357), .B(n356), .Z(n363) );
  XOR2_X1 U422 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n359) );
  XNOR2_X1 U423 ( .A(KEYINPUT73), .B(KEYINPUT76), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n575) );
  XOR2_X1 U427 ( .A(KEYINPUT36), .B(n575), .Z(n598) );
  XOR2_X1 U428 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n365) );
  XNOR2_X1 U429 ( .A(KEYINPUT22), .B(KEYINPUT85), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U431 ( .A(n366), .B(G155GAT), .Z(n368) );
  XOR2_X1 U432 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n446) );
  XNOR2_X1 U433 ( .A(G50GAT), .B(n446), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U435 ( .A(n370), .B(n369), .Z(n374) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U438 ( .A(KEYINPUT86), .B(G211GAT), .Z(n376) );
  NAND2_X1 U439 ( .A1(G228GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U441 ( .A(n378), .B(n377), .Z(n384) );
  XNOR2_X1 U442 ( .A(G204GAT), .B(KEYINPUT89), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n379), .B(KEYINPUT88), .ZN(n380) );
  XOR2_X1 U444 ( .A(n380), .B(KEYINPUT21), .Z(n382) );
  XNOR2_X1 U445 ( .A(G197GAT), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n419) );
  XNOR2_X1 U447 ( .A(n419), .B(KEYINPUT23), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n485) );
  XOR2_X1 U449 ( .A(KEYINPUT17), .B(KEYINPUT83), .Z(n386) );
  XNOR2_X1 U450 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n411) );
  XNOR2_X1 U452 ( .A(G43GAT), .B(KEYINPUT84), .ZN(n388) );
  XOR2_X1 U453 ( .A(n390), .B(G190GAT), .Z(n399) );
  XOR2_X1 U454 ( .A(G15GAT), .B(G71GAT), .Z(n392) );
  NAND2_X1 U455 ( .A1(G227GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U457 ( .A(G169GAT), .B(n393), .ZN(n397) );
  XOR2_X1 U458 ( .A(G127GAT), .B(G176GAT), .Z(n395) );
  XNOR2_X1 U459 ( .A(KEYINPUT20), .B(G183GAT), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U461 ( .A(KEYINPUT82), .B(G134GAT), .Z(n401) );
  XNOR2_X1 U462 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U464 ( .A(G113GAT), .B(n402), .ZN(n436) );
  XNOR2_X1 U465 ( .A(n403), .B(n436), .ZN(n550) );
  INV_X1 U466 ( .A(n550), .ZN(n542) );
  NAND2_X1 U467 ( .A1(n485), .A2(n542), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n404), .B(KEYINPUT26), .ZN(n587) );
  INV_X1 U469 ( .A(n587), .ZN(n422) );
  XOR2_X1 U470 ( .A(n406), .B(n405), .Z(n410) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n415) );
  XOR2_X1 U473 ( .A(KEYINPUT97), .B(n411), .Z(n413) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U476 ( .A(n415), .B(n414), .Z(n421) );
  XOR2_X1 U477 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n417) );
  XNOR2_X1 U478 ( .A(G36GAT), .B(G92GAT), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n540) );
  XOR2_X1 U482 ( .A(n540), .B(KEYINPUT27), .Z(n452) );
  NAND2_X1 U483 ( .A1(n422), .A2(n452), .ZN(n428) );
  NOR2_X1 U484 ( .A1(n542), .A2(n540), .ZN(n423) );
  XOR2_X1 U485 ( .A(KEYINPUT99), .B(n423), .Z(n424) );
  NOR2_X1 U486 ( .A1(n485), .A2(n424), .ZN(n426) );
  NAND2_X1 U487 ( .A1(n428), .A2(n427), .ZN(n451) );
  XOR2_X1 U488 ( .A(KEYINPUT90), .B(G85GAT), .Z(n430) );
  XNOR2_X1 U489 ( .A(G141GAT), .B(G148GAT), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U491 ( .A(n432), .B(n431), .Z(n434) );
  XNOR2_X1 U492 ( .A(G29GAT), .B(G162GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U494 ( .A(n436), .B(n435), .Z(n450) );
  XOR2_X1 U495 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n438) );
  XNOR2_X1 U496 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U498 ( .A(G57GAT), .B(KEYINPUT91), .Z(n440) );
  XNOR2_X1 U499 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U501 ( .A(n442), .B(n441), .Z(n448) );
  XOR2_X1 U502 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n444) );
  NAND2_X1 U503 ( .A1(G225GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n515) );
  INV_X1 U508 ( .A(n515), .ZN(n538) );
  NAND2_X1 U509 ( .A1(n451), .A2(n538), .ZN(n456) );
  NAND2_X1 U510 ( .A1(n515), .A2(n452), .ZN(n548) );
  XOR2_X1 U511 ( .A(n485), .B(KEYINPUT28), .Z(n551) );
  INV_X1 U512 ( .A(n551), .ZN(n512) );
  NOR2_X1 U513 ( .A1(n548), .A2(n512), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n453), .B(KEYINPUT98), .ZN(n454) );
  NAND2_X1 U515 ( .A1(n454), .A2(n542), .ZN(n455) );
  NAND2_X1 U516 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n457), .B(KEYINPUT101), .ZN(n500) );
  NOR2_X1 U518 ( .A1(n598), .A2(n500), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n497), .A2(n458), .ZN(n459) );
  XNOR2_X1 U520 ( .A(KEYINPUT37), .B(n459), .ZN(n537) );
  NAND2_X1 U521 ( .A1(n501), .A2(n537), .ZN(n460) );
  XOR2_X1 U522 ( .A(KEYINPUT38), .B(n460), .Z(n520) );
  NAND2_X1 U523 ( .A1(n520), .A2(n550), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  NAND2_X1 U525 ( .A1(n520), .A2(n512), .ZN(n464) );
  INV_X1 U526 ( .A(KEYINPUT41), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n466), .B(n465), .ZN(n569) );
  INV_X1 U528 ( .A(n569), .ZN(n522) );
  INV_X1 U529 ( .A(KEYINPUT47), .ZN(n472) );
  AND2_X1 U530 ( .A1(n569), .A2(n589), .ZN(n467) );
  XNOR2_X1 U531 ( .A(n467), .B(KEYINPUT46), .ZN(n468) );
  XNOR2_X1 U532 ( .A(KEYINPUT114), .B(n594), .ZN(n582) );
  NOR2_X1 U533 ( .A1(n468), .A2(n582), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n469), .B(KEYINPUT115), .ZN(n470) );
  NOR2_X1 U535 ( .A1(n470), .A2(n575), .ZN(n471) );
  XNOR2_X1 U536 ( .A(n472), .B(n471), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n497), .A2(n598), .ZN(n473) );
  XNOR2_X1 U538 ( .A(n473), .B(KEYINPUT45), .ZN(n475) );
  INV_X1 U539 ( .A(n465), .ZN(n474) );
  NAND2_X1 U540 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U541 ( .A1(n553), .A2(n476), .ZN(n477) );
  XNOR2_X1 U542 ( .A(KEYINPUT116), .B(n477), .ZN(n478) );
  NOR2_X1 U543 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n480), .B(KEYINPUT48), .ZN(n547) );
  NOR2_X1 U545 ( .A1(n547), .A2(n540), .ZN(n481) );
  XOR2_X1 U546 ( .A(KEYINPUT54), .B(n481), .Z(n482) );
  NOR2_X1 U547 ( .A1(n482), .A2(n515), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n484), .B(n483), .ZN(n588) );
  NOR2_X1 U549 ( .A1(n485), .A2(n588), .ZN(n488) );
  INV_X1 U550 ( .A(KEYINPUT124), .ZN(n486) );
  NAND2_X1 U551 ( .A1(n492), .A2(n550), .ZN(n578) );
  NOR2_X1 U552 ( .A1(n522), .A2(n578), .ZN(n491) );
  XNOR2_X1 U553 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n489), .B(G176GAT), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(G1349GAT) );
  AND2_X1 U556 ( .A1(n492), .A2(n550), .ZN(n583) );
  AND2_X1 U557 ( .A1(n583), .A2(n575), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT58), .B(KEYINPUT126), .ZN(n494) );
  INV_X1 U559 ( .A(G190GAT), .ZN(n493) );
  XOR2_X1 U560 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n504) );
  NOR2_X1 U561 ( .A1(n575), .A2(n497), .ZN(n498) );
  XOR2_X1 U562 ( .A(KEYINPUT16), .B(n498), .Z(n499) );
  NOR2_X1 U563 ( .A1(n500), .A2(n499), .ZN(n523) );
  NAND2_X1 U564 ( .A1(n501), .A2(n523), .ZN(n502) );
  XOR2_X1 U565 ( .A(KEYINPUT102), .B(n502), .Z(n513) );
  NAND2_X1 U566 ( .A1(n515), .A2(n513), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G1GAT), .B(n505), .ZN(G1324GAT) );
  INV_X1 U569 ( .A(n540), .ZN(n519) );
  NAND2_X1 U570 ( .A1(n513), .A2(n519), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(KEYINPUT104), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G8GAT), .B(n507), .ZN(G1325GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT35), .B(KEYINPUT106), .Z(n509) );
  NAND2_X1 U574 ( .A1(n513), .A2(n550), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n511) );
  XOR2_X1 U576 ( .A(G15GAT), .B(KEYINPUT105), .Z(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1326GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U580 ( .A1(n520), .A2(n515), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(KEYINPUT107), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(G1328GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G36GAT), .ZN(G1329GAT) );
  NOR2_X1 U586 ( .A1(n589), .A2(n522), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n536), .A2(n523), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(KEYINPUT110), .ZN(n532) );
  NOR2_X1 U589 ( .A1(n538), .A2(n532), .ZN(n528) );
  XOR2_X1 U590 ( .A(KEYINPUT109), .B(KEYINPUT111), .Z(n526) );
  XNOR2_X1 U591 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1332GAT) );
  NOR2_X1 U594 ( .A1(n540), .A2(n532), .ZN(n529) );
  XOR2_X1 U595 ( .A(G64GAT), .B(n529), .Z(G1333GAT) );
  NOR2_X1 U596 ( .A1(n542), .A2(n532), .ZN(n530) );
  XOR2_X1 U597 ( .A(KEYINPUT112), .B(n530), .Z(n531) );
  XNOR2_X1 U598 ( .A(G71GAT), .B(n531), .ZN(G1334GAT) );
  XNOR2_X1 U599 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n534) );
  NOR2_X1 U600 ( .A1(n551), .A2(n532), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U602 ( .A(G78GAT), .B(n535), .Z(G1335GAT) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n544) );
  NOR2_X1 U604 ( .A1(n538), .A2(n544), .ZN(n539) );
  XOR2_X1 U605 ( .A(G85GAT), .B(n539), .Z(G1336GAT) );
  NOR2_X1 U606 ( .A1(n540), .A2(n544), .ZN(n541) );
  XOR2_X1 U607 ( .A(G92GAT), .B(n541), .Z(G1337GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n544), .ZN(n543) );
  XOR2_X1 U609 ( .A(G99GAT), .B(n543), .Z(G1338GAT) );
  NOR2_X1 U610 ( .A1(n551), .A2(n544), .ZN(n545) );
  XOR2_X1 U611 ( .A(KEYINPUT44), .B(n545), .Z(n546) );
  XNOR2_X1 U612 ( .A(G106GAT), .B(n546), .ZN(G1339GAT) );
  NOR2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(KEYINPUT117), .ZN(n565) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U616 ( .A1(n565), .A2(n552), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n562), .A2(n553), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U619 ( .A(G113GAT), .B(n555), .ZN(G1340GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n557) );
  NAND2_X1 U621 ( .A1(n562), .A2(n569), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U623 ( .A(G120GAT), .B(n558), .Z(G1341GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n560) );
  NAND2_X1 U625 ( .A1(n562), .A2(n582), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(G127GAT), .B(n561), .Z(G1342GAT) );
  XOR2_X1 U628 ( .A(G134GAT), .B(KEYINPUT51), .Z(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n575), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1343GAT) );
  NOR2_X1 U631 ( .A1(n587), .A2(n565), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT121), .B(n566), .Z(n576) );
  NAND2_X1 U633 ( .A1(n576), .A2(n589), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G141GAT), .B(n568), .ZN(G1344GAT) );
  XOR2_X1 U636 ( .A(G148GAT), .B(KEYINPUT52), .Z(n571) );
  NAND2_X1 U637 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(G1345GAT) );
  NAND2_X1 U641 ( .A1(n594), .A2(n576), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n577), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G169GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1348GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n586) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n591) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n596) );
  NAND2_X1 U654 ( .A1(n589), .A2(n596), .ZN(n590) );
  XOR2_X1 U655 ( .A(n591), .B(n590), .Z(G1352GAT) );
  XOR2_X1 U656 ( .A(G204GAT), .B(KEYINPUT61), .Z(n593) );
  NAND2_X1 U657 ( .A1(n596), .A2(n465), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1353GAT) );
  NAND2_X1 U659 ( .A1(n594), .A2(n596), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n595), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U661 ( .A(n596), .ZN(n597) );
  NOR2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U663 ( .A(KEYINPUT62), .B(n599), .Z(n600) );
  XNOR2_X1 U664 ( .A(G218GAT), .B(n600), .ZN(G1355GAT) );
endmodule

