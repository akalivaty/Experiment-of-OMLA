//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  AND2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(KEYINPUT26), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n208), .A2(KEYINPUT65), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT65), .B1(new_n208), .B2(new_n209), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n214), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT27), .B(G183gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT64), .B(KEYINPUT28), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(new_n219), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n212), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n213), .ZN(new_n229));
  NAND3_X1  g028(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n204), .A3(new_n205), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n203), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT25), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n231), .A2(new_n235), .A3(KEYINPUT25), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n227), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n240));
  OAI21_X1  g039(.A(G134gat), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G127gat), .ZN(new_n242));
  INV_X1    g041(.A(G134gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n241), .B(new_n244), .C1(KEYINPUT1), .C2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n248));
  INV_X1    g047(.A(G113gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(G120gat), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(G113gat), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n247), .B(new_n248), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n238), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT32), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT33), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G71gat), .B(G99gat), .Z(new_n262));
  XNOR2_X1  g061(.A(G15gat), .B(G43gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n238), .A2(new_n254), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n238), .A2(new_n254), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n256), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT34), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n260), .B1(new_n264), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n271), .B2(new_n264), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT32), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n265), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n256), .B1(new_n266), .B2(new_n267), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT32), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n264), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n276), .A2(KEYINPUT33), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n268), .B(KEYINPUT34), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285));
  INV_X1    g084(.A(G211gat), .ZN(new_n286));
  INV_X1    g085(.A(G218gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT71), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G218gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n286), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(KEYINPUT70), .B(KEYINPUT22), .Z(new_n292));
  OAI21_X1  g091(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT71), .B(G218gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n297), .B1(new_n298), .B2(new_n286), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(new_n294), .A3(new_n285), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n294), .B1(new_n299), .B2(new_n285), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT74), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G141gat), .B(G148gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313));
  INV_X1    g112(.A(G148gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G141gat), .ZN(new_n315));
  INV_X1    g114(.A(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G155gat), .B(G162gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n320));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(KEYINPUT2), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n312), .A2(new_n313), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G228gat), .ZN(new_n328));
  INV_X1    g127(.A(G233gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n319), .B1(new_n318), .B2(new_n322), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n301), .A2(new_n325), .A3(new_n304), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(new_n313), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n312), .A2(new_n323), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT29), .B1(new_n296), .B2(new_n300), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(KEYINPUT3), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n330), .B1(new_n327), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI211_X1 g142(.A(KEYINPUT82), .B(new_n330), .C1(new_n327), .C2(new_n340), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n337), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G22gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT83), .ZN(new_n347));
  INV_X1    g146(.A(G22gat), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n337), .B(new_n348), .C1(new_n343), .C2(new_n344), .ZN(new_n349));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT31), .B(G50gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n346), .A2(new_n347), .A3(new_n349), .A4(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(KEYINPUT83), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n355), .A2(new_n352), .B1(new_n346), .B2(new_n349), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n202), .B(new_n284), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT0), .ZN(new_n359));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n246), .A2(new_n312), .A3(new_n323), .A4(new_n253), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT4), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n334), .A2(new_n368), .A3(new_n253), .A4(new_n246), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(KEYINPUT77), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT4), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n338), .A2(KEYINPUT3), .B1(new_n253), .B2(new_n246), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT75), .B1(new_n374), .B2(new_n324), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT3), .B1(new_n332), .B2(new_n333), .ZN(new_n376));
  AND4_X1   g175(.A1(KEYINPUT75), .A2(new_n376), .A3(new_n324), .A4(new_n254), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n373), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT78), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n369), .A2(new_n370), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n362), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT76), .B1(new_n362), .B2(KEYINPUT4), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT78), .ZN(new_n387));
  INV_X1    g186(.A(new_n373), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n376), .A2(new_n324), .A3(new_n254), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n374), .A2(KEYINPUT75), .A3(new_n324), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n386), .A2(new_n387), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n254), .A2(new_n338), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n369), .A2(new_n370), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n388), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT5), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n379), .A2(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n362), .A2(new_n381), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n404), .B1(new_n380), .B2(KEYINPUT4), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(new_n378), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT6), .B(new_n361), .C1(new_n402), .C2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n361), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n372), .A2(new_n378), .A3(KEYINPUT78), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n387), .B1(new_n386), .B2(new_n393), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT79), .B1(new_n397), .B2(KEYINPUT5), .ZN(new_n413));
  INV_X1    g212(.A(new_n401), .ZN(new_n414));
  OAI22_X1  g213(.A1(new_n411), .A2(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n408), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n410), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n410), .B1(new_n407), .B2(new_n378), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n418), .B1(new_n402), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n409), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n305), .ZN(new_n422));
  NAND2_X1  g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n238), .B2(new_n325), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n231), .A2(new_n235), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT25), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n231), .A2(new_n235), .A3(KEYINPUT25), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n423), .B1(new_n430), .B2(new_n227), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n422), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n238), .A2(new_n424), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT29), .B1(new_n430), .B2(new_n227), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n433), .B(new_n305), .C1(new_n434), .C2(new_n424), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G8gat), .B(G36gat), .Z(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT73), .ZN(new_n438));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT30), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n440), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n421), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT87), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n421), .A2(new_n447), .A3(new_n444), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n357), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n379), .A2(new_n394), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n400), .A2(new_n401), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n419), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n450), .B1(new_n453), .B2(KEYINPUT6), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT80), .B(new_n418), .C1(new_n402), .C2(new_n419), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n361), .B1(new_n402), .B2(new_n408), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT81), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(new_n459), .A3(new_n455), .A4(new_n456), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n460), .A3(new_n409), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n265), .B(new_n274), .C1(KEYINPUT68), .C2(new_n270), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT68), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n280), .A2(new_n463), .A3(new_n281), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n331), .A2(new_n336), .ZN(new_n466));
  INV_X1    g265(.A(new_n300), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n325), .B1(new_n467), .B2(new_n302), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n334), .B1(new_n468), .B2(new_n313), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n301), .A2(new_n304), .B1(new_n325), .B2(new_n324), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT82), .B1(new_n471), .B2(new_n330), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n341), .A2(new_n342), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n347), .B1(new_n474), .B2(new_n348), .ZN(new_n475));
  INV_X1    g274(.A(new_n352), .ZN(new_n476));
  INV_X1    g275(.A(new_n349), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n472), .A2(new_n473), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n348), .B1(new_n478), .B2(new_n337), .ZN(new_n479));
  OAI22_X1  g278(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n465), .B1(new_n480), .B2(new_n353), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n444), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n449), .B1(new_n482), .B2(KEYINPUT35), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT84), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n354), .B2(new_n356), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(KEYINPUT84), .A3(new_n353), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n461), .B2(new_n444), .ZN(new_n488));
  INV_X1    g287(.A(new_n419), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT6), .B1(new_n415), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n456), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT38), .ZN(new_n492));
  INV_X1    g291(.A(new_n440), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n432), .A2(new_n494), .A3(new_n435), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n432), .B2(new_n435), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n492), .B(new_n493), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n442), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n436), .A2(KEYINPUT37), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n432), .A2(new_n494), .A3(new_n435), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n492), .B1(new_n501), .B2(new_n493), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n491), .A2(new_n503), .A3(new_n409), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n480), .A2(new_n353), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n403), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n375), .A2(new_n377), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n388), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT39), .ZN(new_n511));
  INV_X1    g310(.A(new_n396), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n373), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n391), .A2(new_n392), .ZN(new_n515));
  AOI211_X1 g314(.A(KEYINPUT39), .B(new_n373), .C1(new_n405), .C2(new_n515), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n516), .A2(KEYINPUT85), .A3(new_n361), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT85), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n511), .B(new_n388), .C1(new_n508), .C2(new_n509), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(new_n410), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT40), .B(new_n514), .C1(new_n517), .C2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(new_n443), .A3(new_n456), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT86), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT85), .B1(new_n516), .B2(new_n361), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n518), .A3(new_n410), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n524), .A2(new_n525), .B1(new_n510), .B2(new_n513), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n523), .B1(new_n526), .B2(KEYINPUT40), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n514), .B1(new_n517), .B2(new_n520), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT40), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(KEYINPUT86), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n522), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g330(.A(KEYINPUT69), .B(KEYINPUT36), .C1(new_n275), .C2(new_n282), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT36), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT36), .B1(new_n275), .B2(new_n282), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT69), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI22_X1  g335(.A1(new_n506), .A2(new_n531), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n488), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT88), .B1(new_n483), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n536), .A2(new_n532), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n504), .A2(new_n505), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n527), .A2(new_n530), .ZN(new_n542));
  INV_X1    g341(.A(new_n522), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n540), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n457), .A2(KEYINPUT81), .B1(KEYINPUT6), .B2(new_n417), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n443), .B1(new_n546), .B2(new_n460), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n547), .B2(new_n487), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT88), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n202), .B1(new_n547), .B2(new_n481), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n449), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n539), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G113gat), .B(G141gat), .Z(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT89), .B(G197gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT11), .B(G169gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n555), .B(new_n556), .Z(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT12), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G15gat), .B(G22gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT16), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(G1gat), .ZN(new_n562));
  INV_X1    g361(.A(G8gat), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n562), .B(new_n563), .C1(G1gat), .C2(new_n560), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT91), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n560), .A2(G1gat), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n562), .B1(new_n566), .B2(KEYINPUT90), .ZN(new_n568));
  OAI21_X1  g367(.A(G8gat), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G29gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT14), .ZN(new_n572));
  INV_X1    g371(.A(G36gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G43gat), .B(G50gat), .Z(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n571), .A2(KEYINPUT14), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n575), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(KEYINPUT15), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n582), .A2(new_n574), .A3(new_n577), .A4(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n570), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT13), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n565), .A2(new_n569), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(KEYINPUT17), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n584), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n570), .A2(new_n584), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(KEYINPUT92), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(new_n592), .A3(new_n598), .A4(new_n594), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n597), .A2(new_n599), .B1(G229gat), .B2(G233gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n590), .B1(new_n600), .B2(KEYINPUT18), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(KEYINPUT92), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n604), .A2(KEYINPUT18), .A3(new_n587), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n559), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n587), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT18), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n600), .A2(KEYINPUT18), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n590), .A4(new_n558), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  XOR2_X1   g413(.A(G57gat), .B(G64gat), .Z(new_n615));
  AOI21_X1  g414(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(KEYINPUT93), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(KEYINPUT93), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G71gat), .B(G78gat), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n619), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G99gat), .B(G106gat), .Z(new_n623));
  OR2_X1    g422(.A1(new_n623), .A2(KEYINPUT97), .ZN(new_n624));
  INV_X1    g423(.A(G99gat), .ZN(new_n625));
  INV_X1    g424(.A(G106gat), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT8), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(G85gat), .B2(G92gat), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n628), .B1(KEYINPUT97), .B2(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(G85gat), .A2(G92gat), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT7), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n630), .B2(KEYINPUT7), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT95), .B1(new_n630), .B2(KEYINPUT7), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n630), .A2(KEYINPUT95), .A3(KEYINPUT7), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n624), .B1(new_n629), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n629), .A2(new_n624), .A3(new_n636), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n622), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n637), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n619), .B(new_n620), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n614), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n638), .B2(new_n637), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n644), .A2(KEYINPUT10), .A3(new_n641), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n639), .A2(new_n642), .A3(new_n649), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(G120gat), .B(G148gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT99), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n650), .A2(new_n651), .A3(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G155gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G183gat), .B(G211gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(G231gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n329), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n641), .A2(KEYINPUT21), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n668), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT21), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n622), .B2(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n669), .A2(new_n672), .A3(G127gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n570), .B1(KEYINPUT21), .B2(new_n641), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G127gat), .B1(new_n669), .B2(new_n672), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n676), .B1(new_n674), .B2(new_n677), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n666), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n680), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n678), .A3(new_n665), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(G232gat), .A2(G233gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(KEYINPUT41), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT94), .ZN(new_n688));
  XNOR2_X1  g487(.A(G134gat), .B(G162gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n644), .A2(new_n646), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n692), .A2(new_n584), .B1(KEYINPUT41), .B2(new_n686), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n592), .A3(new_n594), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(G190gat), .B(G218gat), .Z(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n696), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n693), .A2(new_n698), .A3(new_n694), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n690), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n697), .A2(new_n690), .A3(new_n699), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n661), .A2(new_n684), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n552), .A2(new_n613), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n461), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n443), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT16), .B(G8gat), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n710), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n708), .ZN(new_n711));
  INV_X1    g510(.A(new_n710), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(G1325gat));
  AOI21_X1  g517(.A(G15gat), .B1(new_n704), .B2(new_n284), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n540), .A2(KEYINPUT102), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n540), .A2(KEYINPUT102), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G15gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT103), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n719), .B1(new_n704), .B2(new_n725), .ZN(G1326gat));
  INV_X1    g525(.A(new_n487), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n704), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT43), .B(G22gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731));
  INV_X1    g530(.A(new_n702), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n700), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n539), .A2(new_n551), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n613), .A2(new_n684), .A3(new_n660), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n461), .A2(G29gat), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n731), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n736), .A2(KEYINPUT45), .A3(new_n737), .A4(new_n739), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n737), .B(KEYINPUT104), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT105), .B1(new_n488), .B2(new_n537), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n545), .B(new_n746), .C1(new_n547), .C2(new_n487), .ZN(new_n747));
  AOI211_X1 g546(.A(KEYINPUT106), .B(new_n483), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n747), .ZN(new_n750));
  INV_X1    g549(.A(new_n483), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n734), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n748), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n735), .A2(KEYINPUT44), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n744), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n758), .A2(new_n705), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n741), .B(new_n742), .C1(new_n759), .C2(new_n571), .ZN(G1328gat));
  NOR2_X1   g559(.A1(new_n444), .A2(G36gat), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  OR3_X1    g561(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT46), .B1(new_n738), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n758), .A2(new_n443), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n766), .B(KEYINPUT107), .C1(new_n767), .C2(new_n573), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n573), .B1(new_n758), .B2(new_n443), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(new_n765), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(G1329gat));
  NOR3_X1   g571(.A1(new_n738), .A2(G43gat), .A3(new_n283), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n723), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(G43gat), .ZN(new_n775));
  INV_X1    g574(.A(G43gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n758), .B2(new_n540), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n775), .A2(KEYINPUT47), .B1(new_n777), .B2(new_n779), .ZN(G1330gat));
  NOR3_X1   g579(.A1(new_n738), .A2(G50gat), .A3(new_n487), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n758), .A2(new_n727), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n782), .B2(G50gat), .ZN(new_n783));
  INV_X1    g582(.A(G50gat), .ZN(new_n784));
  INV_X1    g583(.A(new_n505), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n758), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT48), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n783), .A2(KEYINPUT48), .B1(new_n786), .B2(new_n788), .ZN(G1331gat));
  NOR2_X1   g588(.A1(new_n612), .A2(new_n661), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(new_n684), .A3(new_n733), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n748), .A2(new_n752), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n461), .ZN(new_n793));
  XOR2_X1   g592(.A(KEYINPUT108), .B(G57gat), .Z(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1332gat));
  AOI21_X1  g594(.A(new_n444), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n792), .A2(KEYINPUT109), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT109), .B1(new_n792), .B2(new_n797), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1333gat));
  OAI21_X1  g601(.A(G71gat), .B1(new_n792), .B2(new_n722), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n283), .A2(G71gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n792), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g605(.A1(new_n792), .A2(new_n487), .ZN(new_n807));
  XNOR2_X1  g606(.A(KEYINPUT110), .B(G78gat), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1335gat));
  INV_X1    g608(.A(new_n684), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n790), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n757), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n755), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G85gat), .B1(new_n814), .B2(new_n461), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n461), .A2(new_n444), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n727), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n746), .B1(new_n817), .B2(new_n545), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n488), .A2(new_n537), .A3(KEYINPUT105), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n751), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n734), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n483), .B1(new_n745), .B2(new_n747), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT111), .B1(new_n823), .B2(new_n733), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n612), .A2(new_n684), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n822), .A2(new_n824), .A3(KEYINPUT51), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n461), .A2(G85gat), .A3(new_n661), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n832), .ZN(G1336gat));
  OAI21_X1  g632(.A(G92gat), .B1(new_n814), .B2(new_n444), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n661), .A2(G92gat), .A3(new_n444), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n834), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(G1337gat));
  NAND4_X1  g640(.A1(new_n830), .A2(new_n625), .A3(new_n284), .A4(new_n660), .ZN(new_n842));
  OAI21_X1  g641(.A(G99gat), .B1(new_n814), .B2(new_n722), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1338gat));
  AOI21_X1  g643(.A(new_n811), .B1(new_n756), .B2(new_n757), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n626), .B1(new_n845), .B2(new_n727), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n505), .A2(new_n661), .A3(G106gat), .ZN(new_n847));
  INV_X1    g646(.A(new_n825), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n823), .A2(new_n733), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n821), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT51), .B1(new_n850), .B2(new_n824), .ZN(new_n851));
  INV_X1    g650(.A(new_n829), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n846), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n785), .B(new_n812), .C1(new_n755), .C2(new_n813), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G106gat), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n859));
  AND4_X1   g658(.A1(new_n856), .A2(new_n858), .A3(new_n853), .A4(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT53), .B1(new_n830), .B2(new_n847), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n856), .B1(new_n861), .B2(new_n858), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n855), .B1(new_n860), .B2(new_n862), .ZN(G1339gat));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864));
  INV_X1    g663(.A(new_n649), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n643), .A2(new_n865), .A3(new_n647), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n650), .A2(new_n866), .A3(KEYINPUT54), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n643), .B2(new_n647), .ZN(new_n868));
  XOR2_X1   g667(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n869));
  AOI21_X1  g668(.A(new_n656), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT55), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n659), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n867), .A2(KEYINPUT55), .A3(new_n870), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n612), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n586), .A2(new_n589), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n604), .B2(new_n587), .ZN(new_n877));
  INV_X1    g676(.A(new_n557), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n611), .A2(new_n660), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n734), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n874), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(new_n872), .A3(new_n871), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n611), .B(new_n879), .C1(new_n732), .C2(new_n700), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n864), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n611), .A2(new_n879), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n734), .A2(new_n888), .A3(new_n883), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n883), .A2(new_n612), .B1(new_n888), .B2(new_n660), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT115), .B(new_n889), .C1(new_n890), .C2(new_n734), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n891), .A3(new_n810), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n703), .A2(KEYINPUT113), .A3(new_n612), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT113), .B1(new_n703), .B2(new_n612), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n727), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n461), .A2(new_n443), .A3(new_n283), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n249), .A3(new_n613), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n461), .B1(new_n892), .B2(new_n895), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n900), .A2(new_n444), .A3(new_n481), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n612), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n899), .B1(new_n902), .B2(new_n249), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT116), .ZN(G1340gat));
  NOR3_X1   g703(.A1(new_n898), .A2(new_n251), .A3(new_n661), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n901), .A2(new_n660), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n251), .ZN(G1341gat));
  OR2_X1    g706(.A1(new_n239), .A2(new_n240), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n810), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n896), .A2(new_n684), .A3(new_n897), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n901), .A2(new_n909), .B1(new_n910), .B2(new_n908), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT117), .ZN(G1342gat));
  NAND3_X1  g711(.A1(new_n901), .A2(new_n243), .A3(new_n734), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n914));
  OAI21_X1  g713(.A(G134gat), .B1(new_n898), .B2(new_n733), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(G1343gat));
  XOR2_X1   g716(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n918));
  NAND2_X1  g717(.A1(new_n722), .A2(new_n785), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n443), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n900), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n612), .A2(new_n316), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT120), .Z(new_n924));
  AOI211_X1 g723(.A(KEYINPUT57), .B(new_n505), .C1(new_n892), .C2(new_n895), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n461), .A2(new_n443), .A3(new_n540), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n810), .B1(new_n881), .B2(new_n886), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n487), .B1(new_n927), .B2(new_n895), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT57), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n925), .A2(new_n613), .A3(new_n930), .ZN(new_n931));
  OAI221_X1 g730(.A(new_n918), .B1(new_n922), .B2(new_n924), .C1(new_n316), .C2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(new_n925), .B2(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n892), .A2(new_n895), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n929), .A3(new_n785), .ZN(new_n936));
  INV_X1    g735(.A(new_n926), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n927), .A2(new_n895), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n727), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n939), .B2(KEYINPUT57), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n940), .A3(KEYINPUT118), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n941), .A3(new_n612), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n942), .A2(new_n943), .A3(G141gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n942), .B2(G141gat), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n922), .A2(new_n924), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT58), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n932), .B1(new_n947), .B2(new_n948), .ZN(G1344gat));
  NAND3_X1  g748(.A1(new_n921), .A2(new_n314), .A3(new_n660), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n941), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI211_X1 g751(.A(KEYINPUT59), .B(new_n314), .C1(new_n952), .C2(new_n660), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n927), .B1(new_n612), .B2(new_n703), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n929), .A3(new_n727), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n505), .B1(new_n892), .B2(new_n895), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n929), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n957), .A2(new_n661), .ZN(new_n958));
  OAI21_X1  g757(.A(G148gat), .B1(new_n958), .B2(new_n937), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(KEYINPUT59), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n950), .B1(new_n953), .B2(new_n960), .ZN(G1345gat));
  OAI21_X1  g760(.A(G155gat), .B1(new_n951), .B2(new_n810), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n810), .A2(G155gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n922), .B2(new_n963), .ZN(G1346gat));
  NAND3_X1  g763(.A1(new_n952), .A2(KEYINPUT123), .A3(new_n734), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n966), .B1(new_n951), .B2(new_n733), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n965), .A2(G162gat), .A3(new_n967), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n922), .A2(G162gat), .A3(new_n733), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT122), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(G1347gat));
  AOI21_X1  g770(.A(new_n705), .B1(new_n892), .B2(new_n895), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n481), .A2(new_n443), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(G169gat), .B1(new_n975), .B2(new_n612), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n896), .A2(new_n461), .A3(new_n443), .A4(new_n284), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n977), .A2(new_n204), .A3(new_n613), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n976), .A2(new_n978), .ZN(G1348gat));
  OAI21_X1  g778(.A(G176gat), .B1(new_n977), .B2(new_n661), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n660), .A2(new_n205), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n974), .B2(new_n981), .ZN(G1349gat));
  OAI21_X1  g781(.A(G183gat), .B1(new_n977), .B2(new_n810), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n684), .A2(new_n224), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n974), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g785(.A(G190gat), .B1(new_n977), .B2(new_n733), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n987), .B(KEYINPUT61), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n975), .A2(new_n219), .A3(new_n734), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1351gat));
  NOR2_X1   g789(.A1(new_n919), .A2(new_n444), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n972), .A2(new_n991), .ZN(new_n992));
  OR3_X1    g791(.A1(new_n992), .A2(G197gat), .A3(new_n613), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n722), .A2(new_n461), .A3(new_n443), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n957), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(KEYINPUT124), .B1(new_n995), .B2(new_n613), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(G197gat), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n995), .A2(KEYINPUT124), .A3(new_n613), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n993), .B1(new_n997), .B2(new_n998), .ZN(G1352gat));
  XNOR2_X1  g798(.A(KEYINPUT125), .B(G204gat), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n992), .A2(new_n661), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1001), .B(KEYINPUT62), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1000), .B1(new_n958), .B2(new_n994), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1353gat));
  INV_X1    g803(.A(KEYINPUT63), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n286), .B1(KEYINPUT126), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1006), .B1(new_n995), .B2(new_n810), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT63), .ZN(new_n1009));
  OAI221_X1 g808(.A(new_n1006), .B1(KEYINPUT126), .B2(new_n1005), .C1(new_n995), .C2(new_n810), .ZN(new_n1010));
  INV_X1    g809(.A(new_n992), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1011), .A2(new_n286), .A3(new_n684), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(G1354gat));
  AOI21_X1  g812(.A(G218gat), .B1(new_n1011), .B2(new_n734), .ZN(new_n1014));
  XNOR2_X1  g813(.A(new_n995), .B(KEYINPUT127), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n733), .A2(new_n298), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(G1355gat));
endmodule


