//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(KEYINPUT24), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n203), .A2(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n210), .C1(KEYINPUT24), .C2(new_n202), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT25), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NOR3_X1   g012(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  INV_X1    g015(.A(G169gat), .ZN(new_n217));
  INV_X1    g016(.A(G176gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT27), .B(G183gat), .Z(new_n220));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n204), .A2(KEYINPUT27), .ZN(new_n223));
  AOI21_X1  g022(.A(G190gat), .B1(new_n223), .B2(KEYINPUT64), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT28), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT28), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n220), .A2(new_n226), .A3(G190gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n219), .B(new_n202), .C1(new_n225), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G226gat), .A2(G233gat), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n232), .A3(new_n230), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(G197gat), .A2(G204gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(G197gat), .A2(G204gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G218gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G211gat), .ZN(new_n239));
  INV_X1    g038(.A(G211gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G218gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243));
  OR2_X1    g042(.A1(KEYINPUT68), .A2(G211gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT68), .A2(G211gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(G218gat), .A3(new_n245), .ZN(new_n246));
  AOI211_X1 g045(.A(new_n237), .B(new_n242), .C1(new_n243), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n242), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n243), .ZN(new_n249));
  INV_X1    g048(.A(new_n237), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n234), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253));
  INV_X1    g052(.A(G64gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G92gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n247), .B2(new_n251), .ZN(new_n260));
  AND2_X1   g059(.A1(KEYINPUT68), .A2(G211gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(KEYINPUT68), .A2(G211gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT22), .B1(new_n263), .B2(G218gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n242), .B1(new_n264), .B2(new_n237), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(new_n248), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(KEYINPUT69), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n231), .A2(new_n268), .A3(new_n233), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n252), .A2(new_n258), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT30), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n269), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n257), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n270), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G127gat), .B(G134gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(KEYINPUT1), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G120gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(KEYINPUT1), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n281), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G141gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT73), .B1(new_n285), .B2(G148gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n287));
  INV_X1    g086(.A(G148gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(G141gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(new_n288), .A3(G141gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n285), .A2(KEYINPUT72), .A3(G148gat), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n286), .A2(new_n289), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT2), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  INV_X1    g095(.A(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n294), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n293), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n288), .A2(G141gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n285), .A2(G148gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n294), .ZN(new_n304));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT71), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(new_n298), .B2(new_n294), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n303), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n284), .B(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n281), .B(new_n283), .Z(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n309), .A3(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n316), .B2(new_n310), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n284), .A2(KEYINPUT4), .A3(new_n309), .A4(new_n300), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n321), .A2(new_n312), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n315), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT5), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT5), .B1(new_n313), .B2(new_n314), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n325), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT0), .B(G57gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(G85gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G1gat), .B(G29gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  NOR3_X1   g133(.A1(new_n330), .A2(KEYINPUT84), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT84), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n326), .A2(KEYINPUT5), .B1(new_n328), .B2(new_n325), .ZN(new_n337));
  INV_X1    g136(.A(new_n334), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(G225gat), .A3(G233gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n311), .A2(new_n312), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n342), .A2(KEYINPUT39), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(KEYINPUT39), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n344), .A2(new_n338), .A3(new_n345), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n346), .A2(KEYINPUT40), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(KEYINPUT40), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n278), .A2(new_n340), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n274), .A2(new_n258), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT37), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n234), .B2(new_n268), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n247), .A2(new_n251), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(new_n234), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n252), .A2(new_n353), .A3(new_n269), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n356), .A2(new_n351), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n352), .B1(new_n358), .B2(new_n258), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n337), .A2(KEYINPUT6), .A3(new_n338), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT76), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT6), .B1(new_n330), .B2(new_n334), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n335), .B2(new_n339), .ZN(new_n363));
  INV_X1    g162(.A(new_n357), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n353), .B1(new_n252), .B2(new_n269), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n350), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n359), .A2(new_n361), .A3(new_n363), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT83), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n265), .B2(new_n266), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n310), .B1(new_n369), .B2(KEYINPUT3), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n318), .A2(new_n232), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n260), .A3(new_n267), .ZN(new_n372));
  INV_X1    g171(.A(G228gat), .ZN(new_n373));
  INV_X1    g172(.A(G233gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n370), .A2(new_n372), .A3(KEYINPUT79), .A4(new_n375), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n370), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n371), .A2(new_n355), .ZN(new_n383));
  OAI211_X1 g182(.A(KEYINPUT77), .B(new_n310), .C1(new_n369), .C2(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n375), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT78), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n380), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G22gat), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT81), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n379), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n385), .A2(new_n389), .A3(new_n386), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n389), .B1(new_n385), .B2(new_n386), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(G22gat), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n392), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT80), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n388), .A2(new_n390), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n392), .A4(new_n394), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n393), .A2(new_n399), .A3(new_n401), .A4(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(G78gat), .B(G106gat), .Z(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT31), .ZN(new_n407));
  INV_X1    g206(.A(G50gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n392), .A2(KEYINPUT82), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n412), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n368), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  AOI211_X1 g217(.A(KEYINPUT83), .B(new_n416), .C1(new_n405), .C2(new_n410), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n349), .B(new_n367), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n391), .A2(KEYINPUT81), .A3(new_n392), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n398), .B1(new_n397), .B2(G22gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n401), .A2(new_n404), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n409), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT83), .B1(new_n425), .B2(new_n416), .ZN(new_n426));
  INV_X1    g225(.A(new_n278), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT75), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n428), .B(new_n429), .C1(new_n337), .C2(new_n338), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n334), .B2(new_n330), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n362), .A2(new_n428), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n360), .B(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n427), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n411), .A2(new_n368), .A3(new_n417), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT36), .ZN(new_n439));
  NAND2_X1  g238(.A1(G227gat), .A2(G233gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT67), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n229), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n316), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n316), .B1(new_n229), .B2(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT32), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT34), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n442), .B2(new_n316), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n450), .B2(new_n440), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n450), .A2(new_n449), .A3(new_n440), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n443), .A2(new_n440), .A3(new_n445), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT34), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n449), .A3(new_n440), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n455), .B(new_n456), .C1(new_n447), .C2(new_n446), .ZN(new_n457));
  XNOR2_X1  g256(.A(G15gat), .B(G43gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n446), .B2(KEYINPUT33), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n453), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n453), .B2(new_n457), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n439), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n453), .A2(new_n457), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n461), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n453), .A2(new_n457), .A3(new_n462), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(KEYINPUT36), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n420), .A2(new_n438), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n278), .B1(new_n361), .B2(new_n363), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n472), .B(new_n473), .C1(new_n418), .C2(new_n419), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT35), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n426), .A2(new_n437), .ZN(new_n477));
  INV_X1    g276(.A(new_n436), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(KEYINPUT35), .A3(new_n472), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n471), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT88), .B(G36gat), .ZN(new_n482));
  INV_X1    g281(.A(G29gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G36gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT14), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n483), .A2(new_n485), .B1(new_n486), .B2(KEYINPUT86), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(KEYINPUT86), .B2(new_n486), .ZN(new_n488));
  OR4_X1    g287(.A1(KEYINPUT86), .A2(new_n486), .A3(G29gat), .A4(G36gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT87), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n484), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(KEYINPUT87), .A3(new_n489), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G43gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G50gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n408), .A2(G43gat), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT15), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT89), .B(G50gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n495), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT15), .B1(new_n501), .B2(new_n497), .ZN(new_n502));
  NOR4_X1   g301(.A1(new_n502), .A2(new_n490), .A3(new_n498), .A4(new_n484), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT16), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(G1gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(G1gat), .B2(new_n506), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n509), .B(G8gat), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT93), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n511), .ZN(new_n513));
  INV_X1    g312(.A(new_n498), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n492), .B2(new_n493), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(new_n503), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n510), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n512), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT92), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT13), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT18), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n499), .A2(new_n504), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT17), .B1(new_n515), .B2(new_n503), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n510), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT90), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n526), .A2(KEYINPUT18), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n535), .A3(new_n510), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n533), .A2(new_n513), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n520), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n527), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n531), .B2(new_n510), .ZN(new_n540));
  AOI211_X1 g339(.A(KEYINPUT90), .B(new_n511), .C1(new_n529), .C2(new_n530), .ZN(new_n541));
  INV_X1    g340(.A(new_n513), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(new_n526), .A3(KEYINPUT18), .A4(new_n520), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT11), .B(G169gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G197gat), .ZN(new_n547));
  XOR2_X1   g346(.A(G113gat), .B(G141gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT12), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n525), .A2(new_n539), .A3(new_n544), .A4(new_n550), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n480), .A2(new_n481), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n481), .B1(new_n480), .B2(new_n554), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G57gat), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT96), .B1(new_n558), .B2(G64gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(new_n254), .A3(G57gat), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n559), .B(new_n561), .C1(G57gat), .C2(new_n254), .ZN(new_n562));
  NAND2_X1  g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  OR2_X1    g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT98), .ZN(new_n570));
  XNOR2_X1  g369(.A(G57gat), .B(G64gat), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n563), .B(new_n564), .C1(new_n571), .C2(new_n565), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n570), .B1(new_n569), .B2(new_n572), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n510), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G183gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(new_n240), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n585), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n581), .A2(new_n582), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n576), .A2(new_n577), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT104), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT105), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT100), .ZN(new_n601));
  INV_X1    g400(.A(G85gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n601), .A2(KEYINPUT8), .B1(new_n602), .B2(new_n256), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(G85gat), .A3(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G99gat), .B(G106gat), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610));
  INV_X1    g409(.A(new_n608), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n603), .A2(new_n611), .A3(new_n606), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(KEYINPUT101), .A3(new_n608), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n531), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT102), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n531), .A2(new_n618), .A3(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n597), .A2(KEYINPUT105), .ZN(new_n621));
  NAND3_X1  g420(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n622), .B1(new_n615), .B2(new_n516), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT103), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n625), .B(new_n622), .C1(new_n615), .C2(new_n516), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n620), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n620), .A2(new_n631), .A3(new_n627), .A4(new_n621), .ZN(new_n632));
  XOR2_X1   g431(.A(G134gat), .B(G162gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n630), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n634), .B1(new_n630), .B2(new_n632), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n599), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n630), .A2(new_n632), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n633), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n598), .A3(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n569), .A2(new_n572), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n646), .A2(new_n573), .A3(new_n613), .A4(new_n614), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n569), .A2(new_n609), .A3(new_n572), .A4(new_n612), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n613), .A2(new_n614), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n651), .B(KEYINPUT10), .C1(new_n574), .C2(new_n575), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n653), .B1(new_n650), .B2(new_n652), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n644), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n647), .A2(new_n649), .ZN(new_n657));
  INV_X1    g456(.A(new_n644), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT107), .ZN(new_n662));
  INV_X1    g461(.A(G120gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n656), .A2(new_n659), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n659), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n658), .B1(new_n650), .B2(new_n652), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n594), .A2(new_n643), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n557), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n433), .A2(new_n435), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  INV_X1    g475(.A(new_n557), .ZN(new_n677));
  INV_X1    g476(.A(new_n672), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(new_n278), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n681));
  OR2_X1    g480(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n680), .A2(KEYINPUT42), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(G8gat), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n673), .A2(new_n278), .A3(new_n681), .A4(new_n682), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(G1325gat));
  AOI21_X1  g487(.A(G15gat), .B1(new_n673), .B2(new_n472), .ZN(new_n689));
  INV_X1    g488(.A(new_n470), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G15gat), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT108), .Z(new_n692));
  AOI21_X1  g491(.A(new_n689), .B1(new_n673), .B2(new_n692), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n418), .A2(new_n419), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n673), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  NOR2_X1   g496(.A1(new_n594), .A2(new_n670), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n642), .B(new_n698), .C1(new_n555), .C2(new_n556), .ZN(new_n699));
  INV_X1    g498(.A(new_n674), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n699), .A2(G29gat), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT45), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n480), .A2(KEYINPUT44), .A3(new_n642), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n480), .B2(new_n642), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n554), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n594), .A2(new_n707), .A3(new_n670), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n674), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n703), .B1(new_n709), .B2(G29gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n702), .B1(new_n701), .B2(new_n710), .ZN(G1328gat));
  INV_X1    g510(.A(new_n482), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n699), .A2(new_n712), .A3(new_n427), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n706), .A2(new_n278), .A3(new_n708), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n712), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n714), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(G1329gat));
  NAND2_X1  g518(.A1(new_n472), .A2(new_n495), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n699), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n480), .A2(new_n642), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n480), .A2(KEYINPUT44), .A3(new_n642), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n725), .A2(new_n690), .A3(new_n708), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT111), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G43gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n727), .A2(KEYINPUT111), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n722), .B(KEYINPUT47), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n727), .A2(KEYINPUT110), .A3(G43gat), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT110), .B1(new_n727), .B2(G43gat), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n732), .A2(new_n733), .A3(new_n721), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n735));
  OAI21_X1  g534(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(G1330gat));
  NAND4_X1  g535(.A1(new_n706), .A2(KEYINPUT113), .A3(new_n694), .A4(new_n708), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n725), .A2(new_n694), .A3(new_n708), .A4(new_n726), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n740), .A3(new_n500), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n477), .A2(new_n500), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n699), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT112), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(KEYINPUT112), .B2(KEYINPUT48), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n738), .A2(new_n747), .A3(new_n500), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n745), .A2(KEYINPUT48), .B1(new_n746), .B2(new_n748), .ZN(G1331gat));
  AND2_X1   g548(.A1(new_n480), .A2(new_n670), .ZN(new_n750));
  INV_X1    g549(.A(new_n594), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(new_n554), .A3(new_n642), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n700), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n558), .ZN(G1332gat));
  INV_X1    g554(.A(new_n753), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n278), .B(KEYINPUT114), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT49), .B(G64gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n753), .A2(new_n757), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT115), .B(KEYINPUT116), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1333gat));
  NAND3_X1  g563(.A1(new_n756), .A2(G71gat), .A3(new_n690), .ZN(new_n765));
  INV_X1    g564(.A(new_n472), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n753), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(G71gat), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n756), .A2(new_n694), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g570(.A1(new_n594), .A2(new_n554), .A3(new_n671), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n706), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n773), .A2(new_n602), .A3(new_n700), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n594), .A2(new_n554), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n480), .A2(new_n642), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT51), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n480), .A2(new_n778), .A3(new_n642), .A4(new_n775), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n674), .A3(new_n670), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n774), .B1(new_n602), .B2(new_n781), .ZN(G1336gat));
  AND2_X1   g581(.A1(new_n706), .A2(new_n772), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n256), .B1(new_n783), .B2(new_n278), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n777), .A2(new_n670), .A3(new_n758), .A4(new_n779), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT52), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(KEYINPUT52), .ZN(new_n788));
  OAI21_X1  g587(.A(G92gat), .B1(new_n773), .B2(new_n757), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n773), .B2(new_n470), .ZN(new_n792));
  INV_X1    g591(.A(G99gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n780), .A2(new_n793), .A3(new_n670), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n766), .B2(new_n794), .ZN(G1338gat));
  NAND4_X1  g594(.A1(new_n725), .A2(new_n694), .A3(new_n726), .A4(new_n772), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(new_n797), .A3(G106gat), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n477), .A2(G106gat), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n777), .A2(new_n670), .A3(new_n779), .A4(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n798), .B(new_n800), .C1(KEYINPUT118), .C2(new_n797), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n796), .A2(new_n802), .A3(G106gat), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n800), .A2(KEYINPUT118), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n796), .B2(G106gat), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n801), .B1(new_n806), .B2(new_n797), .ZN(G1339gat));
  NAND3_X1  g606(.A1(new_n650), .A2(new_n658), .A3(new_n652), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n656), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n665), .B1(new_n668), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT119), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n811), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(new_n666), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n812), .A2(new_n818), .A3(new_n813), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n815), .A2(new_n817), .A3(new_n554), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n543), .A2(new_n520), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n519), .A2(new_n522), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n549), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n553), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n670), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n642), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n636), .A2(new_n637), .A3(new_n599), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n598), .B1(new_n640), .B2(new_n635), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n817), .A3(new_n819), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n751), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n594), .A2(new_n707), .A3(new_n643), .A4(new_n671), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n694), .A2(new_n766), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n835), .A2(new_n674), .A3(new_n836), .A4(new_n757), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(G113gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n839), .A3(new_n554), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n700), .B1(new_n833), .B2(new_n834), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(KEYINPUT120), .A3(new_n836), .A4(new_n757), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n554), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n841), .B1(new_n847), .B2(G113gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n837), .A2(new_n842), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n707), .B1(new_n849), .B2(new_n845), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(KEYINPUT121), .A3(new_n839), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n840), .B1(new_n848), .B2(new_n851), .ZN(G1340gat));
  NOR2_X1   g651(.A1(new_n843), .A2(new_n846), .ZN(new_n853));
  OAI21_X1  g652(.A(G120gat), .B1(new_n853), .B2(new_n671), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n663), .A3(new_n670), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1341gat));
  AOI21_X1  g655(.A(G127gat), .B1(new_n838), .B2(new_n594), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n853), .A2(new_n751), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(G127gat), .ZN(G1342gat));
  OAI21_X1  g658(.A(G134gat), .B1(new_n853), .B2(new_n643), .ZN(new_n860));
  INV_X1    g659(.A(G134gat), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n643), .A2(new_n278), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n844), .A2(new_n861), .A3(new_n836), .A4(new_n862), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT56), .Z(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(G1343gat));
  NOR3_X1   g664(.A1(new_n690), .A2(new_n700), .A3(new_n758), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT122), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n835), .A2(new_n694), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n817), .A2(new_n554), .A3(new_n814), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n642), .B1(new_n872), .B2(new_n826), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n751), .B1(new_n832), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n477), .B1(new_n874), .B2(new_n834), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT57), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n867), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n285), .B1(new_n877), .B2(new_n554), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n477), .B1(new_n833), .B2(new_n834), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n866), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(G141gat), .A3(new_n707), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT58), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n867), .ZN(new_n883));
  INV_X1    g682(.A(new_n876), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n879), .A2(new_n869), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886), .B2(new_n707), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  INV_X1    g687(.A(new_n881), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n882), .A2(new_n890), .ZN(G1344gat));
  OAI22_X1  g690(.A1(new_n868), .A2(new_n870), .B1(new_n875), .B2(KEYINPUT57), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n670), .A3(new_n883), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n895), .A3(new_n670), .ZN(new_n896));
  INV_X1    g695(.A(new_n880), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n670), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n894), .B(new_n896), .C1(G148gat), .C2(new_n898), .ZN(G1345gat));
  AOI21_X1  g698(.A(G155gat), .B1(new_n897), .B2(new_n594), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n751), .A2(new_n296), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n877), .B2(new_n901), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n886), .B2(new_n643), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n690), .A2(new_n700), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n879), .A2(new_n297), .A3(new_n862), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1347gat));
  AOI211_X1 g705(.A(new_n674), .B(new_n757), .C1(new_n833), .C2(new_n834), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n836), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n217), .A3(new_n554), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n674), .B1(new_n833), .B2(new_n834), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n836), .A2(new_n278), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n707), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n910), .A2(new_n915), .ZN(G1348gat));
  NOR3_X1   g715(.A1(new_n914), .A2(new_n218), .A3(new_n671), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n218), .B1(new_n908), .B2(new_n671), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n918), .A2(KEYINPUT124), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(KEYINPUT124), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1349gat));
  NAND4_X1  g720(.A1(new_n835), .A2(new_n700), .A3(new_n594), .A4(new_n913), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G183gat), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n751), .A2(new_n220), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n911), .A2(new_n836), .A3(new_n758), .A4(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n924), .B1(new_n923), .B2(new_n926), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n923), .A2(new_n926), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT126), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n933), .A2(new_n927), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n931), .A2(new_n934), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n909), .A2(new_n205), .A3(new_n642), .ZN(new_n936));
  OAI21_X1  g735(.A(G190gat), .B1(new_n914), .B2(new_n643), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1351gat));
  NOR3_X1   g739(.A1(new_n690), .A2(new_n674), .A3(new_n427), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n892), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n554), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G197gat), .ZN(new_n944));
  AND4_X1   g743(.A1(new_n694), .A2(new_n911), .A3(new_n470), .A4(new_n758), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(G197gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n707), .B2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(G204gat), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n907), .A2(new_n949), .A3(new_n694), .A4(new_n470), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT62), .B1(new_n950), .B2(new_n671), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n945), .A2(new_n952), .A3(new_n949), .A4(new_n670), .ZN(new_n953));
  AOI211_X1 g752(.A(new_n477), .B(new_n870), .C1(new_n833), .C2(new_n834), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n872), .A2(new_n826), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n818), .B1(new_n812), .B2(new_n813), .ZN(new_n956));
  AOI211_X1 g755(.A(KEYINPUT119), .B(KEYINPUT55), .C1(new_n809), .C2(new_n811), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n816), .A2(new_n666), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n824), .B1(new_n638), .B2(new_n641), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n955), .A2(new_n643), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n834), .B1(new_n961), .B2(new_n594), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT57), .B1(new_n962), .B2(new_n694), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n670), .B(new_n941), .C1(new_n954), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G204gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n951), .A2(new_n953), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n951), .A2(new_n953), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n892), .A2(new_n594), .A3(new_n941), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n594), .B1(new_n262), .B2(new_n261), .ZN(new_n974));
  OAI22_X1  g773(.A1(new_n972), .A2(new_n973), .B1(new_n946), .B2(new_n974), .ZN(G1354gat));
  NAND3_X1  g774(.A1(new_n945), .A2(new_n238), .A3(new_n642), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n942), .A2(new_n642), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n977), .B2(new_n238), .ZN(G1355gat));
endmodule


