//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT68), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G221), .A3(G218), .A4(G220), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n467), .A2(new_n474), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n467), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n474), .B2(G112), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n478), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT69), .Z(G162));
  NAND4_X1  g059(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n474), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n474), .A2(G2104), .ZN(new_n487));
  INV_X1    g062(.A(G102), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n467), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n489), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(G75), .A2(G543), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g073(.A(G543), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT73), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n496), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT75), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI211_X1 g085(.A(KEYINPUT70), .B(KEYINPUT6), .C1(new_n510), .C2(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n515), .B2(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n505), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT74), .B(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n517), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G50), .A3(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n509), .A2(new_n520), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n518), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n517), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g105(.A(KEYINPUT76), .B(new_n511), .C1(new_n514), .C2(new_n516), .ZN(new_n531));
  AND4_X1   g106(.A1(G51), .A2(new_n530), .A3(G543), .A4(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G63), .ZN(new_n533));
  NOR3_X1   g108(.A1(new_n505), .A2(new_n533), .A3(new_n510), .ZN(new_n534));
  OAI21_X1  g109(.A(KEYINPUT77), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n505), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G63), .A3(G651), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n530), .A2(G51), .A3(G543), .A4(new_n531), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n528), .B1(new_n535), .B2(new_n540), .ZN(G168));
  NAND4_X1  g116(.A1(new_n530), .A2(G52), .A3(G543), .A4(new_n531), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n521), .A2(new_n502), .A3(new_n500), .A4(new_n504), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n500), .A2(G64), .A3(new_n502), .A4(new_n504), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n510), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n536), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n510), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n530), .A2(G543), .A3(new_n531), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n552), .A2(new_n553), .B1(new_n543), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT78), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n505), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n518), .B2(G91), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n530), .A2(G543), .A3(new_n531), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .A3(G53), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n530), .A2(G53), .A3(G543), .A4(new_n531), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n569), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n574), .B1(new_n545), .B2(new_n548), .ZN(new_n575));
  INV_X1    g150(.A(new_n548), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n536), .A2(G90), .A3(new_n521), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n576), .A2(KEYINPUT79), .A3(new_n542), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  NAND2_X1  g155(.A1(new_n568), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n536), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n518), .A2(G87), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n505), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n500), .A2(G86), .A3(new_n502), .A4(new_n504), .ZN(new_n589));
  NAND2_X1  g164(.A1(G48), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(new_n521), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n510), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n518), .A2(G85), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT80), .B(G47), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n568), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n568), .A2(G54), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT10), .B1(new_n543), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n505), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n518), .A2(new_n608), .A3(G92), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n601), .A2(new_n603), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n600), .B1(G868), .B2(new_n611), .ZN(G284));
  OAI21_X1  g187(.A(new_n600), .B1(G868), .B2(new_n611), .ZN(G321));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT81), .B1(new_n614), .B2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  MUX2_X1   g191(.A(KEYINPUT81), .B(new_n615), .S(new_n616), .Z(G297));
  MUX2_X1   g192(.A(KEYINPUT81), .B(new_n615), .S(new_n616), .Z(G280));
  XOR2_X1   g193(.A(KEYINPUT82), .B(G559), .Z(new_n619));
  OAI21_X1  g194(.A(new_n611), .B1(G860), .B2(new_n619), .ZN(G148));
  NAND2_X1  g195(.A1(new_n611), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g199(.A1(new_n467), .A2(new_n487), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT84), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n477), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n479), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n630), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2435), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2438), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  AOI21_X1  g233(.A(KEYINPUT18), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(KEYINPUT18), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n659), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n663), .B(new_n666), .Z(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT88), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT90), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n670), .A2(new_n674), .A3(new_n677), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT22), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  XNOR2_X1  g263(.A(KEYINPUT31), .B(G11), .ZN(new_n689));
  NAND2_X1  g264(.A1(G171), .A2(G16), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G5), .B2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G1961), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT97), .ZN(new_n695));
  OR2_X1    g270(.A1(G29), .A2(G32), .ZN(new_n696));
  AOI22_X1  g271(.A1(G129), .A2(new_n477), .B1(new_n479), .B2(G141), .ZN(new_n697));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT26), .Z(new_n699));
  INV_X1    g274(.A(G105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n697), .B(new_n699), .C1(new_n700), .C2(new_n487), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n696), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT27), .B(G1996), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n694), .A2(new_n695), .B1(KEYINPUT95), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(KEYINPUT95), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n691), .A2(new_n692), .ZN(new_n708));
  NOR2_X1   g283(.A1(G29), .A2(G35), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G162), .B2(G29), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT29), .ZN(new_n711));
  OAI221_X1 g286(.A(new_n708), .B1(new_n694), .B2(new_n695), .C1(new_n711), .C2(G2090), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n635), .A2(new_n702), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n703), .A2(new_n704), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT30), .B(G28), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n713), .B(new_n715), .C1(new_n702), .C2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G34), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(KEYINPUT24), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(KEYINPUT24), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n702), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G160), .B2(new_n702), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G2084), .Z(new_n723));
  AND2_X1   g298(.A1(new_n702), .A2(G33), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n479), .A2(G139), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT25), .Z(new_n727));
  INV_X1    g302(.A(new_n467), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n728), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n725), .B(new_n727), .C1(new_n729), .C2(new_n474), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(G29), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(G2072), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n717), .A2(new_n723), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n707), .A2(new_n712), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G19), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n556), .B2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G1341), .Z(new_n740));
  AND2_X1   g315(.A1(new_n702), .A2(G26), .ZN(new_n741));
  OAI21_X1  g316(.A(G2104), .B1(new_n474), .B2(G116), .ZN(new_n742));
  INV_X1    g317(.A(G104), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n474), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT93), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n477), .A2(G128), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n479), .A2(G140), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(G29), .ZN(new_n749));
  MUX2_X1   g324(.A(new_n741), .B(new_n749), .S(KEYINPUT28), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2067), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n737), .A2(G4), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n611), .B2(new_n737), .ZN(new_n753));
  INV_X1    g328(.A(G1348), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n740), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT94), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT23), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n737), .A2(G20), .ZN(new_n759));
  AOI22_X1  g334(.A1(G299), .A2(G16), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n758), .B2(new_n759), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G1956), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n711), .A2(G2090), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT98), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n756), .A2(KEYINPUT94), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n736), .A2(new_n757), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(KEYINPUT96), .B1(G16), .B2(G21), .ZN(new_n769));
  NAND2_X1  g344(.A1(G168), .A2(G16), .ZN(new_n770));
  MUX2_X1   g345(.A(KEYINPUT96), .B(new_n769), .S(new_n770), .Z(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G1966), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(G1966), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n764), .B2(new_n765), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n768), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n737), .A2(G22), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G166), .B2(new_n737), .ZN(new_n778));
  INV_X1    g353(.A(G1971), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G6), .B(G305), .S(G16), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT91), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT32), .B(G1981), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n785));
  NOR2_X1   g360(.A1(G16), .A2(G23), .ZN(new_n786));
  INV_X1    g361(.A(G288), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n780), .A2(new_n784), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n702), .A2(G25), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n477), .A2(G119), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n479), .A2(G131), .ZN(new_n794));
  OR2_X1    g369(.A1(G95), .A2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n792), .B1(new_n798), .B2(new_n702), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT35), .B(G1991), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n799), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n737), .A2(G24), .ZN(new_n803));
  INV_X1    g378(.A(G290), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n737), .ZN(new_n805));
  INV_X1    g380(.A(G1986), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n791), .A2(new_n802), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT92), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n791), .A2(KEYINPUT92), .A3(new_n802), .A4(new_n807), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n780), .A2(new_n784), .A3(new_n790), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n813), .B1(new_n812), .B2(new_n815), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n689), .B(new_n776), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n702), .A2(G27), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G164), .B2(new_n702), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2078), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(G311));
  OR2_X1    g397(.A1(new_n816), .A2(new_n817), .ZN(new_n823));
  INV_X1    g398(.A(new_n821), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n823), .A2(new_n689), .A3(new_n776), .A4(new_n824), .ZN(G150));
  NAND2_X1  g400(.A1(new_n536), .A2(G67), .ZN(new_n826));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n510), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G55), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n552), .A2(new_n829), .B1(new_n543), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT37), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n556), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n828), .A2(new_n831), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n551), .B2(new_n555), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n611), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n834), .B1(new_n842), .B2(G860), .ZN(G145));
  XNOR2_X1  g418(.A(G160), .B(new_n635), .ZN(new_n844));
  XNOR2_X1  g419(.A(G162), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n748), .B(new_n494), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n730), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n701), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n477), .A2(G130), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n479), .A2(G142), .ZN(new_n850));
  NOR2_X1   g425(.A1(G106), .A2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(new_n474), .B2(G118), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n626), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n797), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT99), .B1(new_n848), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n848), .B(new_n855), .ZN(new_n857));
  AOI211_X1 g432(.A(new_n845), .B(new_n856), .C1(new_n857), .C2(KEYINPUT99), .ZN(new_n858));
  AOI211_X1 g433(.A(G37), .B(new_n858), .C1(new_n845), .C2(new_n857), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(G395));
  XNOR2_X1  g436(.A(G290), .B(new_n787), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(G303), .B(G305), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n863), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT42), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n603), .A2(new_n609), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n570), .B(KEYINPUT9), .ZN(new_n871));
  AOI22_X1  g446(.A1(G54), .A2(new_n568), .B1(new_n606), .B2(G651), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n567), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(G299), .A2(new_n610), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(KEYINPUT41), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n873), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(KEYINPUT100), .A3(new_n879), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n838), .B(new_n621), .ZN(new_n884));
  MUX2_X1   g459(.A(new_n876), .B(new_n883), .S(new_n884), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n869), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(G868), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(G868), .B2(new_n836), .ZN(G295));
  OAI21_X1  g463(.A(new_n887), .B1(G868), .B2(new_n836), .ZN(G331));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n890));
  NAND2_X1  g465(.A1(G301), .A2(G168), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n892));
  NAND2_X1  g467(.A1(G286), .A2(G171), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  NAND3_X1  g469(.A1(G301), .A2(G168), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n838), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n835), .A2(new_n837), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n898), .A2(new_n892), .A3(new_n893), .A4(new_n895), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(KEYINPUT103), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n901), .A3(new_n838), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n883), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n897), .A2(new_n876), .A3(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT104), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n897), .A2(new_n906), .A3(new_n876), .A4(new_n899), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n868), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n890), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI211_X1 g486(.A(KEYINPUT105), .B(G37), .C1(new_n908), .C2(new_n868), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n908), .A2(new_n868), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT43), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n875), .B1(new_n900), .B2(new_n902), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n897), .A2(new_n899), .B1(new_n880), .B2(new_n877), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n868), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND4_X1   g493(.A1(KEYINPUT43), .A2(new_n914), .A3(new_n910), .A4(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT44), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n913), .B2(new_n914), .ZN(new_n923));
  AND4_X1   g498(.A1(new_n922), .A2(new_n914), .A3(new_n910), .A4(new_n918), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n925), .ZN(G397));
  INV_X1    g501(.A(KEYINPUT125), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n787), .A2(G1976), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT52), .ZN(new_n929));
  AOI21_X1  g504(.A(G1384), .B1(new_n486), .B2(new_n493), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n470), .A2(new_n475), .A3(G40), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n932), .A2(G8), .ZN(new_n933));
  INV_X1    g508(.A(G1976), .ZN(new_n934));
  NAND2_X1  g509(.A1(G288), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n928), .A2(new_n929), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n933), .B1(new_n934), .B2(G288), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT52), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n937), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(G305), .A2(G1981), .ZN(new_n943));
  INV_X1    g518(.A(G1981), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n588), .A2(new_n592), .A3(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(KEYINPUT111), .A2(KEYINPUT49), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(KEYINPUT111), .A2(KEYINPUT49), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n943), .A2(KEYINPUT111), .A3(KEYINPUT49), .A4(new_n945), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n933), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n949), .A2(KEYINPUT112), .A3(new_n933), .A4(new_n950), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n942), .A2(new_n955), .A3(KEYINPUT113), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT113), .B1(new_n942), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n931), .B1(new_n930), .B2(KEYINPUT45), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT106), .B(G1384), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n779), .ZN(new_n963));
  INV_X1    g538(.A(new_n931), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(new_n965), .B2(new_n930), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n494), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT50), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n963), .B1(G2090), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G8), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(G303), .B2(G8), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(G303), .A2(G8), .A3(new_n973), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n969), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n930), .A2(new_n965), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT107), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n966), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n963), .B1(G2090), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n963), .B(KEYINPUT108), .C1(G2090), .C2(new_n982), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(G8), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n976), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(new_n974), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n977), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n956), .A2(new_n957), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n982), .A2(KEYINPUT117), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n979), .A2(new_n966), .A3(new_n981), .A4(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT122), .B(G1961), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n962), .B2(G2078), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n958), .B1(KEYINPUT45), .B2(new_n930), .ZN(new_n999));
  INV_X1    g574(.A(G2078), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(KEYINPUT53), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G301), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n494), .A2(new_n960), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1008));
  NAND2_X1  g583(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n997), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1007), .A2(new_n931), .A3(new_n961), .A4(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n996), .A2(G301), .A3(new_n998), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1004), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT124), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n982), .A2(G2084), .B1(new_n999), .B2(G1966), .ZN(new_n1018));
  AND2_X1   g593(.A1(G286), .A2(G8), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1023), .B(G8), .C1(new_n1018), .C2(G286), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1018), .A2(G8), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1019), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(KEYINPUT51), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1013), .A2(KEYINPUT124), .A3(new_n1014), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n991), .A2(new_n1017), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n996), .A2(new_n998), .A3(new_n1011), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G171), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(KEYINPUT54), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n927), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1017), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(KEYINPUT125), .A3(new_n1034), .A4(new_n991), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT116), .B(G2072), .Z(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT56), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n959), .A2(new_n961), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1956), .B1(new_n966), .B2(new_n969), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G299), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT61), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(new_n1056), .A3(new_n1053), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n992), .A2(new_n754), .A3(new_n994), .ZN(new_n1059));
  INV_X1    g634(.A(new_n932), .ZN(new_n1060));
  INV_X1    g635(.A(G2067), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g638(.A1(new_n1063), .A2(KEYINPUT60), .B1(KEYINPUT120), .B2(new_n611), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(KEYINPUT60), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(new_n610), .B(KEYINPUT120), .Z(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT58), .B(G1341), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n962), .A2(G1996), .B1(new_n1060), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n556), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1072), .A2(KEYINPUT119), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(KEYINPUT119), .ZN(new_n1075));
  OR3_X1    g650(.A1(new_n1071), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1058), .A2(new_n1068), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1053), .B1(new_n1063), .B2(new_n610), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1052), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT118), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1036), .A2(new_n1038), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT63), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1025), .A2(G286), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n991), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n987), .A2(new_n989), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n955), .A3(new_n942), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n987), .A2(new_n989), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(new_n955), .A3(new_n942), .A4(new_n1084), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n955), .A2(new_n934), .A3(new_n787), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n945), .ZN(new_n1091));
  AOI22_X1  g666(.A1(KEYINPUT63), .A2(new_n1089), .B1(new_n1091), .B2(new_n933), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1085), .A2(new_n1087), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n956), .A2(new_n957), .ZN(new_n1094));
  INV_X1    g669(.A(new_n990), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1022), .A2(new_n1024), .A3(new_n1096), .A4(new_n1027), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1004), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n991), .A2(new_n1100), .A3(new_n1097), .A4(new_n1101), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT126), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1093), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1082), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n748), .B(new_n1061), .ZN(new_n1107));
  INV_X1    g682(.A(G1996), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n701), .B(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n797), .A2(new_n800), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n798), .A2(new_n801), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n804), .A2(new_n806), .ZN(new_n1114));
  NAND2_X1  g689(.A1(G290), .A2(G1986), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1007), .A2(new_n964), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1106), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1117), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1121), .B(KEYINPUT48), .Z(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1120), .B2(new_n1113), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1107), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1117), .B1(new_n1124), .B2(new_n701), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT46), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1120), .B2(G1996), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1117), .A2(KEYINPUT46), .A3(new_n1108), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT47), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1111), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1110), .A2(new_n1131), .B1(G2067), .B2(new_n748), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1117), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1123), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT127), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1119), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g711(.A1(new_n909), .A2(new_n910), .ZN(new_n1138));
  NAND2_X1  g712(.A1(new_n1138), .A2(KEYINPUT105), .ZN(new_n1139));
  NAND3_X1  g713(.A1(new_n909), .A2(new_n890), .A3(new_n910), .ZN(new_n1140));
  NAND3_X1  g714(.A1(new_n1139), .A2(new_n914), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g715(.A(new_n924), .B1(new_n1141), .B2(KEYINPUT43), .ZN(new_n1142));
  NOR2_X1   g716(.A1(G229), .A2(new_n460), .ZN(new_n1143));
  INV_X1    g717(.A(new_n1143), .ZN(new_n1144));
  OR2_X1    g718(.A1(G401), .A2(G227), .ZN(new_n1145));
  NOR4_X1   g719(.A1(new_n1142), .A2(new_n859), .A3(new_n1144), .A4(new_n1145), .ZN(G308));
  NOR2_X1   g720(.A1(new_n859), .A2(new_n1145), .ZN(new_n1147));
  OAI211_X1 g721(.A(new_n1147), .B(new_n1143), .C1(new_n923), .C2(new_n924), .ZN(G225));
endmodule


