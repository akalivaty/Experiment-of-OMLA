//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n534, new_n536, new_n537,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n595,
    new_n598, new_n600, new_n601, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n458), .A2(G2105), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n462), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT68), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(G136), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(G162));
  NAND4_X1  g053(.A1(new_n459), .A2(new_n461), .A3(G138), .A4(new_n471), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  OR2_X1    g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(KEYINPUT4), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n471), .A2(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  OR3_X1    g063(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n486), .B2(new_n487), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n489), .A2(new_n490), .B1(new_n472), .B2(G126), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n483), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  AND2_X1   g068(.A1(KEYINPUT5), .A2(G543), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G62), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(G651), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  XOR2_X1   g076(.A(KEYINPUT6), .B(G651), .Z(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(new_n496), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G88), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(G50), .A3(G543), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(G303));
  INV_X1    g082(.A(G303), .ZN(G166));
  NAND3_X1  g083(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT7), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G51), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n505), .A2(G89), .ZN(new_n514));
  NAND2_X1  g089(.A1(G63), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n496), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(G168));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n505), .ZN(new_n519));
  INV_X1    g094(.A(G90), .ZN(new_n520));
  INV_X1    g095(.A(G52), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n519), .A2(new_n520), .B1(new_n511), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(G171));
  INV_X1    g101(.A(G81), .ZN(new_n527));
  INV_X1    g102(.A(G43), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n519), .A2(new_n527), .B1(new_n511), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n524), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G860), .ZN(G153));
  AND3_X1   g108(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G36), .ZN(G176));
  NAND2_X1  g110(.A1(G1), .A2(G3), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT8), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(new_n537), .ZN(G188));
  INV_X1    g113(.A(G53), .ZN(new_n539));
  OR3_X1    g114(.A1(new_n511), .A2(KEYINPUT9), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(KEYINPUT9), .B1(new_n511), .B2(new_n539), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n503), .A2(G91), .ZN(new_n543));
  NAND2_X1  g118(.A1(G78), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G65), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n496), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(G651), .B1(new_n546), .B2(new_n547), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n542), .B(new_n543), .C1(new_n548), .C2(new_n549), .ZN(G299));
  INV_X1    g125(.A(G171), .ZN(G301));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n552));
  XNOR2_X1  g127(.A(G168), .B(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(G286));
  OAI21_X1  g129(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n518), .A2(new_n505), .A3(G87), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n505), .A2(G49), .A3(G543), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT73), .Z(G288));
  INV_X1    g134(.A(G86), .ZN(new_n560));
  INV_X1    g135(.A(G48), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n519), .A2(new_n560), .B1(new_n511), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(G61), .B1(new_n494), .B2(new_n495), .ZN(new_n564));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT74), .B1(new_n566), .B2(G651), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  AOI211_X1 g143(.A(new_n568), .B(new_n524), .C1(new_n564), .C2(new_n565), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NOR3_X1   g145(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n565), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n518), .B2(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n568), .B1(new_n573), .B2(new_n524), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n566), .A2(KEYINPUT74), .A3(G651), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT75), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n563), .B1(new_n571), .B2(new_n576), .ZN(G305));
  INV_X1    g152(.A(new_n511), .ZN(new_n578));
  AOI22_X1  g153(.A1(G47), .A2(new_n578), .B1(new_n503), .B2(G85), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n524), .B2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n518), .A2(new_n505), .A3(G92), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT10), .ZN(new_n584));
  NAND2_X1  g159(.A1(G79), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G66), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n496), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(G54), .A2(new_n578), .B1(new_n587), .B2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n582), .B1(new_n590), .B2(G868), .ZN(G321));
  XNOR2_X1  g166(.A(G321), .B(KEYINPUT76), .ZN(G284));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NOR2_X1   g168(.A1(G286), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(G299), .B(KEYINPUT77), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(G297));
  XNOR2_X1  g171(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n590), .B1(new_n598), .B2(G860), .ZN(G148));
  NAND2_X1  g174(.A1(new_n590), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G868), .B2(new_n532), .ZN(G323));
  XNOR2_X1  g177(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g178(.A1(new_n463), .A2(G2104), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT12), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT13), .ZN(new_n606));
  INV_X1    g181(.A(G2100), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n463), .A2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n472), .A2(G123), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n471), .A2(G111), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT79), .B(G2096), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n608), .A2(new_n609), .A3(new_n616), .ZN(G156));
  XOR2_X1   g192(.A(KEYINPUT15), .B(G2435), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2438), .ZN(new_n619));
  XOR2_X1   g194(.A(G2427), .B(G2430), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT82), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n619), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(KEYINPUT14), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(G2443), .B(G2446), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n624), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT81), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(G14), .A3(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(G401));
  INV_X1    g212(.A(KEYINPUT18), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n641), .B2(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2096), .B(G2100), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(G227));
  XNOR2_X1  g226(.A(G1971), .B(G1976), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT84), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(new_n655), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT85), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(new_n653), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n652), .B(KEYINPUT19), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n654), .A2(new_n655), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n658), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G229));
  XNOR2_X1  g249(.A(KEYINPUT87), .B(G1971), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(G88), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n506), .B1(new_n519), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n518), .A2(G62), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n524), .B1(new_n679), .B2(new_n499), .ZN(new_n680));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(G16), .A2(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n676), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n683), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n685), .B(new_n675), .C1(G303), .C2(new_n681), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n558), .A2(KEYINPUT86), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(G16), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(G16), .A2(G23), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT33), .B(G1976), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(new_n693), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n687), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  NAND2_X1  g274(.A1(G305), .A2(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n681), .A2(G6), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n570), .B1(new_n567), .B2(new_n569), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n574), .A2(KEYINPUT75), .A3(new_n575), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n562), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n701), .B(new_n699), .C1(new_n705), .C2(new_n681), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n698), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT34), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n710), .B(new_n698), .C1(new_n702), .C2(new_n707), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n681), .A2(G24), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G290), .B2(G16), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G1986), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(G1986), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n463), .A2(G131), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n472), .A2(G119), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n471), .A2(G107), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(G25), .B(new_n721), .S(G29), .Z(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n715), .A2(new_n716), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n711), .A2(new_n712), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n712), .B1(new_n711), .B2(new_n726), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n709), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(KEYINPUT89), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(new_n709), .C1(new_n727), .C2(new_n728), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT36), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n463), .A2(G141), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n472), .A2(G129), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n464), .A2(G105), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT26), .Z(new_n739));
  NAND4_X1  g314(.A1(new_n735), .A2(new_n736), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G32), .B(new_n740), .S(G29), .Z(new_n741));
  XOR2_X1   g316(.A(KEYINPUT27), .B(G1996), .Z(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT99), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n681), .A2(G19), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n532), .B2(new_n681), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G1341), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n463), .A2(G140), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n472), .A2(G128), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n471), .A2(G116), .ZN(new_n750));
  OAI21_X1  g325(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT24), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n755), .B1(new_n761), .B2(G34), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n761), .B2(G34), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G160), .B2(G29), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(G2084), .ZN(new_n765));
  INV_X1    g340(.A(G28), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(KEYINPUT30), .ZN(new_n767));
  AOI21_X1  g342(.A(G29), .B1(new_n766), .B2(KEYINPUT30), .ZN(new_n768));
  OR2_X1    g343(.A1(KEYINPUT31), .A2(G11), .ZN(new_n769));
  NAND2_X1  g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n767), .A2(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n614), .B2(new_n755), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n741), .A2(new_n742), .B1(new_n764), .B2(G2084), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n747), .A2(new_n760), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G171), .A2(new_n681), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G5), .B2(new_n681), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n681), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n681), .ZN(new_n780));
  OAI22_X1  g355(.A1(new_n777), .A2(new_n778), .B1(G1966), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(new_n778), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  INV_X1    g358(.A(new_n780), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n744), .A2(new_n775), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G27), .A2(G29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G164), .B2(G29), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(G2078), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n681), .A2(G20), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT23), .Z(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1956), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n755), .A2(G35), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT100), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G162), .B2(new_n755), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT29), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT29), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(new_n796), .C1(G162), .C2(new_n755), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n789), .B(new_n794), .C1(G2090), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(G2090), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n788), .A2(G2078), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n786), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n755), .A2(G33), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT95), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT25), .ZN(new_n810));
  NAND2_X1  g385(.A1(G115), .A2(G2104), .ZN(new_n811));
  INV_X1    g386(.A(G127), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n462), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n813), .A2(G2105), .B1(new_n463), .B2(G139), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT96), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n807), .B1(new_n816), .B2(G29), .ZN(new_n817));
  INV_X1    g392(.A(G2072), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  NOR2_X1   g395(.A1(G4), .A2(G16), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT91), .Z(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n589), .B2(new_n681), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT93), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT92), .B(G1348), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n817), .A2(new_n818), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT98), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n806), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n734), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(new_n709), .C1(new_n727), .C2(new_n728), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT90), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n832), .B1(new_n729), .B2(KEYINPUT89), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n733), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n831), .A2(new_n836), .ZN(G311));
  OAI21_X1  g412(.A(KEYINPUT101), .B1(new_n831), .B2(new_n836), .ZN(new_n838));
  INV_X1    g413(.A(new_n834), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n711), .A2(new_n726), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT88), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n711), .A2(new_n712), .A3(new_n726), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n841), .A2(new_n842), .B1(KEYINPUT34), .B2(new_n708), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT36), .B1(new_n843), .B2(new_n732), .ZN(new_n844));
  INV_X1    g419(.A(new_n733), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n839), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n734), .A4(new_n830), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n838), .A2(new_n848), .ZN(G150));
  NAND2_X1  g424(.A1(new_n590), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n524), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT102), .ZN(new_n854));
  AOI22_X1  g429(.A1(G55), .A2(new_n578), .B1(new_n503), .B2(G93), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n531), .B2(new_n529), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n532), .A3(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n851), .B(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT103), .B(G860), .Z(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n854), .B2(new_n855), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(G145));
  INV_X1    g443(.A(KEYINPUT108), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n721), .B(KEYINPUT107), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n605), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n463), .A2(G142), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT105), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n472), .A2(G130), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n471), .A2(KEYINPUT106), .A3(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT106), .B1(new_n471), .B2(G118), .ZN(new_n876));
  OR2_X1    g451(.A1(G106), .A2(G2105), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(G2104), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n874), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n871), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n492), .A2(KEYINPUT104), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n483), .A2(new_n491), .A3(new_n884), .A4(new_n485), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n752), .B(new_n740), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n888), .A2(new_n816), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n815), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n882), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n871), .B(new_n880), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n890), .A2(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(G160), .B(new_n614), .Z(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(G162), .Z(new_n898));
  OAI21_X1  g473(.A(new_n869), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n892), .A2(KEYINPUT108), .A3(new_n895), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n896), .B2(new_n898), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT40), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(G395));
  XNOR2_X1  g481(.A(new_n859), .B(new_n600), .ZN(new_n907));
  XNOR2_X1  g482(.A(G299), .B(new_n589), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OR3_X1    g484(.A1(new_n908), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT109), .B1(new_n908), .B2(KEYINPUT41), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(KEYINPUT41), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n688), .A2(new_n690), .ZN(new_n916));
  XNOR2_X1  g491(.A(G305), .B(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G290), .B(G166), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n917), .B(new_n918), .Z(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n915), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n915), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(G868), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n856), .A2(new_n593), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(G295));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n924), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  OR3_X1    g502(.A1(new_n553), .A2(KEYINPUT110), .A3(G301), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n553), .A2(G301), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT110), .B1(G301), .B2(G168), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n860), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n859), .B(new_n928), .C1(new_n929), .C2(new_n930), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n913), .ZN(new_n935));
  INV_X1    g510(.A(new_n919), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n935), .B(new_n936), .C1(new_n908), .C2(new_n934), .ZN(new_n937));
  INV_X1    g512(.A(G37), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n934), .ZN(new_n940));
  INV_X1    g515(.A(new_n908), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n936), .B1(new_n942), .B2(new_n935), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n927), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n934), .A2(new_n908), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n908), .A2(KEYINPUT41), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n932), .A2(new_n933), .B1(new_n946), .B2(new_n912), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n919), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n948), .A2(new_n937), .A3(KEYINPUT43), .A4(new_n938), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT44), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT43), .B1(new_n939), .B2(new_n943), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n948), .A2(new_n937), .A3(new_n927), .A4(new_n938), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n883), .A2(new_n958), .A3(new_n885), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n465), .A2(G40), .A3(new_n469), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(G290), .A2(G1986), .ZN(new_n965));
  AND2_X1   g540(.A1(G290), .A2(G1986), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1996), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT111), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n964), .A2(KEYINPUT111), .A3(new_n968), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n740), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n752), .B(G2067), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n964), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n964), .A2(new_n740), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n975), .B2(new_n968), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT112), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n978));
  INV_X1    g553(.A(new_n976), .ZN(new_n979));
  INV_X1    g554(.A(new_n971), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(new_n969), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n978), .B(new_n979), .C1(new_n981), .C2(new_n740), .ZN(new_n982));
  INV_X1    g557(.A(new_n723), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n721), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n721), .A2(new_n983), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n964), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AND4_X1   g561(.A1(new_n967), .A2(new_n977), .A3(new_n982), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n916), .A2(G1976), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n492), .A2(new_n962), .A3(new_n958), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT116), .B(G8), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1976), .ZN(new_n993));
  AND2_X1   g568(.A1(G288), .A2(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n992), .A2(new_n994), .A3(KEYINPUT52), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(KEYINPUT52), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT117), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n992), .A2(new_n998), .A3(KEYINPUT52), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n995), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1981), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n705), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n574), .A2(new_n575), .ZN(new_n1003));
  OAI21_X1  g578(.A(G1981), .B1(new_n1003), .B2(new_n562), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT118), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT49), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(KEYINPUT118), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n989), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(new_n990), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1000), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n492), .A2(new_n958), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n963), .B1(new_n1015), .B2(new_n960), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n492), .A2(KEYINPUT45), .A3(new_n958), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n492), .A2(new_n1020), .A3(new_n958), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n962), .A3(new_n1021), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n1018), .A2(G1966), .B1(G2084), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(new_n553), .A3(new_n991), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT63), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n883), .A2(KEYINPUT45), .A3(new_n958), .A4(new_n885), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1016), .A2(new_n1027), .ZN(new_n1028));
  OAI22_X1  g603(.A1(new_n1028), .A2(G1971), .B1(G2090), .B2(new_n1022), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  NAND4_X1  g605(.A1(G303), .A2(new_n1030), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT55), .B(G8), .C1(new_n678), .C2(new_n680), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT113), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1031), .A2(new_n1033), .A3(KEYINPUT114), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1036), .A2(KEYINPUT115), .A3(new_n1037), .A4(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1029), .A2(G8), .A3(new_n1041), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1041), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1022), .A2(G2090), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1971), .B1(new_n1016), .B2(new_n1027), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1014), .A2(new_n1026), .A3(new_n1045), .A4(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1045), .A2(new_n1012), .A3(new_n1000), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1046), .B1(new_n1049), .B2(new_n990), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1053), .A2(new_n1055), .A3(new_n1024), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1052), .B1(new_n1056), .B2(KEYINPUT63), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G168), .A2(new_n990), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1023), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1022), .A2(G2084), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1966), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1058), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1060), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1060), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1023), .B2(new_n991), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1059), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT62), .ZN(new_n1069));
  INV_X1    g644(.A(G2078), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1016), .A2(new_n1027), .A3(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1072));
  AOI22_X1  g647(.A1(new_n1071), .A2(new_n1072), .B1(new_n778), .B2(new_n1022), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(KEYINPUT53), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1016), .A2(new_n1075), .A3(new_n1017), .ZN(new_n1076));
  AOI21_X1  g651(.A(G301), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  AND4_X1   g652(.A1(new_n1054), .A2(new_n1045), .A3(new_n1012), .A4(new_n1000), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n1059), .C1(new_n1065), .C2(new_n1067), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1069), .A2(new_n1077), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1002), .B(KEYINPUT119), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G288), .A2(G1976), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1012), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1011), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n1084), .A2(new_n1085), .B1(new_n1013), .B2(new_n1045), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI221_X1 g663(.A(KEYINPUT120), .B1(new_n1013), .B2(new_n1045), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1057), .A2(new_n1081), .A3(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n961), .A2(new_n962), .A3(new_n1027), .A4(new_n1075), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1073), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1092), .B1(new_n1095), .B2(new_n1077), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(G171), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1073), .A2(G301), .A3(new_n1076), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(KEYINPUT54), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1078), .A2(new_n1096), .A3(new_n1099), .A4(new_n1068), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1022), .A2(new_n1101), .B1(new_n759), .B2(new_n1010), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT60), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT122), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1105), .A3(KEYINPUT60), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n590), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(KEYINPUT122), .A3(new_n589), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1102), .A2(KEYINPUT60), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1016), .A2(new_n1027), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT58), .B(G1341), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1111), .A2(G1996), .B1(new_n1010), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n532), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1116), .A3(new_n532), .ZN(new_n1117));
  XOR2_X1   g692(.A(G299), .B(KEYINPUT57), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1022), .A2(new_n793), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1016), .A2(new_n1027), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1119), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1115), .A2(new_n1117), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1122), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1110), .B(new_n1126), .C1(KEYINPUT61), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1102), .A2(new_n589), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1122), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1100), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n987), .B1(new_n1091), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n964), .A2(new_n965), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT48), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n977), .A2(new_n982), .A3(new_n986), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT46), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n980), .A2(new_n969), .B1(KEYINPUT125), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n970), .A2(new_n971), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n974), .A2(new_n975), .A3(new_n1145), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n964), .B(KEYINPUT126), .C1(new_n740), .C2(new_n973), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1146), .A2(new_n1147), .B1(KEYINPUT125), .B2(new_n1140), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT47), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1144), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1139), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n977), .A2(new_n982), .A3(new_n985), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n752), .A2(G2067), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1152), .B1(new_n964), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1136), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g732(.A1(new_n649), .A2(G319), .A3(new_n650), .ZN(new_n1159));
  XNOR2_X1  g733(.A(new_n1159), .B(KEYINPUT127), .ZN(new_n1160));
  NOR2_X1   g734(.A1(G401), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n673), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g736(.A(new_n1162), .B1(new_n902), .B2(new_n903), .ZN(new_n1163));
  AND2_X1   g737(.A1(new_n1163), .A2(new_n954), .ZN(G308));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n954), .ZN(G225));
endmodule


