//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  XOR2_X1   g000(.A(KEYINPUT72), .B(G217), .Z(new_n187));
  INV_X1    g001(.A(G234), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  OAI211_X1 g006(.A(G119), .B(new_n191), .C1(new_n192), .C2(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT73), .B1(new_n195), .B2(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G110), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT24), .B(G110), .Z(new_n200));
  XNOR2_X1  g014(.A(G119), .B(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G125), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n204), .A2(G146), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(G146), .B1(new_n204), .B2(new_n207), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n199), .B(new_n202), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  OAI22_X1  g024(.A1(new_n198), .A2(G110), .B1(new_n201), .B2(new_n200), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n204), .A2(G146), .A3(new_n207), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n203), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT74), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT74), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n210), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G137), .ZN(new_n220));
  INV_X1    g034(.A(G221), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n221), .A2(new_n188), .A3(G953), .ZN(new_n222));
  XOR2_X1   g036(.A(new_n220), .B(new_n222), .Z(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n217), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n216), .A2(KEYINPUT74), .A3(new_n223), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT25), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n230));
  AOI211_X1 g044(.A(new_n230), .B(G902), .C1(new_n225), .C2(new_n226), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n190), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n190), .A2(G902), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(G472), .A2(G902), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT2), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT2), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G113), .ZN(new_n241));
  INV_X1    g055(.A(G116), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(G119), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n195), .A2(G116), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n239), .B(new_n241), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n241), .ZN(new_n246));
  XNOR2_X1  g060(.A(G116), .B(G119), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n245), .A2(new_n248), .A3(KEYINPUT66), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT66), .B1(new_n245), .B2(new_n248), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT30), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n253));
  INV_X1    g067(.A(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT11), .A2(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT65), .A2(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT11), .A2(G134), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT11), .A2(G134), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G137), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n255), .A2(new_n264), .A3(new_n257), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n262), .B1(G134), .B2(G137), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n263), .A2(KEYINPUT67), .A3(new_n267), .ZN(new_n271));
  INV_X1    g085(.A(G143), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT1), .B1(new_n272), .B2(G146), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(G146), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n213), .A2(G143), .ZN(new_n275));
  OAI211_X1 g089(.A(G128), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n213), .A2(G143), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(G146), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n277), .B(new_n278), .C1(KEYINPUT1), .C2(new_n191), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n270), .A2(new_n271), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT0), .A2(G128), .ZN(new_n282));
  NOR2_X1   g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(KEYINPUT64), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n277), .A2(new_n278), .B1(new_n283), .B2(KEYINPUT64), .ZN(new_n286));
  INV_X1    g100(.A(new_n282), .ZN(new_n287));
  XNOR2_X1  g101(.A(G143), .B(G146), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n285), .A2(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n263), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n262), .B1(new_n258), .B2(new_n261), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n252), .B1(new_n281), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n288), .A2(new_n287), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n283), .A2(KEYINPUT64), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n274), .B2(new_n275), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n296), .B2(new_n284), .ZN(new_n297));
  INV_X1    g111(.A(new_n291), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(new_n263), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n276), .A2(new_n279), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n268), .A2(new_n300), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n299), .A2(new_n301), .A3(KEYINPUT30), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n251), .B1(new_n293), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT31), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n300), .B1(new_n268), .B2(new_n269), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n263), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n305), .A2(new_n271), .B1(new_n306), .B2(new_n289), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n245), .A2(new_n248), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n245), .A2(new_n248), .A3(KEYINPUT66), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G237), .A2(G953), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G210), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT27), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G101), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n303), .A2(new_n304), .A3(new_n313), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n281), .A2(new_n312), .A3(new_n292), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n292), .B(new_n252), .C1(new_n268), .C2(new_n300), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n307), .B2(new_n252), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n321), .B1(new_n323), .B2(new_n251), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT68), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n304), .A4(new_n318), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n303), .A2(new_n313), .A3(new_n318), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT31), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n321), .A2(KEYINPUT28), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n251), .B1(new_n299), .B2(new_n301), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT69), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT69), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n251), .B(new_n333), .C1(new_n299), .C2(new_n301), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n313), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n330), .B1(new_n335), .B2(KEYINPUT28), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n329), .B1(new_n318), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n237), .B1(new_n327), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n339));
  INV_X1    g153(.A(new_n237), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(KEYINPUT28), .ZN(new_n341));
  INV_X1    g155(.A(new_n330), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n318), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n343), .A2(new_n344), .B1(KEYINPUT31), .B2(new_n328), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n320), .A2(new_n326), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n339), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n281), .A2(new_n292), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n251), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n313), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT28), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n355), .A2(new_n342), .A3(KEYINPUT29), .A4(new_n318), .ZN(new_n356));
  AOI211_X1 g170(.A(new_n318), .B(new_n321), .C1(new_n323), .C2(new_n251), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n343), .B2(new_n318), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n356), .B(new_n228), .C1(new_n358), .C2(KEYINPUT29), .ZN(new_n359));
  AOI22_X1  g173(.A1(G472), .A2(new_n359), .B1(new_n347), .B2(KEYINPUT32), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n236), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G122), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n364), .A2(KEYINPUT3), .A3(G107), .ZN(new_n365));
  AND2_X1   g179(.A1(KEYINPUT75), .A2(G104), .ZN(new_n366));
  NOR2_X1   g180(.A1(KEYINPUT75), .A2(G104), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n365), .B1(new_n368), .B2(G107), .ZN(new_n369));
  INV_X1    g183(.A(G107), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n366), .B2(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT3), .ZN(new_n372));
  XOR2_X1   g186(.A(KEYINPUT76), .B(G101), .Z(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n371), .B1(G104), .B2(new_n370), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G101), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT78), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n242), .A2(KEYINPUT5), .A3(G119), .ZN(new_n381));
  AOI211_X1 g195(.A(new_n238), .B(new_n381), .C1(KEYINPUT5), .C2(new_n247), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n247), .B2(new_n246), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  OR2_X1    g199(.A1(KEYINPUT75), .A2(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT75), .A2(G104), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n385), .B1(new_n388), .B2(new_n370), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(G107), .A3(new_n387), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(new_n370), .A3(G104), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n374), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n395), .B(G101), .C1(new_n389), .C2(new_n392), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n251), .A3(KEYINPUT80), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n384), .A2(new_n397), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n396), .A2(new_n310), .A3(new_n311), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT80), .B1(new_n399), .B2(new_n394), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n363), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n251), .A3(new_n396), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(new_n362), .A3(new_n384), .A4(new_n397), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n407), .B(new_n363), .C1(new_n398), .C2(new_n400), .ZN(new_n408));
  INV_X1    g222(.A(G125), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n280), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n289), .A2(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G953), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G224), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n412), .B(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n406), .A2(new_n408), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(KEYINPUT7), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT81), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT81), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n420), .B(new_n417), .C1(new_n410), .C2(new_n411), .ZN(new_n421));
  OAI22_X1  g235(.A1(new_n419), .A2(new_n421), .B1(new_n412), .B2(new_n418), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n362), .B(KEYINPUT8), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n383), .B2(new_n377), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n377), .B2(new_n383), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(G902), .B1(new_n426), .B2(new_n405), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G210), .B1(G237), .B2(G902), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT82), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n430), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n416), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(G237), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n413), .A3(G214), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n272), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n314), .A2(G143), .A3(G214), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT18), .A3(G131), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n203), .B(new_n213), .ZN(new_n442));
  NAND2_X1  g256(.A1(KEYINPUT18), .A2(G131), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n262), .B1(new_n438), .B2(new_n439), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n446), .A2(KEYINPUT84), .A3(KEYINPUT17), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT84), .B1(new_n446), .B2(KEYINPUT17), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n439), .ZN(new_n450));
  AOI21_X1  g264(.A(G143), .B1(new_n314), .B2(G214), .ZN(new_n451));
  OAI21_X1  g265(.A(G131), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT17), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n438), .A2(new_n262), .A3(new_n439), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n209), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n212), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n445), .B1(new_n449), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G113), .B(G122), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n364), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(KEYINPUT85), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n208), .A2(new_n209), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n464), .B(new_n455), .C1(new_n447), .C2(new_n448), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n445), .A3(new_n461), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n228), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n463), .A2(KEYINPUT86), .A3(new_n228), .A4(new_n466), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(G475), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n458), .A2(new_n460), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n452), .A2(new_n454), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n203), .B(KEYINPUT19), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n212), .B(new_n473), .C1(new_n475), .C2(G146), .ZN(new_n476));
  INV_X1    g290(.A(new_n460), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n445), .ZN(new_n478));
  NOR2_X1   g292(.A1(G475), .A2(G902), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n472), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n472), .A2(new_n484), .A3(new_n478), .A4(new_n479), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(G234), .A2(G237), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(G952), .A3(new_n413), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT21), .B(G898), .Z(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(G902), .A3(G953), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n491), .B(KEYINPUT88), .Z(new_n492));
  NAND3_X1  g306(.A1(new_n471), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G478), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT9), .B(G234), .Z(new_n497));
  AND3_X1   g311(.A1(new_n187), .A2(new_n497), .A3(new_n413), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n242), .A2(G122), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n242), .A2(G122), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(KEYINPUT14), .ZN(new_n502));
  INV_X1    g316(.A(G122), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(G116), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(G116), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT87), .B1(new_n500), .B2(KEYINPUT14), .ZN(new_n508));
  OAI211_X1 g322(.A(G107), .B(new_n502), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n500), .A3(new_n370), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n272), .A2(G128), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n191), .A2(G143), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n511), .A2(new_n512), .A3(new_n264), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n264), .B1(new_n511), .B2(new_n512), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n509), .B(new_n510), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G107), .B1(new_n501), .B2(new_n504), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n513), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT13), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n272), .A2(KEYINPUT13), .A3(G128), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n519), .A2(new_n520), .A3(new_n512), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n517), .B1(new_n264), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n498), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n515), .A2(new_n522), .A3(new_n498), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n496), .B1(new_n526), .B2(new_n228), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n228), .A3(new_n496), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n493), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n434), .A2(new_n435), .A3(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n374), .A2(new_n280), .A3(new_n376), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n280), .B1(new_n374), .B2(new_n376), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n306), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(KEYINPUT12), .B(new_n306), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT10), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n300), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n378), .A2(new_n380), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n374), .A2(new_n280), .A3(new_n376), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n540), .ZN(new_n544));
  INV_X1    g358(.A(G101), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n369), .B2(new_n372), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n297), .B1(new_n546), .B2(new_n395), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n547), .A2(new_n394), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n547), .B2(new_n394), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n542), .B(new_n544), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n539), .B1(new_n551), .B2(new_n306), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G140), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n413), .A2(G227), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n306), .ZN(new_n557));
  INV_X1    g371(.A(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n551), .B2(new_n306), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n559), .B2(KEYINPUT79), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT79), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n547), .A2(new_n394), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT77), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n547), .A2(new_n394), .A3(new_n548), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n374), .A2(new_n376), .A3(new_n379), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n379), .B1(new_n374), .B2(new_n376), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n568), .A2(new_n541), .B1(new_n540), .B2(new_n543), .ZN(new_n569));
  INV_X1    g383(.A(new_n306), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n565), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n561), .B1(new_n571), .B2(new_n558), .ZN(new_n572));
  OAI211_X1 g386(.A(G469), .B(new_n556), .C1(new_n560), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G469), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n558), .A3(new_n539), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n558), .B1(new_n557), .B2(new_n571), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n574), .B(new_n228), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n574), .A2(new_n228), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n221), .B1(new_n497), .B2(new_n228), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n532), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n361), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n586), .B(new_n373), .Z(G3));
  NOR2_X1   g401(.A1(new_n584), .A2(new_n236), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n228), .B1(new_n327), .B2(new_n337), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G472), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n590), .A2(new_n339), .A3(new_n349), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n429), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n416), .A2(new_n427), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n435), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n428), .B2(new_n429), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n471), .A2(new_n486), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n526), .A2(new_n494), .A3(new_n228), .ZN(new_n598));
  NAND2_X1  g412(.A1(G478), .A2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n526), .A2(KEYINPUT33), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n524), .A2(new_n602), .A3(new_n525), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n600), .B1(new_n604), .B2(G478), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n597), .A2(new_n492), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n592), .A2(new_n594), .A3(new_n596), .A4(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT34), .B(G104), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  AOI21_X1  g424(.A(new_n477), .B1(new_n465), .B2(new_n445), .ZN(new_n611));
  INV_X1    g425(.A(new_n478), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n481), .A3(new_n479), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n483), .A3(KEYINPUT89), .ZN(new_n615));
  OR3_X1    g429(.A1(new_n480), .A2(KEYINPUT89), .A3(new_n482), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n530), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n596), .A2(new_n471), .A3(new_n594), .A4(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n592), .A2(new_n492), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  NOR2_X1   g437(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n216), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n233), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n232), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n585), .A2(new_n591), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT37), .B(G110), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G12));
  NAND2_X1  g444(.A1(new_n351), .A2(new_n360), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n581), .A2(new_n583), .A3(new_n627), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n428), .A2(new_n429), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n435), .A3(new_n594), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n490), .A2(G900), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n488), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n471), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n617), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT90), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n631), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G128), .ZN(G30));
  AND3_X1   g456(.A1(new_n416), .A2(new_n427), .A3(new_n432), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n432), .B1(new_n416), .B2(new_n427), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT92), .Z(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n647), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n434), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n597), .A2(new_n530), .ZN(new_n652));
  NOR4_X1   g466(.A1(new_n651), .A2(new_n595), .A3(new_n627), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT94), .B(KEYINPUT39), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n637), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n581), .A2(new_n583), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT95), .B(KEYINPUT40), .Z(new_n657));
  OR2_X1    g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n347), .A2(KEYINPUT32), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n354), .A2(new_n344), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n328), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT93), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n228), .B1(new_n661), .B2(new_n662), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n351), .A2(new_n659), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n656), .A2(new_n657), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n653), .A2(new_n658), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT96), .B(G143), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G45));
  AND2_X1   g484(.A1(new_n597), .A2(new_n605), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT97), .B1(new_n671), .B2(new_n637), .ZN(new_n672));
  AND4_X1   g486(.A1(KEYINPUT97), .A2(new_n597), .A3(new_n605), .A4(new_n637), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n631), .A2(new_n635), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  OAI21_X1  g490(.A(new_n228), .B1(new_n576), .B2(new_n577), .ZN(new_n677));
  NAND2_X1  g491(.A1(KEYINPUT98), .A2(G469), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n551), .A2(new_n306), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n570), .B1(new_n565), .B2(new_n569), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n555), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(G902), .B1(new_n683), .B2(new_n575), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n678), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n680), .A2(new_n685), .A3(new_n583), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n686), .A2(new_n634), .A3(new_n606), .ZN(new_n687));
  INV_X1    g501(.A(new_n236), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n631), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT99), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n361), .A2(new_n691), .A3(new_n687), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT41), .B(G113), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  INV_X1    g509(.A(new_n492), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n619), .A2(new_n686), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n361), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  NAND2_X1  g513(.A1(new_n531), .A2(new_n627), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n686), .A2(new_n700), .A3(new_n634), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n631), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT100), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n631), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  XOR2_X1   g521(.A(KEYINPUT101), .B(G472), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n589), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n355), .A2(new_n342), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n710), .A2(new_n344), .B1(new_n328), .B2(KEYINPUT31), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n340), .B1(new_n711), .B2(new_n346), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n709), .A2(new_n688), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT102), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n712), .B1(new_n589), .B2(new_n708), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n688), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n652), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n597), .A2(KEYINPUT103), .A3(new_n530), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n596), .A3(new_n594), .A4(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n696), .A3(new_n686), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  AND2_X1   g540(.A1(new_n716), .A2(new_n627), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n686), .A2(new_n634), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n674), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  NAND2_X1  g544(.A1(new_n359), .A2(G472), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n659), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n347), .A2(KEYINPUT32), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n688), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT106), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n736), .B(new_n688), .C1(new_n732), .C2(new_n733), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n643), .A2(new_n644), .A3(new_n595), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n559), .A2(KEYINPUT79), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n571), .A2(new_n561), .A3(new_n558), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n557), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n556), .A2(KEYINPUT104), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n552), .A2(new_n744), .A3(new_n555), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n743), .A3(G469), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n578), .A3(new_n580), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n739), .A2(new_n747), .A3(new_n583), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n748), .A2(KEYINPUT42), .A3(new_n674), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n738), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n631), .A2(new_n748), .A3(new_n688), .A4(new_n674), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(KEYINPUT105), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n361), .A2(new_n753), .A3(new_n674), .A4(new_n748), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n750), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G131), .ZN(G33));
  NAND4_X1  g572(.A1(new_n631), .A2(new_n748), .A3(new_n688), .A4(new_n640), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n605), .A2(new_n486), .A3(new_n471), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT43), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n605), .A2(new_n765), .A3(new_n486), .A4(new_n471), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n764), .B1(new_n763), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n627), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n761), .B1(new_n769), .B2(new_n591), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n769), .A2(new_n761), .A3(new_n591), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n773), .B(new_n761), .C1(new_n769), .C2(new_n591), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n771), .A2(new_n739), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT107), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT45), .A4(new_n745), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n742), .A2(new_n556), .ZN(new_n778));
  OAI211_X1 g592(.A(G469), .B(new_n777), .C1(new_n778), .C2(KEYINPUT45), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n580), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n776), .B1(new_n780), .B2(KEYINPUT46), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n580), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(KEYINPUT107), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(KEYINPUT46), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n781), .A2(new_n578), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n583), .A3(new_n655), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n775), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  XOR2_X1   g603(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(new_n583), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n674), .A2(new_n236), .A3(new_n739), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n631), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n785), .A2(new_n578), .A3(new_n784), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n582), .B1(new_n794), .B2(new_n781), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(KEYINPUT47), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n791), .B(new_n793), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  OR2_X1    g613(.A1(G952), .A2(G953), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n631), .A2(new_n701), .A3(new_n704), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n704), .B1(new_n631), .B2(new_n701), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n725), .B(new_n698), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n691), .A2(new_n631), .A3(new_n688), .A4(new_n687), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n691), .B1(new_n361), .B2(new_n687), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n801), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n719), .A2(new_n724), .B1(new_n361), .B2(new_n697), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n693), .A2(new_n706), .A3(KEYINPUT111), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n645), .A2(new_n595), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n588), .A2(new_n591), .A3(new_n812), .A4(new_n607), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n586), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n815));
  INV_X1    g629(.A(new_n529), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n527), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n528), .A2(KEYINPUT112), .A3(new_n529), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n493), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n434), .A2(new_n820), .A3(new_n435), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n434), .A2(new_n820), .A3(new_n823), .A4(new_n435), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n588), .A2(new_n822), .A3(new_n591), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n628), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT114), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n628), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n814), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n811), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n748), .A2(new_n727), .A3(new_n674), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n818), .A2(new_n817), .A3(new_n615), .A4(new_n616), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n638), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n739), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n632), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n631), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n759), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n723), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n232), .A2(new_n626), .A3(new_n637), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n579), .B1(new_n684), .B2(new_n574), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n582), .B(new_n840), .C1(new_n841), .C2(new_n746), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n339), .A2(new_n349), .A3(new_n350), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n659), .A2(new_n665), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n839), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n641), .A2(new_n675), .A3(new_n845), .A4(new_n729), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n838), .B1(new_n846), .B2(KEYINPUT52), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n641), .A2(new_n729), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n675), .A4(new_n845), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n757), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n641), .A2(new_n729), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT53), .B1(new_n852), .B2(KEYINPUT52), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n831), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n814), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n825), .A2(new_n828), .A3(new_n628), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n828), .B1(new_n825), .B2(new_n628), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n808), .B2(new_n810), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n757), .A2(new_n847), .A3(new_n850), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT53), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT54), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT115), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n804), .B2(new_n807), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n693), .A2(new_n706), .A3(KEYINPUT116), .A4(new_n809), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n852), .B2(KEYINPUT52), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n865), .A2(new_n830), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n851), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n861), .A2(new_n870), .A3(KEYINPUT54), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n873), .B(KEYINPUT54), .C1(new_n854), .C2(new_n861), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n863), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n488), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n766), .A2(new_n763), .A3(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n719), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n686), .A2(new_n435), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n651), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n680), .A2(new_n685), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(new_n583), .A3(new_n595), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n648), .A2(new_n650), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT117), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n878), .A2(KEYINPUT50), .A3(new_n881), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT50), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n881), .A2(new_n885), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n719), .A2(new_n877), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n645), .A2(new_n435), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n686), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n893), .A2(new_n877), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n727), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(KEYINPUT118), .A3(new_n727), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n893), .A2(new_n688), .A3(new_n876), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n666), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n597), .A2(new_n605), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n897), .A2(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT119), .B1(new_n891), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n791), .B1(new_n795), .B2(new_n797), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n882), .A2(new_n582), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n878), .A2(new_n739), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n891), .A2(new_n902), .A3(KEYINPUT119), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT51), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n738), .A2(new_n894), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT48), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n900), .A2(new_n671), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(G952), .A3(new_n413), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n728), .B2(new_n878), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n907), .B1(new_n904), .B2(new_n905), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n891), .A2(new_n902), .A3(KEYINPUT51), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n913), .B(new_n916), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT120), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n913), .ZN(new_n921));
  INV_X1    g735(.A(new_n917), .ZN(new_n922));
  INV_X1    g736(.A(new_n918), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  INV_X1    g739(.A(new_n910), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n917), .A2(new_n926), .A3(new_n903), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n924), .B(new_n925), .C1(new_n927), .C2(KEYINPUT51), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n920), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n800), .B1(new_n875), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT49), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n882), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n882), .A2(new_n931), .ZN(new_n933));
  NOR4_X1   g747(.A1(new_n762), .A2(new_n236), .A3(new_n582), .A4(new_n595), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OR3_X1    g749(.A1(new_n935), .A2(new_n666), .A3(new_n884), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n930), .A2(new_n936), .ZN(G75));
  OAI211_X1 g751(.A(G210), .B(G902), .C1(new_n861), .C2(new_n870), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n406), .A2(new_n408), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n415), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n944), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n938), .A2(new_n939), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n413), .A2(G952), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n945), .A2(KEYINPUT122), .A3(new_n947), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(G51));
  XNOR2_X1  g768(.A(new_n579), .B(KEYINPUT57), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n861), .A2(new_n870), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT54), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n955), .B1(new_n958), .B2(new_n871), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n577), .B2(new_n576), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n861), .A2(new_n870), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(G902), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(new_n779), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n948), .B1(new_n960), .B2(new_n963), .ZN(G54));
  INV_X1    g778(.A(new_n613), .ZN(new_n965));
  NAND2_X1  g779(.A1(KEYINPUT58), .A2(G475), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n949), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(G60));
  INV_X1    g784(.A(new_n604), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n599), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n971), .B(new_n973), .C1(new_n958), .C2(new_n871), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n949), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n875), .A2(new_n973), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n604), .ZN(G63));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT60), .Z(new_n979));
  OAI211_X1 g793(.A(new_n625), .B(new_n979), .C1(new_n861), .C2(new_n870), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT61), .B1(new_n980), .B2(KEYINPUT124), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n227), .B1(new_n961), .B2(new_n979), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n949), .ZN(new_n983));
  OR3_X1    g797(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G66));
  NAND2_X1  g800(.A1(new_n489), .A2(G224), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(G953), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n859), .B2(G953), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n941), .B1(G898), .B2(new_n413), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  AOI21_X1  g805(.A(new_n413), .B1(G227), .B2(G900), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n323), .B(new_n475), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n994));
  INV_X1    g808(.A(new_n798), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n848), .A2(new_n675), .A3(new_n759), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n723), .B1(new_n735), .B2(new_n737), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n786), .A2(new_n997), .A3(new_n583), .A4(new_n655), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n996), .B(new_n998), .C1(new_n775), .C2(new_n787), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(G953), .B1(new_n1000), .B2(new_n757), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n413), .A2(G900), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT125), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n994), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n999), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n757), .A3(new_n798), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n413), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1008), .A2(KEYINPUT126), .A3(new_n1003), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n993), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n993), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n668), .A2(new_n675), .A3(new_n848), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT62), .Z(new_n1013));
  NAND2_X1  g827(.A1(new_n597), .A2(new_n605), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n819), .A2(new_n597), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n892), .B(new_n656), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n361), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1013), .A2(new_n788), .A3(new_n798), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1011), .B1(new_n1018), .B2(new_n413), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n992), .B1(new_n1010), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(KEYINPUT126), .B1(new_n1008), .B2(new_n1003), .ZN(new_n1021));
  AOI211_X1 g835(.A(new_n994), .B(new_n1004), .C1(new_n1007), .C2(new_n413), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1011), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n992), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1019), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1020), .A2(new_n1026), .ZN(G72));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  OAI21_X1  g843(.A(new_n1029), .B1(new_n1018), .B2(new_n831), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n324), .A2(new_n344), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1029), .B1(new_n1007), .B2(new_n831), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n357), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1032), .A2(new_n1034), .A3(new_n949), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n854), .A2(new_n861), .ZN(new_n1036));
  INV_X1    g850(.A(new_n357), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(new_n1029), .ZN(new_n1038));
  OR2_X1    g852(.A1(new_n1038), .A2(new_n1031), .ZN(new_n1039));
  OAI21_X1  g853(.A(KEYINPUT127), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  OR3_X1    g854(.A1(new_n1036), .A2(KEYINPUT127), .A3(new_n1039), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1035), .B1(new_n1040), .B2(new_n1041), .ZN(G57));
endmodule


