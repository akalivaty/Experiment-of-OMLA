//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT84), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n204));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n206));
  OR2_X1    g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n205), .B1(new_n209), .B2(KEYINPUT72), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT72), .ZN(new_n211));
  XOR2_X1   g010(.A(G197gat), .B(G204gat), .Z(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(new_n206), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(KEYINPUT72), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n210), .B1(new_n215), .B2(new_n205), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n204), .B1(new_n216), .B2(KEYINPUT29), .ZN(new_n217));
  AND2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G141gat), .B(G148gat), .Z(new_n221));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT76), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT76), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n218), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n221), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n229), .A2(KEYINPUT77), .A3(new_n218), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n220), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n233));
  NAND2_X1  g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT80), .B1(new_n218), .B2(new_n219), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(KEYINPUT2), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G141gat), .ZN(new_n239));
  OR3_X1    g038(.A1(new_n239), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT79), .B1(new_n239), .B2(G148gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT78), .B(G141gat), .ZN(new_n242));
  INV_X1    g041(.A(G148gat), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n240), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n231), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n217), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT77), .B1(new_n229), .B2(new_n218), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n223), .A2(new_n225), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(new_n227), .A3(new_n234), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n250), .A3(new_n221), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n251), .A2(new_n220), .B1(new_n238), .B2(new_n244), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT29), .B1(new_n252), .B2(new_n204), .ZN(new_n253));
  INV_X1    g052(.A(new_n216), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n203), .B1(new_n247), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT86), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n202), .B1(new_n217), .B2(new_n246), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n216), .B1(new_n253), .B2(KEYINPUT85), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT85), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n257), .B(new_n258), .C1(new_n259), .C2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n262), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n253), .A2(KEYINPUT85), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n216), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n257), .B1(new_n268), .B2(new_n258), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n256), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT31), .B(G50gat), .Z(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G78gat), .B(G106gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(G22gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n271), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n256), .B(new_n275), .C1(new_n265), .C2(new_n269), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(new_n274), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G113gat), .ZN(new_n281));
  INV_X1    g080(.A(G120gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284));
  NAND2_X1  g083(.A1(G113gat), .A2(G120gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(G127gat), .A2(G134gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(G127gat), .A2(G134gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT68), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G127gat), .B(G134gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT1), .B1(new_n281), .B2(new_n282), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n285), .A4(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT67), .B(G134gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G127gat), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n288), .B1(new_n293), .B2(new_n285), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n290), .A2(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT23), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n306), .A2(KEYINPUT25), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n305), .A2(new_n314), .A3(KEYINPUT23), .ZN(new_n315));
  INV_X1    g114(.A(new_n309), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n305), .B2(KEYINPUT23), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(new_n306), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n301), .A2(KEYINPUT64), .A3(new_n302), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n313), .A2(new_n315), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n311), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n309), .B1(new_n305), .B2(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n300), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT27), .B(G183gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT66), .ZN(new_n329));
  INV_X1    g128(.A(G183gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT27), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n332));
  INV_X1    g131(.A(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n327), .B1(new_n329), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n333), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n326), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n298), .B1(new_n322), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n298), .ZN(new_n339));
  INV_X1    g138(.A(new_n326), .ZN(new_n340));
  XOR2_X1   g139(.A(KEYINPUT27), .B(G183gat), .Z(new_n341));
  INV_X1    g140(.A(KEYINPUT66), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(G190gat), .B1(new_n331), .B2(KEYINPUT66), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT28), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n336), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n301), .A2(KEYINPUT64), .A3(new_n302), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT64), .B1(new_n301), .B2(new_n302), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G169gat), .ZN(new_n351));
  INV_X1    g150(.A(G176gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT23), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n306), .B1(new_n353), .B2(KEYINPUT65), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n354), .A2(new_n315), .A3(new_n309), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT25), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n339), .B(new_n347), .C1(new_n356), .C2(new_n311), .ZN(new_n357));
  INV_X1    g156(.A(G227gat), .ZN(new_n358));
  INV_X1    g157(.A(G233gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n338), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT32), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT69), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n364), .A3(KEYINPUT32), .ZN(new_n365));
  XNOR2_X1  g164(.A(G15gat), .B(G43gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G71gat), .B(G99gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n361), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n363), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n360), .B1(new_n338), .B2(new_n357), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT70), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n361), .B(KEYINPUT32), .C1(new_n369), .C2(new_n368), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n371), .B2(new_n375), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT34), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n372), .B2(new_n373), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n379), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n371), .A2(new_n375), .ZN(new_n382));
  INV_X1    g181(.A(new_n374), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n277), .B(new_n280), .C1(new_n380), .C2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  OAI21_X1  g189(.A(new_n260), .B1(new_n322), .B2(new_n337), .ZN(new_n391));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n392), .B(KEYINPUT73), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n347), .B1(new_n356), .B2(new_n311), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n393), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n254), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n320), .A2(new_n321), .ZN(new_n400));
  INV_X1    g199(.A(new_n311), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n337), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n399), .B1(new_n402), .B2(new_n394), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(KEYINPUT74), .A3(new_n393), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n403), .A2(new_n404), .B1(new_n394), .B2(new_n391), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n390), .B(new_n398), .C1(new_n405), .C2(new_n254), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT30), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n403), .A2(new_n404), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n254), .B1(new_n409), .B2(new_n395), .ZN(new_n410));
  INV_X1    g209(.A(new_n398), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT75), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n390), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT75), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n414), .B(new_n398), .C1(new_n405), .C2(new_n254), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n406), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n408), .B1(new_n417), .B2(KEYINPUT30), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT35), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n420), .A2(KEYINPUT81), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n231), .A2(new_n298), .A3(new_n245), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n298), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n339), .B1(new_n252), .B2(new_n204), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n231), .A2(new_n204), .A3(new_n245), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n424), .B(new_n425), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n421), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n246), .A2(new_n339), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n422), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n420), .B1(new_n433), .B2(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G1gat), .B(G29gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT0), .ZN(new_n437));
  XNOR2_X1  g236(.A(G57gat), .B(G85gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(new_n430), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT5), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n252), .A2(new_n204), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n339), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n445), .A2(new_n429), .A3(new_n424), .A4(new_n425), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(new_n446), .A3(new_n421), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n435), .A2(new_n440), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449));
  OR3_X1    g248(.A1(new_n448), .A2(KEYINPUT83), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT83), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n431), .A2(new_n434), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n442), .B1(new_n446), .B2(new_n421), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n439), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n449), .A3(new_n448), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n418), .A2(new_n419), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n387), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n448), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n435), .A2(new_n447), .A3(KEYINPUT82), .A4(new_n440), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(new_n449), .A3(new_n454), .A4(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n450), .A3(new_n451), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n418), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT35), .B1(new_n387), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(KEYINPUT89), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n274), .B1(new_n272), .B2(new_n276), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n379), .B1(new_n376), .B2(new_n377), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n384), .A2(new_n385), .A3(new_n381), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n469), .A2(new_n472), .A3(new_n463), .A4(new_n418), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT35), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n280), .A2(new_n277), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n464), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT71), .A4(KEYINPUT36), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT36), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT71), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT39), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n428), .A2(new_n483), .A3(new_n430), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n428), .A2(new_n430), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT39), .B1(new_n433), .B2(new_n430), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n439), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT87), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n448), .B1(new_n488), .B2(KEYINPUT40), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(KEYINPUT40), .B2(new_n488), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n417), .A2(KEYINPUT30), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(new_n408), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n398), .B1(new_n405), .B2(new_n254), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n494), .A2(KEYINPUT37), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n412), .A2(KEYINPUT37), .A3(new_n415), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n413), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(KEYINPUT88), .A3(new_n413), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n493), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n405), .A2(new_n216), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n395), .A2(new_n397), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(new_n216), .ZN(new_n506));
  AOI211_X1 g305(.A(KEYINPUT38), .B(new_n390), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n407), .B1(new_n507), .B2(new_n495), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n508), .A2(new_n450), .A3(new_n451), .A4(new_n455), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n492), .B(new_n469), .C1(new_n502), .C2(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n466), .A2(new_n475), .B1(new_n482), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n513), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  NOR3_X1   g313(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT90), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  OAI221_X1 g317(.A(new_n514), .B1(KEYINPUT15), .B2(new_n513), .C1(new_n516), .C2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  OAI22_X1  g320(.A1(new_n518), .A2(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(KEYINPUT15), .A3(new_n513), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G1gat), .B2(new_n526), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n524), .B(KEYINPUT17), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(new_n531), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(KEYINPUT18), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(KEYINPUT18), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n524), .B(new_n531), .Z(new_n539));
  XOR2_X1   g338(.A(new_n535), .B(KEYINPUT13), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G197gat), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT11), .B(G169gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n546), .B(KEYINPUT12), .Z(new_n547));
  OR2_X1    g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G57gat), .B(G64gat), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n552));
  OR2_X1    g351(.A1(G71gat), .A2(G78gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT9), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n554), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G57gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n558), .B(new_n560), .C1(new_n551), .C2(KEYINPUT91), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n565));
  AND2_X1   g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G127gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n531), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n564), .B2(KEYINPUT21), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n568), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G155gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n575), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT93), .ZN(new_n580));
  XOR2_X1   g379(.A(G134gat), .B(G162gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT7), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(KEYINPUT8), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n585), .B1(new_n525), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT95), .Z(new_n597));
  XOR2_X1   g396(.A(new_n594), .B(KEYINPUT94), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n533), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n584), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n597), .A2(new_n584), .A3(new_n599), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n582), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT96), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n600), .A2(KEYINPUT97), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(KEYINPUT97), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n605), .A2(new_n606), .A3(new_n582), .A4(new_n602), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n578), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n564), .A2(new_n595), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n562), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT10), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT98), .Z(new_n613));
  NAND3_X1  g412(.A1(new_n564), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT99), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT100), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n610), .A2(new_n611), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n621), .A2(new_n616), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n615), .A2(new_n623), .A3(new_n618), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n620), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n616), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(new_n622), .A3(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n512), .A2(new_n550), .A3(new_n609), .A4(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(new_n463), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT101), .B(G1gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1324gat));
  INV_X1    g437(.A(new_n635), .ZN(new_n639));
  INV_X1    g438(.A(new_n418), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n530), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT16), .B(G8gat), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n635), .A2(new_n418), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT42), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n644), .B1(KEYINPUT42), .B2(new_n643), .ZN(G1325gat));
  AND2_X1   g444(.A1(new_n481), .A2(new_n478), .ZN(new_n646));
  OAI21_X1  g445(.A(G15gat), .B1(new_n635), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n472), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n648), .A2(G15gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n635), .B2(new_n649), .ZN(G1326gat));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n469), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT43), .B(G22gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1327gat));
  INV_X1    g452(.A(new_n608), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n465), .A2(KEYINPUT89), .ZN(new_n655));
  INV_X1    g454(.A(new_n458), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n475), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n482), .A2(new_n510), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n578), .ZN(new_n660));
  INV_X1    g459(.A(new_n550), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n660), .A2(new_n661), .A3(new_n633), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n463), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n520), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT45), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT35), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n474), .B1(new_n473), .B2(KEYINPUT35), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n669), .A2(new_n670), .A3(new_n458), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n510), .A2(new_n646), .A3(new_n477), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n608), .B(new_n668), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n659), .A2(KEYINPUT104), .A3(new_n668), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n659), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(KEYINPUT102), .B(KEYINPUT44), .C1(new_n511), .C2(new_n654), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n662), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n683), .A2(new_n463), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n666), .B1(new_n685), .B2(new_n520), .ZN(G1328gat));
  NAND3_X1  g485(.A1(new_n663), .A2(new_n521), .A3(new_n640), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n688));
  NAND2_X1  g487(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  NOR3_X1   g489(.A1(new_n683), .A2(new_n418), .A3(new_n684), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(new_n521), .ZN(G1329gat));
  NOR3_X1   g491(.A1(new_n683), .A2(new_n646), .A3(new_n684), .ZN(new_n693));
  INV_X1    g492(.A(G43gat), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT106), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n663), .A2(new_n694), .A3(new_n472), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n693), .B2(new_n694), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n695), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n699), .A2(new_n700), .ZN(G1330gat));
  INV_X1    g500(.A(G50gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n663), .A2(new_n702), .A3(new_n476), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n683), .A2(new_n469), .A3(new_n684), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G50gat), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  OAI211_X1 g506(.A(KEYINPUT48), .B(new_n703), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n703), .B1(new_n704), .B2(new_n702), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n709), .A2(KEYINPUT107), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT107), .B1(new_n709), .B2(new_n710), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n708), .B1(new_n711), .B2(new_n712), .ZN(G1331gat));
  NAND4_X1  g512(.A1(new_n512), .A2(new_n661), .A3(new_n609), .A4(new_n633), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n463), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n559), .ZN(G1332gat));
  XOR2_X1   g515(.A(new_n714), .B(KEYINPUT109), .Z(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n640), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT49), .B(G64gat), .Z(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n718), .B2(new_n720), .ZN(G1333gat));
  INV_X1    g520(.A(G71gat), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n646), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n714), .B2(new_n648), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n717), .A2(new_n476), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g528(.A1(new_n659), .A2(new_n661), .A3(new_n578), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n732), .A2(KEYINPUT110), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n730), .A2(new_n731), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(new_n589), .A3(new_n664), .A4(new_n633), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n578), .A2(new_n661), .A3(new_n633), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n677), .B2(new_n682), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n463), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n742), .ZN(G1336gat));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n634), .A2(G92gat), .A3(new_n418), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n735), .A2(new_n736), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n741), .A2(new_n418), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748));
  OAI21_X1  g547(.A(G92gat), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n741), .A2(KEYINPUT111), .A3(new_n418), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n744), .B(new_n746), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n747), .A2(new_n590), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n734), .A2(new_n732), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(new_n745), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(G1337gat));
  NOR3_X1   g555(.A1(new_n634), .A2(G99gat), .A3(new_n648), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n737), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G99gat), .B1(new_n741), .B2(new_n646), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1338gat));
  NOR3_X1   g559(.A1(new_n634), .A2(G106gat), .A3(new_n469), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n735), .A2(new_n736), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763));
  INV_X1    g562(.A(G106gat), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n469), .B(new_n739), .C1(new_n677), .C2(new_n682), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n753), .A2(new_n761), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n764), .B1(new_n740), .B2(new_n476), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n765), .A2(KEYINPUT112), .A3(new_n764), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n767), .B(KEYINPUT53), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT112), .B1(new_n765), .B2(new_n764), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n740), .A2(new_n476), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n770), .A3(G106gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n775), .A2(new_n777), .A3(new_n768), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n767), .B1(new_n778), .B2(KEYINPUT53), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n766), .B1(new_n774), .B2(new_n779), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT54), .B1(new_n620), .B2(new_n624), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n615), .B2(new_n616), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n613), .A2(new_n617), .A3(new_n614), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n629), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n781), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n624), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n623), .B1(new_n615), .B2(new_n618), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n783), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n629), .A4(new_n786), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n788), .A2(new_n792), .A3(new_n550), .A4(new_n632), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n534), .A2(new_n535), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n539), .A2(new_n540), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n546), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n633), .A2(new_n548), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n654), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n548), .A2(new_n796), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n604), .B2(new_n607), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n801), .A2(new_n788), .A3(new_n632), .A4(new_n792), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(KEYINPUT114), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n608), .B1(new_n793), .B2(new_n797), .ZN(new_n805));
  INV_X1    g604(.A(new_n802), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n803), .A2(new_n578), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n609), .A2(new_n661), .A3(new_n634), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n664), .A3(new_n469), .A4(new_n472), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n418), .A3(new_n550), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT115), .B1(new_n810), .B2(new_n469), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  AOI211_X1 g615(.A(new_n816), .B(new_n476), .C1(new_n808), .C2(new_n809), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n648), .A2(new_n640), .A3(new_n463), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n661), .A2(new_n281), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n814), .A2(new_n281), .B1(new_n821), .B2(new_n822), .ZN(G1340gat));
  OAI211_X1 g622(.A(new_n633), .B(new_n819), .C1(new_n815), .C2(new_n817), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(KEYINPUT117), .A3(G120gat), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT117), .B1(new_n824), .B2(G120gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n813), .A2(new_n418), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n633), .A2(new_n282), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n825), .A2(new_n826), .B1(new_n827), .B2(new_n828), .ZN(G1341gat));
  OAI21_X1  g628(.A(G127gat), .B1(new_n820), .B2(new_n578), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n578), .A2(G127gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n827), .B2(new_n831), .ZN(G1342gat));
  NOR2_X1   g631(.A1(new_n654), .A2(new_n295), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n418), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT56), .ZN(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n820), .B2(new_n654), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n813), .A2(new_n837), .A3(new_n418), .A4(new_n833), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(G1343gat));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n463), .B1(new_n808), .B2(new_n809), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n646), .A2(new_n476), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n846), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n843), .B1(new_n841), .B2(KEYINPUT119), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(KEYINPUT120), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n661), .A2(G141gat), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n847), .A2(new_n850), .A3(new_n418), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n798), .A2(KEYINPUT118), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n793), .A2(new_n797), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n654), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n660), .B1(new_n856), .B2(new_n802), .ZN(new_n857));
  INV_X1    g656(.A(new_n809), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n476), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT57), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n810), .A2(new_n861), .A3(new_n476), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n646), .A2(new_n664), .A3(new_n418), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n860), .A2(new_n550), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT58), .B1(new_n864), .B2(new_n242), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n852), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n864), .A2(new_n242), .ZN(new_n867));
  AND4_X1   g666(.A1(new_n418), .A2(new_n848), .A3(new_n849), .A4(new_n851), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT58), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n634), .A2(G148gat), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n847), .A2(new_n850), .A3(new_n418), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n634), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(KEYINPUT59), .A3(new_n243), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n809), .A2(KEYINPUT121), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n609), .A2(new_n878), .A3(new_n661), .A4(new_n634), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n855), .A2(new_n654), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n854), .B1(new_n793), .B2(new_n797), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n802), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n883), .B2(new_n578), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT122), .B(new_n861), .C1(new_n884), .C2(new_n469), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n810), .A2(KEYINPUT57), .A3(new_n476), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n476), .B1(new_n857), .B2(new_n880), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT122), .B1(new_n888), .B2(new_n861), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n633), .B(new_n863), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n876), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n872), .B1(new_n875), .B2(new_n891), .ZN(G1345gat));
  NOR2_X1   g691(.A1(new_n578), .A2(G155gat), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n847), .A2(new_n850), .A3(new_n418), .A4(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G155gat), .B1(new_n873), .B2(new_n578), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1346gat));
  NOR2_X1   g695(.A1(new_n654), .A2(G162gat), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n847), .A2(new_n850), .A3(new_n418), .A4(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G162gat), .B1(new_n873), .B2(new_n654), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1347gat));
  AOI21_X1  g699(.A(new_n664), .B1(new_n808), .B2(new_n809), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n387), .A2(new_n418), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n550), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n648), .A2(new_n664), .A3(new_n418), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n818), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n661), .A2(new_n351), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G1348gat));
  OAI211_X1 g707(.A(new_n633), .B(new_n905), .C1(new_n815), .C2(new_n817), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G176gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n903), .A2(new_n352), .A3(new_n633), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT123), .ZN(G1349gat));
  OAI211_X1 g712(.A(new_n660), .B(new_n905), .C1(new_n815), .C2(new_n817), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G183gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n903), .A2(new_n328), .A3(new_n660), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  OAI211_X1 g717(.A(new_n608), .B(new_n905), .C1(new_n815), .C2(new_n817), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G190gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n922), .A3(G190gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(KEYINPUT61), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n903), .A2(new_n333), .A3(new_n608), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT124), .Z(new_n926));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n920), .A2(KEYINPUT125), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(G1351gat));
  AND3_X1   g728(.A1(new_n901), .A2(new_n640), .A3(new_n844), .ZN(new_n930));
  INV_X1    g729(.A(G197gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(new_n550), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n646), .A2(new_n463), .A3(new_n640), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n550), .B(new_n933), .C1(new_n887), .C2(new_n889), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G197gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n934), .A2(new_n935), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(G1352gat));
  OR2_X1    g738(.A1(new_n887), .A2(new_n889), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n633), .A3(new_n933), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G204gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  AOI21_X1  g742(.A(G204gat), .B1(new_n943), .B2(KEYINPUT62), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n930), .A2(new_n633), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n942), .A2(new_n947), .ZN(G1353gat));
  INV_X1    g747(.A(G211gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n949), .A3(new_n660), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n660), .B(new_n933), .C1(new_n887), .C2(new_n889), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n951), .B2(G211gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1354gat));
  INV_X1    g753(.A(G218gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n930), .A2(new_n955), .A3(new_n608), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n608), .A3(new_n933), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n958), .B2(new_n955), .ZN(G1355gat));
endmodule


