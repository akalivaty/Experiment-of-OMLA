//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n467), .A2(new_n468), .A3(G137), .A4(new_n462), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n462), .B1(new_n474), .B2(new_n475), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT69), .Z(new_n486));
  NAND2_X1  g061(.A1(new_n467), .A2(new_n462), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI211_X1 g063(.A(new_n483), .B(new_n486), .C1(G136), .C2(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n463), .B2(new_n464), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT70), .B(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n496), .B(new_n500), .C1(new_n464), .C2(new_n463), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n494), .B1(new_n499), .B2(new_n501), .ZN(G164));
  AND2_X1   g077(.A1(KEYINPUT71), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT71), .A2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NOR3_X1   g080(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n505), .A2(KEYINPUT72), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n512), .A2(G88), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n512), .A2(G50), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n503), .A2(new_n504), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(G62), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(KEYINPUT73), .B1(G75), .B2(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n519), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n518), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n515), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n508), .ZN(new_n537));
  NAND2_X1  g112(.A1(KEYINPUT71), .A2(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(KEYINPUT6), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n539), .A2(G543), .A3(new_n510), .A4(new_n509), .ZN(new_n540));
  INV_X1    g115(.A(G51), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n509), .A2(new_n510), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n542), .A2(new_n515), .A3(new_n539), .ZN(new_n543));
  INV_X1    g118(.A(G89), .ZN(new_n544));
  OAI221_X1 g119(.A(new_n535), .B1(new_n540), .B2(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G168));
  INV_X1    g121(.A(new_n543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G90), .ZN(new_n548));
  INV_X1    g123(.A(new_n540), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G52), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n519), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(new_n547), .A2(G81), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n549), .A2(G43), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n519), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n524), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n543), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n512), .A2(new_n573), .A3(G53), .A4(G543), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n540), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n572), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n545), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n547), .A2(G89), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n549), .A2(G51), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n581), .A2(KEYINPUT74), .A3(new_n582), .A4(new_n535), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G286));
  INV_X1    g160(.A(new_n519), .ZN(new_n586));
  INV_X1    g161(.A(new_n528), .ZN(new_n587));
  NAND2_X1  g162(.A1(G75), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(new_n526), .B2(new_n527), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n586), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n590), .A2(new_n516), .A3(new_n517), .ZN(G303));
  OAI21_X1  g166(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n592));
  INV_X1    g167(.A(G49), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI221_X1 g169(.A(new_n592), .B1(new_n540), .B2(new_n593), .C1(new_n543), .C2(new_n594), .ZN(G288));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n524), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n586), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n542), .A2(G48), .A3(G543), .A4(new_n539), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n542), .A2(G86), .A3(new_n515), .A4(new_n539), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G305));
  NAND2_X1  g180(.A1(new_n547), .A2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n549), .A2(G47), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(new_n519), .C2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT76), .B(KEYINPUT10), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n543), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n543), .B2(new_n611), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n524), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n549), .A2(G54), .B1(G651), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n610), .B1(new_n620), .B2(G868), .ZN(G321));
  XOR2_X1   g196(.A(G321), .B(KEYINPUT77), .Z(G284));
  NOR2_X1   g197(.A1(G299), .A2(G868), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n584), .ZN(G297));
  AOI21_X1  g199(.A(new_n623), .B1(G868), .B2(new_n584), .ZN(G280));
  XNOR2_X1  g200(.A(KEYINPUT78), .B(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n620), .B1(G860), .B2(new_n626), .ZN(G148));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n559), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n620), .A2(new_n626), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n629), .B1(new_n631), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n484), .A2(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n462), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G135), .ZN(new_n637));
  OAI221_X1 g212(.A(new_n634), .B1(new_n635), .B2(new_n636), .C1(new_n637), .C2(new_n487), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND3_X1  g214(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n639), .A2(new_n644), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT80), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT17), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n664), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n670), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n668), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n666), .A3(new_n664), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  NAND3_X1  g251(.A1(new_n665), .A2(new_n670), .A3(new_n667), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n684), .A2(new_n685), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n683), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n683), .A2(new_n691), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n689), .A2(new_n690), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n696), .A2(new_n697), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n681), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n696), .A2(new_n697), .ZN(new_n703));
  INV_X1    g278(.A(new_n681), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n703), .A2(new_n704), .A3(new_n698), .ZN(new_n705));
  AND3_X1   g280(.A1(new_n701), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n702), .B1(new_n701), .B2(new_n705), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(G229));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G35), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G162), .B2(new_n709), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT29), .Z(new_n712));
  INV_X1    g287(.A(G2090), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT91), .B(KEYINPUT23), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT92), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G20), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n716), .B(new_n718), .Z(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G299), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT93), .B(G1956), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n714), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n725));
  NAND3_X1  g300(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G139), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n487), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(new_n462), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(new_n709), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n709), .B2(G33), .ZN(new_n734));
  INV_X1    g309(.A(G2072), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n709), .A2(G26), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n488), .A2(G140), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n484), .A2(G128), .ZN(new_n740));
  OR2_X1    g315(.A1(G104), .A2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n741), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n738), .B1(new_n744), .B2(new_n709), .ZN(new_n745));
  INV_X1    g320(.A(G2067), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT31), .B(G11), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(G28), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n709), .B1(new_n749), .B2(G28), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n748), .B1(new_n750), .B2(new_n751), .C1(new_n638), .C2(new_n709), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n709), .A2(G32), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT26), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n484), .A2(G129), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n758));
  INV_X1    g333(.A(G141), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n487), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n753), .B1(new_n761), .B2(new_n709), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT27), .B(G1996), .Z(new_n763));
  AOI21_X1  g338(.A(new_n752), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n736), .A2(new_n747), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n620), .A2(new_n717), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G4), .B2(new_n717), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT86), .B(G1348), .Z(new_n769));
  AOI21_X1  g344(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n712), .B2(new_n713), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n723), .A2(new_n724), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n734), .A2(new_n735), .ZN(new_n774));
  INV_X1    g349(.A(G2078), .ZN(new_n775));
  NOR2_X1   g350(.A1(G164), .A2(new_n709), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G27), .B2(new_n709), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n559), .A2(G16), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n717), .A2(G19), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n779), .B1(G1341), .B2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT24), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n709), .B1(new_n785), .B2(G34), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(KEYINPUT88), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(KEYINPUT88), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n785), .B2(G34), .ZN(new_n789));
  AOI22_X1  g364(.A1(G160), .A2(G29), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2084), .ZN(new_n791));
  NOR2_X1   g366(.A1(G5), .A2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT90), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G301), .B2(new_n717), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1961), .Z(new_n795));
  NOR2_X1   g370(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G1341), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n717), .A2(G21), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G168), .B2(new_n717), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n782), .A2(new_n797), .B1(G1966), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n784), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(G1966), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT89), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n773), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G24), .B(G290), .S(G16), .Z(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(G1986), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n484), .A2(G119), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n462), .A2(G107), .ZN(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n809));
  INV_X1    g384(.A(G131), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n807), .B1(new_n808), .B2(new_n809), .C1(new_n810), .C2(new_n487), .ZN(new_n811));
  MUX2_X1   g386(.A(G25), .B(new_n811), .S(G29), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n717), .A2(G6), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n604), .B2(new_n717), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT32), .B(G1981), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n717), .A2(G22), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G166), .B2(new_n717), .ZN(new_n820));
  INV_X1    g395(.A(G1971), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  MUX2_X1   g397(.A(G23), .B(G288), .S(G16), .Z(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT33), .B(G1976), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n816), .A2(new_n817), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n818), .A2(new_n822), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n806), .B(new_n814), .C1(new_n827), .C2(KEYINPUT34), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT84), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT85), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n804), .B1(new_n832), .B2(KEYINPUT36), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(G311));
  OR2_X1    g410(.A1(new_n833), .A2(new_n834), .ZN(G150));
  NAND2_X1  g411(.A1(new_n620), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(new_n519), .ZN(new_n840));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n543), .A2(new_n841), .B1(new_n540), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n559), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n838), .B(new_n848), .Z(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n850), .A2(new_n851), .A3(G860), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n847), .A2(G860), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  XOR2_X1   g430(.A(new_n479), .B(new_n638), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G162), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n490), .A2(new_n493), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n462), .A2(G138), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n474), .B2(new_n475), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT70), .B(KEYINPUT4), .Z(new_n861));
  OAI211_X1 g436(.A(new_n501), .B(KEYINPUT95), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT95), .B1(new_n499), .B2(new_n501), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n744), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n501), .B1(new_n860), .B2(new_n861), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n494), .B1(new_n869), .B2(new_n862), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n743), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n761), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n866), .A2(new_n871), .A3(new_n761), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(KEYINPUT96), .ZN(new_n877));
  INV_X1    g452(.A(new_n732), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n876), .B2(KEYINPUT96), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n484), .A2(G130), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n462), .A2(G118), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(G142), .B2(new_n488), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n641), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n811), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n888));
  INV_X1    g463(.A(new_n875), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n761), .B1(new_n866), .B2(new_n871), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT97), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n874), .A2(new_n892), .A3(new_n875), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n888), .B1(new_n894), .B2(new_n878), .ZN(new_n895));
  AOI211_X1 g470(.A(KEYINPUT98), .B(new_n732), .C1(new_n891), .C2(new_n893), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n880), .B(new_n887), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT99), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n889), .A2(KEYINPUT97), .A3(new_n890), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n892), .B1(new_n874), .B2(new_n875), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n878), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT98), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n894), .A2(new_n888), .A3(new_n878), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n902), .A2(new_n903), .B1(new_n877), .B2(new_n879), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT100), .B1(new_n904), .B2(new_n887), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n880), .B1(new_n895), .B2(new_n896), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n907));
  INV_X1    g482(.A(new_n887), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n857), .B1(new_n898), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n897), .B(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n857), .B1(new_n906), .B2(new_n908), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n911), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n911), .B2(new_n915), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(G395));
  XNOR2_X1  g494(.A(new_n848), .B(new_n631), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n619), .B(G299), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT102), .B1(new_n921), .B2(KEYINPUT41), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n921), .B(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n920), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n604), .B(G290), .ZN(new_n932));
  XNOR2_X1  g507(.A(G303), .B(G288), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n931), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n931), .B2(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n847), .A2(new_n628), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(G295));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n941), .ZN(G331));
  XNOR2_X1  g518(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(G171), .A2(G168), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(G171), .B2(new_n584), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n848), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n848), .A2(new_n947), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n921), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n928), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n949), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n951), .B(new_n936), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G37), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n953), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n950), .B1(new_n957), .B2(new_n928), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n936), .A2(KEYINPUT104), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n934), .B2(new_n935), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n945), .B1(new_n956), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n958), .B2(new_n936), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(new_n961), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n953), .A2(new_n926), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(new_n967), .B2(new_n950), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n944), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT44), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n965), .A2(new_n968), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n965), .B(new_n944), .C1(new_n958), .C2(new_n962), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n971), .A2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1966), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT45), .B1(new_n865), .B2(new_n979), .ZN(new_n980));
  AND4_X1   g555(.A1(G40), .A2(new_n470), .A3(new_n478), .A4(new_n471), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n858), .A2(new_n867), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n979), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n981), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n978), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n858), .B2(new_n867), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT105), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n990), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G2084), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n865), .A2(new_n988), .A3(new_n979), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n981), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n986), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n545), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n986), .A2(new_n995), .A3(G168), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(G8), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT51), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1002), .A3(G8), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1001), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n865), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n470), .A2(G40), .A3(new_n478), .A4(new_n471), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n984), .B2(new_n982), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1008), .A3(new_n775), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT121), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT121), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n992), .A2(new_n981), .A3(new_n994), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT120), .B(G1961), .Z(new_n1016));
  AOI22_X1  g591(.A1(new_n1012), .A2(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n980), .A2(new_n985), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1010), .A2(G2078), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(G301), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n870), .A2(new_n982), .A3(G1384), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n981), .B1(KEYINPUT45), .B2(new_n987), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n821), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n992), .A2(new_n713), .A3(new_n994), .A4(new_n981), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(G166), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n602), .A2(G1981), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n599), .A2(new_n600), .A3(new_n601), .A4(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(KEYINPUT106), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT106), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n602), .A2(new_n1037), .A3(G1981), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT49), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1041), .A3(new_n1038), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n869), .A2(new_n862), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1384), .B1(new_n1043), .B2(new_n858), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1028), .B1(new_n1044), .B2(new_n981), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n547), .A2(G87), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n549), .A2(G49), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(G1976), .A3(new_n1049), .A4(new_n592), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1047), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n981), .A2(new_n865), .A3(new_n979), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  AND4_X1   g629(.A1(G8), .A2(new_n1052), .A3(new_n1054), .A4(new_n1050), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1032), .A2(new_n1046), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT107), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n988), .B1(new_n865), .B2(new_n979), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n983), .A2(new_n988), .A3(new_n979), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n981), .A2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1060), .A2(new_n1062), .A3(G2090), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1971), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1059), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1007), .B1(new_n988), .B2(new_n987), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1066), .B(new_n713), .C1(new_n1044), .C2(new_n988), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1024), .A2(KEYINPUT107), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(G8), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1031), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1021), .A2(new_n1058), .A3(new_n1071), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1004), .A2(new_n1005), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n584), .A2(G8), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n986), .B2(new_n995), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1028), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1075), .B(KEYINPUT63), .C1(new_n1076), .C2(new_n1031), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1057), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1024), .A2(new_n1067), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1028), .B1(new_n1080), .B2(new_n1059), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1031), .B1(new_n1081), .B2(new_n1068), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1075), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1082), .A2(new_n1057), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(new_n1084), .B2(KEYINPUT63), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT108), .ZN(new_n1086));
  INV_X1    g661(.A(G288), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1046), .A2(new_n1053), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1035), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1045), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1055), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT52), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1046), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1032), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1085), .A2(new_n1086), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1071), .A2(new_n1032), .A3(new_n1094), .A4(new_n1075), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1078), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT108), .B1(new_n1102), .B2(new_n1097), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1073), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1058), .A2(new_n1071), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1003), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n999), .B2(KEYINPUT51), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1017), .A2(G301), .A3(new_n1020), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1014), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1013), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1006), .A2(new_n1019), .ZN(new_n1114));
  INV_X1    g689(.A(new_n980), .ZN(new_n1115));
  OR3_X1    g690(.A1(new_n476), .A2(KEYINPUT122), .A3(new_n477), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT122), .B1(new_n476), .B2(new_n477), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(G2105), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n472), .A2(new_n1118), .A3(G40), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT123), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n980), .A2(new_n1122), .A3(new_n1119), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1114), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT124), .B(new_n1114), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1113), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT54), .B(new_n1109), .C1(new_n1128), .C2(G301), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n1130));
  OAI211_X1 g705(.A(G301), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1130), .B1(new_n1132), .B2(new_n1021), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1108), .A2(new_n1129), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n572), .A2(new_n577), .A3(KEYINPUT57), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT112), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n571), .B1(new_n577), .B2(KEYINPUT110), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT110), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n574), .A2(new_n576), .A3(new_n1138), .ZN(new_n1139));
  AOI211_X1 g714(.A(KEYINPUT111), .B(KEYINPUT57), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT111), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n577), .A2(KEYINPUT110), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1142), .A2(new_n572), .A3(new_n1139), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1136), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT113), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT56), .B(G2072), .Z(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT114), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1066), .B1(new_n1044), .B2(new_n988), .ZN(new_n1152));
  INV_X1    g727(.A(G1956), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(KEYINPUT109), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT109), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1151), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT113), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1158), .B(new_n1136), .C1(new_n1140), .C2(new_n1145), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1147), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1157), .B1(new_n1147), .B2(new_n1159), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1052), .A2(G2067), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n1015), .B2(new_n769), .ZN(new_n1163));
  OR3_X1    g738(.A1(new_n1163), .A2(KEYINPUT115), .A3(new_n619), .ZN(new_n1164));
  INV_X1    g739(.A(new_n769), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1007), .B1(new_n1044), .B2(new_n988), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n992), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n620), .B1(new_n1167), .B2(new_n1162), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT115), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1164), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1160), .B1(new_n1161), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1156), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1172), .A2(new_n1154), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT111), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1143), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1158), .B1(new_n1177), .B2(new_n1136), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1159), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1173), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1161), .A2(KEYINPUT61), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1163), .A2(new_n619), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1168), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n619), .A2(KEYINPUT60), .ZN(new_n1187));
  AOI22_X1  g762(.A1(new_n1186), .A2(KEYINPUT60), .B1(new_n1163), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(G1996), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1006), .A2(new_n1008), .A3(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(KEYINPUT58), .B(G1341), .Z(new_n1191));
  NAND2_X1  g766(.A1(new_n1052), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n559), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT117), .B1(new_n1194), .B2(KEYINPUT59), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT117), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT59), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1193), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(KEYINPUT116), .B1(new_n1194), .B2(KEYINPUT59), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT116), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1193), .A2(new_n1200), .A3(new_n1197), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1195), .B(new_n1198), .C1(new_n1199), .C2(new_n1201), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1188), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1171), .B1(new_n1184), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT118), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1134), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g781(.A(KEYINPUT118), .B(new_n1171), .C1(new_n1184), .C2(new_n1203), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1104), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n980), .A2(new_n981), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n761), .B(G1996), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n743), .B(new_n746), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n811), .B(new_n813), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g790(.A(G290), .B(G1986), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1210), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1208), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1209), .B1(new_n761), .B2(new_n1212), .ZN(new_n1219));
  OR3_X1    g794(.A1(new_n1209), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1220));
  OAI21_X1  g795(.A(KEYINPUT46), .B1(new_n1209), .B2(G1996), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g797(.A(new_n1222), .B(KEYINPUT47), .Z(new_n1223));
  INV_X1    g798(.A(new_n813), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n811), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1213), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n744), .A2(new_n746), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1209), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  OR3_X1    g803(.A1(new_n1209), .A2(G1986), .A3(G290), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1229), .ZN(new_n1230));
  OR2_X1    g805(.A1(new_n1230), .A2(KEYINPUT48), .ZN(new_n1231));
  AOI22_X1  g806(.A1(new_n1230), .A2(KEYINPUT48), .B1(new_n1210), .B2(new_n1215), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1228), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1223), .A2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g809(.A(new_n1234), .B(KEYINPUT125), .Z(new_n1235));
  NAND2_X1  g810(.A1(new_n1218), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g811(.A(G319), .ZN(new_n1238));
  NOR3_X1   g812(.A1(G401), .A2(G227), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g813(.A(new_n1239), .B1(new_n706), .B2(new_n707), .ZN(new_n1240));
  XNOR2_X1  g814(.A(new_n1240), .B(KEYINPUT126), .ZN(new_n1241));
  NAND2_X1  g815(.A1(new_n911), .A2(new_n915), .ZN(new_n1242));
  NAND3_X1  g816(.A1(new_n1241), .A2(new_n1242), .A3(new_n970), .ZN(G225));
  INV_X1    g817(.A(G225), .ZN(G308));
endmodule


