

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724;

  AND2_X1 U364 ( .A1(n410), .A2(n392), .ZN(n391) );
  NOR2_X1 U365 ( .A1(n554), .A2(n551), .ZN(n538) );
  NOR2_X1 U366 ( .A1(n520), .A2(n530), .ZN(n663) );
  XNOR2_X1 U367 ( .A(n448), .B(n468), .ZN(n704) );
  XNOR2_X1 U368 ( .A(n445), .B(n429), .ZN(n708) );
  XNOR2_X1 U369 ( .A(n342), .B(n359), .ZN(n372) );
  NAND2_X1 U370 ( .A1(n371), .A2(n367), .ZN(n342) );
  NAND2_X1 U371 ( .A1(n685), .A2(G469), .ZN(n646) );
  AND2_X4 U372 ( .A1(n369), .A2(n390), .ZN(n685) );
  XNOR2_X2 U373 ( .A(n428), .B(G143), .ZN(n445) );
  XNOR2_X2 U374 ( .A(n474), .B(n473), .ZN(n481) );
  INV_X1 U375 ( .A(G953), .ZN(n710) );
  AND2_X2 U376 ( .A1(n381), .A2(n382), .ZN(n380) );
  XNOR2_X2 U377 ( .A(n545), .B(n544), .ZN(n560) );
  OR2_X2 U378 ( .A1(n643), .A2(G902), .ZN(n400) );
  XNOR2_X2 U379 ( .A(n510), .B(n509), .ZN(n576) );
  NAND2_X1 U380 ( .A1(n355), .A2(n594), .ZN(n413) );
  NAND2_X1 U381 ( .A1(n385), .A2(n384), .ZN(n379) );
  OR2_X1 U382 ( .A1(n580), .A2(n357), .ZN(n569) );
  XNOR2_X1 U383 ( .A(n562), .B(n561), .ZN(n580) );
  XNOR2_X1 U384 ( .A(n462), .B(n461), .ZN(n530) );
  XNOR2_X1 U385 ( .A(n389), .B(n387), .ZN(n609) );
  XOR2_X1 U386 ( .A(G146), .B(G125), .Z(n468) );
  OR2_X2 U387 ( .A1(n563), .A2(n605), .ZN(n577) );
  XNOR2_X1 U388 ( .A(n708), .B(n418), .ZN(n474) );
  XNOR2_X1 U389 ( .A(KEYINPUT66), .B(G101), .ZN(n418) );
  XNOR2_X1 U390 ( .A(n692), .B(KEYINPUT75), .ZN(n473) );
  XNOR2_X1 U391 ( .A(n447), .B(G140), .ZN(n448) );
  XOR2_X1 U392 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n447) );
  INV_X1 U393 ( .A(n671), .ZN(n411) );
  XNOR2_X1 U394 ( .A(KEYINPUT85), .B(KEYINPUT0), .ZN(n561) );
  NOR2_X1 U395 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U396 ( .A(n388), .B(n483), .ZN(n387) );
  OR2_X1 U397 ( .A1(n687), .A2(G902), .ZN(n389) );
  NAND2_X1 U398 ( .A1(n685), .A2(G472), .ZN(n370) );
  NOR2_X1 U399 ( .A1(n722), .A2(n723), .ZN(n534) );
  INV_X1 U400 ( .A(n721), .ZN(n368) );
  OR2_X1 U401 ( .A1(G237), .A2(G902), .ZN(n506) );
  AND2_X1 U402 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U403 ( .A(n386), .B(KEYINPUT88), .ZN(n595) );
  XNOR2_X1 U404 ( .A(G902), .B(KEYINPUT15), .ZN(n386) );
  INV_X1 U405 ( .A(G469), .ZN(n399) );
  XNOR2_X1 U406 ( .A(n481), .B(n475), .ZN(n675) );
  NOR2_X1 U407 ( .A1(n516), .A2(n513), .ZN(n514) );
  XNOR2_X1 U408 ( .A(KEYINPUT6), .B(n576), .ZN(n587) );
  NAND2_X1 U409 ( .A1(n568), .A2(n358), .ZN(n357) );
  INV_X1 U410 ( .A(n610), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n495), .B(n494), .ZN(n687) );
  NAND2_X1 U412 ( .A1(n409), .A2(n408), .ZN(n390) );
  INV_X1 U413 ( .A(KEYINPUT76), .ZN(n375) );
  NOR2_X1 U414 ( .A1(n402), .A2(n401), .ZN(n378) );
  XNOR2_X1 U415 ( .A(G116), .B(KEYINPUT72), .ZN(n423) );
  XNOR2_X1 U416 ( .A(G113), .B(G119), .ZN(n425) );
  XOR2_X1 U417 ( .A(G134), .B(n449), .Z(n477) );
  XNOR2_X1 U418 ( .A(G146), .B(G137), .ZN(n430) );
  INV_X1 U419 ( .A(KEYINPUT4), .ZN(n429) );
  XNOR2_X1 U420 ( .A(n398), .B(n397), .ZN(n463) );
  XNOR2_X1 U421 ( .A(n424), .B(KEYINPUT73), .ZN(n397) );
  XNOR2_X1 U422 ( .A(n425), .B(n423), .ZN(n398) );
  INV_X1 U423 ( .A(KEYINPUT3), .ZN(n424) );
  XOR2_X1 U424 ( .A(G137), .B(KEYINPUT70), .Z(n490) );
  AND2_X1 U425 ( .A1(n550), .A2(n541), .ZN(n371) );
  AND2_X1 U426 ( .A1(n542), .A2(n368), .ZN(n367) );
  INV_X1 U427 ( .A(KEYINPUT48), .ZN(n359) );
  XOR2_X1 U428 ( .A(G146), .B(G140), .Z(n479) );
  XNOR2_X1 U429 ( .A(n467), .B(n365), .ZN(n470) );
  INV_X1 U430 ( .A(n468), .ZN(n365) );
  XNOR2_X1 U431 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n465) );
  NAND2_X1 U432 ( .A1(n621), .A2(n620), .ZN(n625) );
  XNOR2_X1 U433 ( .A(n543), .B(n356), .ZN(n621) );
  INV_X1 U434 ( .A(KEYINPUT38), .ZN(n356) );
  INV_X1 U435 ( .A(KEYINPUT33), .ZN(n403) );
  INV_X1 U436 ( .A(n587), .ZN(n405) );
  AND2_X1 U437 ( .A1(n496), .A2(G217), .ZN(n388) );
  INV_X1 U438 ( .A(KEYINPUT45), .ZN(n412) );
  AND2_X1 U439 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U440 ( .A(G104), .B(G110), .Z(n472) );
  XNOR2_X1 U441 ( .A(n463), .B(n396), .ZN(n690) );
  XNOR2_X1 U442 ( .A(n464), .B(G122), .ZN(n396) );
  XOR2_X1 U443 ( .A(KEYINPUT16), .B(KEYINPUT77), .Z(n464) );
  XNOR2_X1 U444 ( .A(G110), .B(KEYINPUT91), .ZN(n484) );
  INV_X1 U445 ( .A(n595), .ZN(n392) );
  XNOR2_X1 U446 ( .A(G122), .B(KEYINPUT7), .ZN(n437) );
  XOR2_X1 U447 ( .A(KEYINPUT9), .B(KEYINPUT98), .Z(n438) );
  XNOR2_X1 U448 ( .A(G116), .B(G134), .ZN(n436) );
  XNOR2_X1 U449 ( .A(n459), .B(n458), .ZN(n680) );
  XNOR2_X1 U450 ( .A(n457), .B(n456), .ZN(n458) );
  INV_X1 U451 ( .A(G113), .ZN(n456) );
  NOR2_X1 U452 ( .A1(n580), .A2(KEYINPUT34), .ZN(n384) );
  INV_X1 U453 ( .A(KEYINPUT19), .ZN(n544) );
  INV_X1 U454 ( .A(n609), .ZN(n570) );
  INV_X1 U455 ( .A(KEYINPUT123), .ZN(n416) );
  XNOR2_X1 U456 ( .A(n533), .B(KEYINPUT42), .ZN(n722) );
  XNOR2_X1 U457 ( .A(n522), .B(KEYINPUT40), .ZN(n723) );
  XNOR2_X1 U458 ( .A(n579), .B(n366), .ZN(n668) );
  INV_X1 U459 ( .A(KEYINPUT31), .ZN(n366) );
  NOR2_X1 U460 ( .A1(n560), .A2(n546), .ZN(n664) );
  NAND2_X1 U461 ( .A1(n607), .A2(n527), .ZN(n395) );
  NOR2_X1 U462 ( .A1(n589), .A2(n588), .ZN(n650) );
  XNOR2_X1 U463 ( .A(n370), .B(n351), .ZN(n422) );
  XNOR2_X1 U464 ( .A(n686), .B(n362), .ZN(n688) );
  XNOR2_X1 U465 ( .A(n687), .B(KEYINPUT124), .ZN(n362) );
  NOR2_X1 U466 ( .A1(n414), .A2(n689), .ZN(G63) );
  XNOR2_X1 U467 ( .A(n417), .B(n415), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n684), .B(n416), .ZN(n415) );
  NAND2_X1 U469 ( .A1(n685), .A2(G478), .ZN(n417) );
  INV_X1 U470 ( .A(KEYINPUT56), .ZN(n363) );
  NOR2_X1 U471 ( .A1(n639), .A2(n638), .ZN(n642) );
  OR2_X1 U472 ( .A1(n563), .A2(n567), .ZN(n343) );
  NOR2_X1 U473 ( .A1(n699), .A2(n709), .ZN(n344) );
  NOR2_X1 U474 ( .A1(n585), .A2(n570), .ZN(n345) );
  OR2_X1 U475 ( .A1(n343), .A2(n570), .ZN(n346) );
  XOR2_X1 U476 ( .A(KEYINPUT30), .B(n511), .Z(n347) );
  AND2_X1 U477 ( .A1(G210), .A2(n506), .ZN(n348) );
  AND2_X1 U478 ( .A1(n673), .A2(n411), .ZN(n349) );
  OR2_X1 U479 ( .A1(n605), .A2(n395), .ZN(n350) );
  XOR2_X1 U480 ( .A(n435), .B(n434), .Z(n351) );
  XNOR2_X1 U481 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n352) );
  XNOR2_X1 U482 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n353) );
  XOR2_X1 U483 ( .A(KEYINPUT60), .B(KEYINPUT122), .Z(n354) );
  XNOR2_X2 U484 ( .A(n581), .B(KEYINPUT1), .ZN(n563) );
  NAND2_X1 U485 ( .A1(n675), .A2(n595), .ZN(n476) );
  NOR2_X1 U486 ( .A1(n521), .A2(n666), .ZN(n522) );
  NAND2_X1 U487 ( .A1(n543), .A2(n620), .ZN(n545) );
  XNOR2_X2 U488 ( .A(n476), .B(n348), .ZN(n543) );
  AND2_X2 U489 ( .A1(n373), .A2(n377), .ZN(n355) );
  NAND2_X1 U490 ( .A1(n347), .A2(n512), .ZN(n516) );
  XNOR2_X1 U491 ( .A(n361), .B(n354), .ZN(G60) );
  NAND2_X1 U492 ( .A1(n683), .A2(n596), .ZN(n361) );
  XNOR2_X1 U493 ( .A(n376), .B(n375), .ZN(n374) );
  XNOR2_X1 U494 ( .A(n364), .B(n363), .ZN(G51) );
  NAND2_X1 U495 ( .A1(n678), .A2(n596), .ZN(n364) );
  NAND2_X1 U496 ( .A1(n699), .A2(n598), .ZN(n393) );
  XNOR2_X1 U497 ( .A(n394), .B(n353), .ZN(n724) );
  NAND2_X1 U498 ( .A1(n668), .A2(n653), .ZN(n583) );
  AND2_X2 U499 ( .A1(n393), .A2(n391), .ZN(n369) );
  NOR2_X2 U500 ( .A1(n647), .A2(n689), .ZN(n649) );
  XNOR2_X1 U501 ( .A(n505), .B(KEYINPUT78), .ZN(n512) );
  XOR2_X2 U502 ( .A(KEYINPUT69), .B(G131), .Z(n449) );
  NAND2_X1 U503 ( .A1(n372), .A2(n349), .ZN(n709) );
  NAND2_X1 U504 ( .A1(n374), .A2(n572), .ZN(n373) );
  NAND2_X1 U505 ( .A1(n402), .A2(n401), .ZN(n376) );
  XNOR2_X1 U506 ( .A(n378), .B(n573), .ZN(n377) );
  NAND2_X2 U507 ( .A1(n380), .A2(n379), .ZN(n566) );
  NAND2_X1 U508 ( .A1(n600), .A2(KEYINPUT34), .ZN(n381) );
  AND2_X1 U509 ( .A1(n383), .A2(n565), .ZN(n382) );
  NAND2_X1 U510 ( .A1(n580), .A2(KEYINPUT34), .ZN(n383) );
  INV_X1 U511 ( .A(n600), .ZN(n385) );
  XNOR2_X2 U512 ( .A(n404), .B(n403), .ZN(n600) );
  INV_X1 U513 ( .A(n699), .ZN(n409) );
  NOR2_X1 U514 ( .A1(n585), .A2(n346), .ZN(n394) );
  NAND2_X1 U515 ( .A1(n724), .A2(n657), .ZN(n575) );
  NOR2_X1 U516 ( .A1(n580), .A2(n350), .ZN(n582) );
  NOR2_X1 U517 ( .A1(n709), .A2(n598), .ZN(n408) );
  XNOR2_X2 U518 ( .A(n400), .B(n399), .ZN(n581) );
  XNOR2_X1 U519 ( .A(n481), .B(n420), .ZN(n643) );
  INV_X1 U520 ( .A(KEYINPUT44), .ZN(n401) );
  XNOR2_X1 U521 ( .A(n402), .B(G122), .ZN(G24) );
  XNOR2_X2 U522 ( .A(n566), .B(n352), .ZN(n402) );
  NAND2_X1 U523 ( .A1(n406), .A2(n405), .ZN(n404) );
  XNOR2_X1 U524 ( .A(n577), .B(n407), .ZN(n406) );
  INV_X1 U525 ( .A(KEYINPUT100), .ZN(n407) );
  NAND2_X1 U526 ( .A1(n709), .A2(n598), .ZN(n410) );
  XNOR2_X2 U527 ( .A(n413), .B(n412), .ZN(n699) );
  XOR2_X1 U528 ( .A(n431), .B(n430), .Z(n419) );
  XOR2_X1 U529 ( .A(n705), .B(n480), .Z(n420) );
  XOR2_X1 U530 ( .A(n645), .B(n644), .Z(n421) );
  BUF_X1 U531 ( .A(n600), .Z(n629) );
  INV_X1 U532 ( .A(G472), .ZN(n508) );
  XNOR2_X1 U533 ( .A(n460), .B(G475), .ZN(n461) );
  XNOR2_X1 U534 ( .A(n508), .B(KEYINPUT94), .ZN(n509) );
  XNOR2_X1 U535 ( .A(n680), .B(n679), .ZN(n681) );
  INV_X1 U536 ( .A(n689), .ZN(n596) );
  XNOR2_X1 U537 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U538 ( .A1(n422), .A2(n596), .ZN(n597) );
  NOR2_X1 U539 ( .A1(G952), .A2(n710), .ZN(n689) );
  XNOR2_X1 U540 ( .A(n642), .B(n641), .ZN(G75) );
  XOR2_X1 U541 ( .A(KEYINPUT86), .B(KEYINPUT62), .Z(n435) );
  XOR2_X1 U542 ( .A(n477), .B(n463), .Z(n427) );
  NOR2_X1 U543 ( .A1(G953), .A2(G237), .ZN(n452) );
  NAND2_X1 U544 ( .A1(n452), .A2(G210), .ZN(n426) );
  XNOR2_X1 U545 ( .A(n427), .B(n426), .ZN(n433) );
  XNOR2_X2 U546 ( .A(G128), .B(KEYINPUT64), .ZN(n428) );
  XOR2_X1 U547 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n431) );
  XNOR2_X1 U548 ( .A(n474), .B(n419), .ZN(n432) );
  XNOR2_X1 U549 ( .A(n433), .B(n432), .ZN(n507) );
  XOR2_X1 U550 ( .A(n507), .B(KEYINPUT108), .Z(n434) );
  XNOR2_X1 U551 ( .A(n436), .B(G107), .ZN(n440) );
  XNOR2_X1 U552 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U553 ( .A(n440), .B(n439), .Z(n443) );
  NAND2_X1 U554 ( .A1(G234), .A2(n710), .ZN(n441) );
  XOR2_X1 U555 ( .A(KEYINPUT8), .B(n441), .Z(n491) );
  NAND2_X1 U556 ( .A1(G217), .A2(n491), .ZN(n442) );
  XNOR2_X1 U557 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U558 ( .A(n445), .B(n444), .ZN(n684) );
  NOR2_X1 U559 ( .A1(G902), .A2(n684), .ZN(n446) );
  XOR2_X1 U560 ( .A(G478), .B(n446), .Z(n520) );
  XNOR2_X1 U561 ( .A(G143), .B(n449), .ZN(n450) );
  XNOR2_X1 U562 ( .A(n450), .B(G104), .ZN(n451) );
  XOR2_X1 U563 ( .A(n704), .B(n451), .Z(n454) );
  NAND2_X1 U564 ( .A1(G214), .A2(n452), .ZN(n453) );
  XNOR2_X1 U565 ( .A(n454), .B(n453), .ZN(n459) );
  XOR2_X1 U566 ( .A(G122), .B(KEYINPUT11), .Z(n455) );
  XNOR2_X1 U567 ( .A(KEYINPUT12), .B(n455), .ZN(n457) );
  NOR2_X1 U568 ( .A1(G902), .A2(n680), .ZN(n462) );
  XNOR2_X1 U569 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n460) );
  NAND2_X1 U570 ( .A1(n520), .A2(n530), .ZN(n669) );
  XOR2_X1 U571 ( .A(KEYINPUT89), .B(KEYINPUT80), .Z(n466) );
  XNOR2_X1 U572 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U573 ( .A1(G224), .A2(n710), .ZN(n469) );
  XNOR2_X1 U574 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U575 ( .A(n690), .B(n471), .ZN(n475) );
  XNOR2_X1 U576 ( .A(G107), .B(n472), .ZN(n692) );
  INV_X1 U577 ( .A(n621), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n477), .B(n490), .ZN(n705) );
  NAND2_X1 U579 ( .A1(G227), .A2(n710), .ZN(n478) );
  XNOR2_X1 U580 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U581 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n483) );
  NAND2_X1 U582 ( .A1(n595), .A2(G234), .ZN(n482) );
  XNOR2_X1 U583 ( .A(KEYINPUT20), .B(n482), .ZN(n496) );
  XOR2_X1 U584 ( .A(KEYINPUT79), .B(KEYINPUT24), .Z(n485) );
  XNOR2_X1 U585 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U586 ( .A(n704), .B(n486), .ZN(n495) );
  XOR2_X1 U587 ( .A(KEYINPUT74), .B(KEYINPUT23), .Z(n488) );
  XNOR2_X1 U588 ( .A(G128), .B(G119), .ZN(n487) );
  XNOR2_X1 U589 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U590 ( .A(n490), .B(n489), .Z(n493) );
  NAND2_X1 U591 ( .A1(G221), .A2(n491), .ZN(n492) );
  XNOR2_X1 U592 ( .A(n493), .B(n492), .ZN(n494) );
  NAND2_X1 U593 ( .A1(n496), .A2(G221), .ZN(n497) );
  XNOR2_X1 U594 ( .A(n497), .B(KEYINPUT21), .ZN(n610) );
  XOR2_X1 U595 ( .A(KEYINPUT14), .B(KEYINPUT90), .Z(n499) );
  NAND2_X1 U596 ( .A1(G234), .A2(G237), .ZN(n498) );
  XOR2_X1 U597 ( .A(n499), .B(n498), .Z(n500) );
  NAND2_X1 U598 ( .A1(G952), .A2(n500), .ZN(n636) );
  NOR2_X1 U599 ( .A1(G953), .A2(n636), .ZN(n558) );
  AND2_X1 U600 ( .A1(n500), .A2(G953), .ZN(n501) );
  NAND2_X1 U601 ( .A1(G902), .A2(n501), .ZN(n556) );
  NOR2_X1 U602 ( .A1(n556), .A2(G900), .ZN(n502) );
  NOR2_X1 U603 ( .A1(n558), .A2(n502), .ZN(n503) );
  NOR2_X1 U604 ( .A1(n610), .A2(n503), .ZN(n523) );
  NAND2_X1 U605 ( .A1(n570), .A2(n523), .ZN(n504) );
  NOR2_X1 U606 ( .A1(n581), .A2(n504), .ZN(n505) );
  NAND2_X1 U607 ( .A1(G214), .A2(n506), .ZN(n620) );
  NOR2_X1 U608 ( .A1(G902), .A2(n507), .ZN(n510) );
  NAND2_X1 U609 ( .A1(n620), .A2(n576), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n514), .B(KEYINPUT39), .ZN(n521) );
  NOR2_X1 U611 ( .A1(n669), .A2(n521), .ZN(n671) );
  INV_X1 U612 ( .A(n520), .ZN(n529) );
  NOR2_X1 U613 ( .A1(n529), .A2(n530), .ZN(n515) );
  XNOR2_X1 U614 ( .A(n515), .B(KEYINPUT101), .ZN(n564) );
  INV_X1 U615 ( .A(n543), .ZN(n554) );
  NOR2_X1 U616 ( .A1(n554), .A2(n516), .ZN(n517) );
  XNOR2_X1 U617 ( .A(n517), .B(KEYINPUT103), .ZN(n518) );
  NOR2_X1 U618 ( .A1(n564), .A2(n518), .ZN(n519) );
  XNOR2_X1 U619 ( .A(KEYINPUT104), .B(n519), .ZN(n721) );
  INV_X1 U620 ( .A(n663), .ZN(n666) );
  XNOR2_X1 U621 ( .A(KEYINPUT71), .B(n523), .ZN(n524) );
  NOR2_X1 U622 ( .A1(n570), .A2(n524), .ZN(n535) );
  NAND2_X1 U623 ( .A1(n576), .A2(n535), .ZN(n525) );
  XNOR2_X1 U624 ( .A(n525), .B(KEYINPUT105), .ZN(n526) );
  XNOR2_X1 U625 ( .A(KEYINPUT28), .B(n526), .ZN(n528) );
  INV_X1 U626 ( .A(n581), .ZN(n527) );
  NAND2_X1 U627 ( .A1(n528), .A2(n527), .ZN(n546) );
  NAND2_X1 U628 ( .A1(n530), .A2(n529), .ZN(n623) );
  NOR2_X1 U629 ( .A1(n623), .A2(n625), .ZN(n532) );
  XNOR2_X1 U630 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n531) );
  XNOR2_X1 U631 ( .A(n532), .B(n531), .ZN(n619) );
  NOR2_X1 U632 ( .A1(n546), .A2(n619), .ZN(n533) );
  XNOR2_X1 U633 ( .A(n534), .B(KEYINPUT46), .ZN(n542) );
  NAND2_X1 U634 ( .A1(n663), .A2(n535), .ZN(n536) );
  NOR2_X1 U635 ( .A1(n587), .A2(n536), .ZN(n537) );
  NAND2_X1 U636 ( .A1(n537), .A2(n620), .ZN(n551) );
  XNOR2_X1 U637 ( .A(KEYINPUT36), .B(n538), .ZN(n539) );
  INV_X1 U638 ( .A(n563), .ZN(n589) );
  NAND2_X1 U639 ( .A1(n539), .A2(n589), .ZN(n540) );
  XNOR2_X1 U640 ( .A(n540), .B(KEYINPUT107), .ZN(n717) );
  INV_X1 U641 ( .A(n717), .ZN(n541) );
  INV_X1 U642 ( .A(n669), .ZN(n659) );
  NOR2_X1 U643 ( .A1(n659), .A2(n663), .ZN(n547) );
  XNOR2_X1 U644 ( .A(n547), .B(KEYINPUT99), .ZN(n624) );
  NAND2_X1 U645 ( .A1(n664), .A2(n624), .ZN(n548) );
  NOR2_X1 U646 ( .A1(KEYINPUT67), .A2(n548), .ZN(n549) );
  XNOR2_X1 U647 ( .A(n549), .B(KEYINPUT47), .ZN(n550) );
  OR2_X1 U648 ( .A1(n551), .A2(n589), .ZN(n552) );
  XNOR2_X1 U649 ( .A(n552), .B(KEYINPUT43), .ZN(n553) );
  XNOR2_X1 U650 ( .A(n553), .B(KEYINPUT102), .ZN(n555) );
  NAND2_X1 U651 ( .A1(n555), .A2(n554), .ZN(n673) );
  NOR2_X1 U652 ( .A1(G898), .A2(n556), .ZN(n557) );
  NOR2_X1 U653 ( .A1(n558), .A2(n557), .ZN(n559) );
  OR2_X1 U654 ( .A1(n610), .A2(n609), .ZN(n605) );
  INV_X1 U655 ( .A(n564), .ZN(n565) );
  XOR2_X1 U656 ( .A(KEYINPUT82), .B(n587), .Z(n567) );
  INV_X1 U657 ( .A(n623), .ZN(n568) );
  XNOR2_X1 U658 ( .A(KEYINPUT22), .B(n569), .ZN(n585) );
  NOR2_X1 U659 ( .A1(n589), .A2(n576), .ZN(n571) );
  NAND2_X1 U660 ( .A1(n345), .A2(n571), .ZN(n657) );
  INV_X1 U661 ( .A(n575), .ZN(n572) );
  INV_X1 U662 ( .A(KEYINPUT84), .ZN(n573) );
  NAND2_X1 U663 ( .A1(KEYINPUT76), .A2(n401), .ZN(n574) );
  NAND2_X1 U664 ( .A1(n575), .A2(n574), .ZN(n593) );
  INV_X1 U665 ( .A(n580), .ZN(n578) );
  INV_X1 U666 ( .A(n576), .ZN(n607) );
  NOR2_X1 U667 ( .A1(n607), .A2(n577), .ZN(n616) );
  NAND2_X1 U668 ( .A1(n578), .A2(n616), .ZN(n579) );
  XNOR2_X1 U669 ( .A(n582), .B(KEYINPUT95), .ZN(n653) );
  XNOR2_X1 U670 ( .A(KEYINPUT96), .B(n583), .ZN(n584) );
  NAND2_X1 U671 ( .A1(n584), .A2(n624), .ZN(n591) );
  NOR2_X1 U672 ( .A1(n585), .A2(n609), .ZN(n586) );
  NAND2_X1 U673 ( .A1(n587), .A2(n586), .ZN(n588) );
  INV_X1 U674 ( .A(n650), .ZN(n590) );
  XNOR2_X1 U675 ( .A(n597), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U676 ( .A1(n344), .A2(KEYINPUT83), .ZN(n599) );
  INV_X1 U677 ( .A(KEYINPUT2), .ZN(n598) );
  XNOR2_X1 U678 ( .A(n599), .B(n598), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n619), .A2(n629), .ZN(n601) );
  XNOR2_X1 U680 ( .A(KEYINPUT118), .B(n601), .ZN(n602) );
  NOR2_X1 U681 ( .A1(G953), .A2(n602), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n639) );
  NAND2_X1 U683 ( .A1(n563), .A2(n605), .ZN(n606) );
  XNOR2_X1 U684 ( .A(KEYINPUT50), .B(n606), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U687 ( .A(KEYINPUT49), .B(n611), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U689 ( .A(KEYINPUT115), .B(n614), .Z(n615) );
  NOR2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U691 ( .A(KEYINPUT51), .B(n617), .Z(n618) );
  NOR2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n632) );
  NOR2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n628) );
  INV_X1 U695 ( .A(n624), .ZN(n626) );
  NOR2_X1 U696 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U697 ( .A1(n628), .A2(n627), .ZN(n630) );
  NOR2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U700 ( .A(n633), .B(KEYINPUT52), .ZN(n634) );
  XNOR2_X1 U701 ( .A(KEYINPUT116), .B(n634), .ZN(n635) );
  NOR2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U703 ( .A(n637), .B(KEYINPUT117), .Z(n638) );
  INV_X1 U704 ( .A(KEYINPUT119), .ZN(n640) );
  XNOR2_X1 U705 ( .A(n640), .B(KEYINPUT53), .ZN(n641) );
  XNOR2_X1 U706 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n645) );
  XNOR2_X1 U707 ( .A(n643), .B(KEYINPUT57), .ZN(n644) );
  XNOR2_X1 U708 ( .A(n646), .B(n421), .ZN(n647) );
  INV_X1 U709 ( .A(KEYINPUT121), .ZN(n648) );
  XNOR2_X1 U710 ( .A(n649), .B(n648), .ZN(G54) );
  XNOR2_X1 U711 ( .A(G101), .B(n650), .ZN(n651) );
  XNOR2_X1 U712 ( .A(n651), .B(KEYINPUT109), .ZN(G3) );
  NOR2_X1 U713 ( .A1(n666), .A2(n653), .ZN(n652) );
  XOR2_X1 U714 ( .A(G104), .B(n652), .Z(G6) );
  NOR2_X1 U715 ( .A1(n669), .A2(n653), .ZN(n655) );
  XNOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n654) );
  XNOR2_X1 U717 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U718 ( .A(G107), .B(n656), .ZN(G9) );
  XNOR2_X1 U719 ( .A(G110), .B(KEYINPUT110), .ZN(n658) );
  XNOR2_X1 U720 ( .A(n658), .B(n657), .ZN(G12) );
  XOR2_X1 U721 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n661) );
  NAND2_X1 U722 ( .A1(n664), .A2(n659), .ZN(n660) );
  XNOR2_X1 U723 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U724 ( .A(G128), .B(n662), .Z(G30) );
  NAND2_X1 U725 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U726 ( .A(n665), .B(G146), .ZN(G48) );
  NOR2_X1 U727 ( .A1(n666), .A2(n668), .ZN(n667) );
  XOR2_X1 U728 ( .A(G113), .B(n667), .Z(G15) );
  NOR2_X1 U729 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U730 ( .A(G116), .B(n670), .Z(G18) );
  XOR2_X1 U731 ( .A(G134), .B(n671), .Z(n672) );
  XNOR2_X1 U732 ( .A(KEYINPUT114), .B(n672), .ZN(G36) );
  XNOR2_X1 U733 ( .A(G140), .B(n673), .ZN(G42) );
  NAND2_X1 U734 ( .A1(n685), .A2(G210), .ZN(n677) );
  XOR2_X1 U735 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n674) );
  XNOR2_X1 U736 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U737 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U738 ( .A1(n685), .A2(G475), .ZN(n682) );
  XOR2_X1 U739 ( .A(KEYINPUT59), .B(KEYINPUT87), .Z(n679) );
  NAND2_X1 U740 ( .A1(n685), .A2(G217), .ZN(n686) );
  NOR2_X1 U741 ( .A1(n689), .A2(n688), .ZN(G66) );
  XOR2_X1 U742 ( .A(G101), .B(n690), .Z(n691) );
  XNOR2_X1 U743 ( .A(n692), .B(n691), .ZN(n694) );
  NOR2_X1 U744 ( .A1(G898), .A2(n710), .ZN(n693) );
  NOR2_X1 U745 ( .A1(n694), .A2(n693), .ZN(n703) );
  INV_X1 U746 ( .A(G898), .ZN(n698) );
  NAND2_X1 U747 ( .A1(G224), .A2(G953), .ZN(n695) );
  XNOR2_X1 U748 ( .A(n695), .B(KEYINPUT125), .ZN(n696) );
  XNOR2_X1 U749 ( .A(n696), .B(KEYINPUT61), .ZN(n697) );
  NOR2_X1 U750 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U751 ( .A1(G953), .A2(n699), .ZN(n700) );
  NOR2_X1 U752 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U753 ( .A(n703), .B(n702), .Z(G69) );
  XNOR2_X1 U754 ( .A(n704), .B(KEYINPUT126), .ZN(n706) );
  XNOR2_X1 U755 ( .A(n705), .B(n706), .ZN(n707) );
  XNOR2_X1 U756 ( .A(n708), .B(n707), .ZN(n712) );
  XNOR2_X1 U757 ( .A(n709), .B(n712), .ZN(n711) );
  NAND2_X1 U758 ( .A1(n711), .A2(n710), .ZN(n716) );
  XNOR2_X1 U759 ( .A(G227), .B(n712), .ZN(n713) );
  NAND2_X1 U760 ( .A1(n713), .A2(G900), .ZN(n714) );
  NAND2_X1 U761 ( .A1(n714), .A2(G953), .ZN(n715) );
  NAND2_X1 U762 ( .A1(n716), .A2(n715), .ZN(G72) );
  XOR2_X1 U763 ( .A(KEYINPUT113), .B(KEYINPUT37), .Z(n719) );
  XNOR2_X1 U764 ( .A(n717), .B(G125), .ZN(n718) );
  XNOR2_X1 U765 ( .A(n719), .B(n718), .ZN(G27) );
  XOR2_X1 U766 ( .A(G143), .B(KEYINPUT112), .Z(n720) );
  XNOR2_X1 U767 ( .A(n721), .B(n720), .ZN(G45) );
  XOR2_X1 U768 ( .A(G137), .B(n722), .Z(G39) );
  XOR2_X1 U769 ( .A(n723), .B(G131), .Z(G33) );
  XNOR2_X1 U770 ( .A(n724), .B(G119), .ZN(G21) );
endmodule

