//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994;
  INV_X1    g000(.A(G230gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G57gat), .B(G64gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G71gat), .ZN(new_n208));
  INV_X1    g007(.A(G78gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G71gat), .A2(G78gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n207), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n211), .B(new_n210), .C1(new_n206), .C2(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G85gat), .ZN(new_n219));
  INV_X1    g018(.A(G92gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(G85gat), .A3(G92gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT98), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT98), .A2(G99gat), .A3(G106gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT8), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n220), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT99), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n225), .ZN(new_n235));
  INV_X1    g034(.A(new_n225), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT99), .B1(new_n236), .B2(new_n232), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n238), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n231), .A2(new_n238), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n231), .A2(new_n238), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n217), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT10), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n218), .A2(KEYINPUT10), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT100), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n242), .B2(new_n243), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n239), .A2(KEYINPUT100), .A3(new_n240), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n205), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n241), .A2(new_n244), .A3(new_n204), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G120gat), .B(G148gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT105), .ZN(new_n255));
  INV_X1    g054(.A(G176gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G204gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n259), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(G113gat), .B2(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(G113gat), .A2(G120gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G113gat), .ZN(new_n272));
  INV_X1    g071(.A(G120gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(new_n265), .A3(new_n267), .ZN(new_n275));
  AND2_X1   g074(.A1(G127gat), .A2(G134gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(G127gat), .A2(G134gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n275), .A2(KEYINPUT71), .A3(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(KEYINPUT72), .A2(G120gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(KEYINPUT72), .A2(G120gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(G113gat), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n266), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n271), .A2(new_n279), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  AND2_X1   g085(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(KEYINPUT70), .B(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n298));
  INV_X1    g097(.A(G169gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n256), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n297), .B(new_n298), .C1(KEYINPUT26), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n291), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n304));
  OAI211_X1 g103(.A(G183gat), .B(G190gat), .C1(KEYINPUT67), .C2(KEYINPUT24), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G183gat), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n309), .A2(new_n286), .A3(KEYINPUT68), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT68), .B1(new_n309), .B2(new_n286), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n305), .B(new_n308), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n300), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n314), .A2(G176gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(new_n299), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n312), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT64), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n320), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n302), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT64), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n286), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n325), .A2(new_n320), .A3(KEYINPUT24), .A4(new_n302), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n256), .A2(KEYINPUT23), .ZN(new_n329));
  OR2_X1    g128(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n292), .B1(new_n293), .B2(KEYINPUT23), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n328), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n317), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n315), .A2(new_n337), .A3(KEYINPUT66), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n327), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  AOI211_X1 g138(.A(new_n304), .B(new_n319), .C1(new_n316), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n316), .ZN(new_n341));
  INV_X1    g140(.A(new_n319), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT69), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n285), .B(new_n303), .C1(new_n340), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n332), .A2(new_n328), .A3(new_n333), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT66), .B1(new_n315), .B2(new_n337), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT25), .B1(new_n349), .B2(new_n327), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n304), .B1(new_n350), .B2(new_n319), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n319), .B1(new_n339), .B2(new_n316), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT69), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n354), .A2(KEYINPUT73), .A3(new_n285), .A4(new_n303), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n303), .B1(new_n340), .B2(new_n343), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n280), .A2(new_n281), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n284), .B(new_n270), .C1(new_n357), .C2(new_n272), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n269), .A2(new_n264), .A3(new_n270), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT71), .B1(new_n275), .B2(new_n278), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n355), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT33), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G15gat), .B(G43gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(new_n208), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(G99gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n367), .B1(new_n372), .B2(KEYINPUT33), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n366), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n366), .A2(KEYINPUT74), .A3(new_n374), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n373), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n346), .A2(new_n355), .A3(new_n362), .A4(new_n364), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n380), .B(KEYINPUT34), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n381), .A2(new_n373), .A3(new_n377), .A4(new_n378), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(KEYINPUT75), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT36), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n379), .A2(new_n387), .A3(new_n382), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(KEYINPUT36), .A3(new_n384), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT77), .ZN(new_n393));
  INV_X1    g192(.A(G64gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(new_n220), .ZN(new_n396));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n356), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400));
  INV_X1    g199(.A(new_n303), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n352), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n397), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT76), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n405), .A3(new_n397), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G197gat), .B(G204gat), .ZN(new_n408));
  INV_X1    g207(.A(G211gat), .ZN(new_n409));
  INV_X1    g208(.A(G218gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n408), .B1(KEYINPUT22), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G211gat), .B(G218gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n398), .A2(KEYINPUT29), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n356), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n398), .B(new_n303), .C1(new_n350), .C2(new_n319), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n414), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n396), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT37), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n402), .A2(new_n405), .A3(new_n397), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n405), .B1(new_n402), .B2(new_n397), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n414), .B1(new_n426), .B2(new_n399), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n416), .A2(KEYINPUT37), .A3(new_n421), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n396), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n422), .B1(new_n431), .B2(KEYINPUT38), .ZN(new_n432));
  XNOR2_X1  g231(.A(G155gat), .B(G162gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G141gat), .B(G148gat), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n434), .B1(KEYINPUT2), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT79), .ZN(new_n437));
  INV_X1    g236(.A(G148gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(G141gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(G141gat), .ZN(new_n440));
  INV_X1    g239(.A(G141gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G162gat), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT2), .B1(new_n444), .B2(KEYINPUT80), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n433), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n436), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n271), .A2(new_n279), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(new_n436), .A3(new_n446), .A4(new_n358), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT4), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n436), .A2(new_n446), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n285), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT84), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n447), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT3), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n436), .A2(new_n446), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n361), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n454), .A2(new_n458), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n468));
  INV_X1    g267(.A(new_n463), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n361), .A2(new_n447), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n451), .A2(new_n358), .B1(new_n436), .B2(new_n446), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT81), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n361), .A2(new_n447), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n452), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT81), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n469), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n466), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n463), .B(new_n462), .C1(new_n448), .C2(new_n457), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n468), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n476), .B1(new_n475), .B2(new_n469), .ZN(new_n481));
  AOI211_X1 g280(.A(KEYINPUT81), .B(new_n463), .C1(new_n474), .C2(new_n452), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n479), .B(new_n465), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n467), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT0), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G57gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(new_n219), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n485), .A2(KEYINPUT6), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT89), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n485), .A2(new_n493), .A3(KEYINPUT6), .A4(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n485), .A2(new_n490), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497));
  INV_X1    g296(.A(new_n467), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n478), .A2(new_n468), .A3(new_n479), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n489), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT38), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n418), .A2(new_n415), .A3(new_n419), .ZN(new_n505));
  OAI211_X1 g304(.A(KEYINPUT37), .B(new_n505), .C1(new_n407), .C2(new_n415), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n429), .A2(new_n504), .A3(new_n396), .A4(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n432), .A2(new_n495), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n415), .A2(new_n400), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n460), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n447), .ZN(new_n511));
  AND2_X1   g310(.A1(G228gat), .A2(G233gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n461), .A2(new_n400), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT85), .Z(new_n514));
  OAI211_X1 g313(.A(new_n511), .B(new_n512), .C1(new_n514), .C2(new_n415), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n510), .A2(new_n447), .B1(new_n414), .B2(new_n513), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT86), .B(G22gat), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT87), .A3(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G78gat), .B(G106gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT31), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n523), .B(G50gat), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n517), .A2(new_n526), .A3(new_n518), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n521), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n517), .A2(G22gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n519), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT30), .B1(new_n422), .B2(KEYINPUT78), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n428), .B1(new_n415), .B2(new_n407), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n396), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT78), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n535), .B(new_n536), .C1(new_n533), .C2(new_n396), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n454), .A2(new_n462), .A3(new_n458), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n469), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n475), .A2(new_n469), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT39), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT88), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OR3_X1    g342(.A1(new_n541), .A2(KEYINPUT88), .A3(new_n542), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n540), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n489), .B1(new_n540), .B2(KEYINPUT39), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT40), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n538), .A2(new_n549), .A3(new_n496), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n508), .A2(new_n531), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n531), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n503), .A2(new_n491), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(new_n538), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n391), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n385), .A2(new_n388), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n501), .A2(new_n489), .ZN(new_n557));
  AOI211_X1 g356(.A(new_n490), .B(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n492), .A2(new_n494), .B1(new_n559), .B2(new_n497), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n560), .A2(KEYINPUT35), .A3(new_n538), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n531), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n553), .ZN(new_n563));
  INV_X1    g362(.A(new_n538), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n531), .A2(new_n383), .A3(new_n384), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT35), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n555), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT94), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT18), .ZN(new_n571));
  NOR2_X1   g370(.A1(G15gat), .A2(G22gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G1gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(G15gat), .A2(G22gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(KEYINPUT16), .ZN(new_n577));
  INV_X1    g376(.A(new_n575), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(new_n572), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n579), .A3(KEYINPUT91), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n581), .B(new_n577), .C1(new_n578), .C2(new_n572), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(G8gat), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(KEYINPUT92), .B(G8gat), .Z(new_n584));
  NAND3_X1  g383(.A1(new_n576), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(G29gat), .A2(G36gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT14), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G29gat), .A2(G36gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G43gat), .B(G50gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT15), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G43gat), .B(G50gat), .Z(new_n596));
  INV_X1    g395(.A(KEYINPUT15), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT90), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n590), .B(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n598), .A2(new_n589), .A3(new_n593), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n586), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT13), .Z(new_n605));
  AOI21_X1  g404(.A(new_n571), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n570), .A2(KEYINPUT18), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n586), .A2(new_n602), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT93), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n583), .A2(new_n610), .A3(new_n585), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n583), .B2(new_n585), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n595), .A2(new_n601), .A3(KEYINPUT17), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT17), .B1(new_n595), .B2(new_n601), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n609), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n607), .B1(new_n618), .B2(new_n604), .ZN(new_n619));
  INV_X1    g418(.A(new_n613), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n595), .A2(new_n601), .A3(KEYINPUT17), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n620), .A2(new_n622), .A3(new_n623), .A4(new_n611), .ZN(new_n624));
  AND4_X1   g423(.A1(new_n608), .A2(new_n624), .A3(new_n604), .A4(new_n607), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n606), .B1(new_n619), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G197gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT11), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n299), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n629), .B(G169gat), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT12), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n626), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n635), .B(new_n606), .C1(new_n619), .C2(new_n625), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n248), .A2(new_n249), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n602), .ZN(new_n643));
  NAND3_X1  g442(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(KEYINPUT102), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n595), .A2(new_n601), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n248), .B2(new_n249), .ZN(new_n648));
  INV_X1    g447(.A(new_n644), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G190gat), .B(G218gat), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n622), .A2(new_n623), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n642), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n617), .A2(KEYINPUT101), .A3(new_n249), .A4(new_n248), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n651), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n652), .B1(new_n651), .B2(new_n657), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n641), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT102), .B1(new_n643), .B2(new_n644), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n648), .A2(new_n646), .A3(new_n649), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n652), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n651), .A2(new_n652), .A3(new_n657), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(KEYINPUT103), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G162gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT97), .B(G134gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n660), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n671), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n665), .A2(KEYINPUT103), .A3(new_n666), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(G127gat), .B(G155gat), .Z(new_n676));
  INV_X1    g475(.A(KEYINPUT21), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n583), .B(new_n585), .C1(new_n217), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n218), .A2(KEYINPUT21), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n680), .B2(new_n682), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n676), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  INV_X1    g486(.A(new_n676), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n683), .ZN(new_n689));
  XOR2_X1   g488(.A(G183gat), .B(G211gat), .Z(new_n690));
  NAND2_X1  g489(.A1(G231gat), .A2(G233gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n692), .B(new_n693), .Z(new_n694));
  AND3_X1   g493(.A1(new_n686), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n686), .B2(new_n689), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n640), .B1(new_n675), .B2(new_n698), .ZN(new_n699));
  AOI211_X1 g498(.A(KEYINPUT104), .B(new_n697), .C1(new_n672), .C2(new_n674), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND4_X1   g500(.A1(new_n263), .A2(new_n569), .A3(new_n639), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n553), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g503(.A1(new_n551), .A2(new_n554), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n705), .A2(new_n391), .B1(new_n562), .B2(new_n567), .ZN(new_n706));
  INV_X1    g505(.A(new_n639), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n263), .A3(new_n701), .ZN(new_n709));
  OAI21_X1  g508(.A(G8gat), .B1(new_n709), .B2(new_n564), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n711));
  OR2_X1    g510(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n702), .A2(new_n538), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n714), .A2(KEYINPUT106), .A3(new_n711), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT106), .B1(new_n714), .B2(new_n711), .ZN(new_n716));
  OAI221_X1 g515(.A(new_n710), .B1(new_n711), .B2(new_n714), .C1(new_n715), .C2(new_n716), .ZN(G1325gat));
  AOI21_X1  g516(.A(G15gat), .B1(new_n702), .B2(new_n556), .ZN(new_n718));
  INV_X1    g517(.A(G15gat), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n709), .A2(new_n719), .A3(new_n391), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(G1326gat));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n709), .B2(new_n531), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n702), .A2(new_n723), .A3(new_n552), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT43), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n722), .A2(new_n727), .A3(new_n724), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n726), .A2(G22gat), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(G22gat), .B1(new_n726), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(G1327gat));
  AND2_X1   g530(.A1(new_n672), .A2(new_n674), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n698), .A2(new_n262), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n708), .A2(new_n553), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n739), .A2(KEYINPUT45), .A3(G29gat), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT45), .B1(new_n739), .B2(G29gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n675), .B1(new_n555), .B2(new_n568), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n706), .A2(KEYINPUT44), .A3(new_n675), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n639), .B(new_n733), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G29gat), .B1(new_n747), .B2(new_n563), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n742), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1328gat));
  OAI21_X1  g552(.A(G36gat), .B1(new_n747), .B2(new_n564), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n708), .A2(new_n736), .A3(new_n738), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(G36gat), .A3(new_n564), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n755), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n758), .A2(KEYINPUT110), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(KEYINPUT110), .ZN(new_n760));
  OAI221_X1 g559(.A(new_n754), .B1(new_n755), .B2(new_n757), .C1(new_n759), .C2(new_n760), .ZN(G1329gat));
  INV_X1    g560(.A(G43gat), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n708), .A2(new_n762), .A3(new_n736), .A4(new_n738), .ZN(new_n763));
  INV_X1    g562(.A(new_n556), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n763), .A2(KEYINPUT111), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT111), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G43gat), .B1(new_n747), .B2(new_n391), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(KEYINPUT47), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1330gat));
  OAI21_X1  g572(.A(G50gat), .B1(new_n747), .B2(new_n531), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n756), .A2(G50gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n531), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT48), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1331gat));
  NOR2_X1   g577(.A1(new_n706), .A2(new_n263), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n699), .A2(new_n700), .A3(new_n639), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n553), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n538), .B1(new_n785), .B2(new_n394), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT112), .Z(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n394), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1333gat));
  OAI21_X1  g589(.A(G71gat), .B1(new_n781), .B2(new_n391), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n556), .A2(new_n208), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n781), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g593(.A1(new_n781), .A2(new_n531), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(new_n209), .ZN(G1335gat));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(KEYINPUT113), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n698), .A2(new_n639), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(KEYINPUT113), .B2(new_n797), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n799), .B1(new_n743), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n802), .ZN(new_n804));
  NOR4_X1   g603(.A1(new_n706), .A2(new_n675), .A3(new_n798), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n806), .A2(new_n219), .A3(new_n553), .A4(new_n262), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n801), .A2(new_n263), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n745), .B2(new_n746), .ZN(new_n809));
  OAI21_X1  g608(.A(G85gat), .B1(new_n809), .B2(new_n563), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(G1336gat));
  OAI211_X1 g610(.A(new_n538), .B(new_n808), .C1(new_n745), .C2(new_n746), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G92gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n551), .A2(new_n554), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n390), .B2(new_n389), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n552), .B1(new_n385), .B2(new_n388), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n553), .A2(new_n538), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n817), .A2(new_n384), .A3(new_n383), .A4(new_n531), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n816), .A2(new_n561), .B1(new_n818), .B2(KEYINPUT35), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n732), .B(new_n802), .C1(new_n815), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n798), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n743), .A2(new_n799), .A3(new_n802), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n564), .A2(G92gat), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n821), .A2(new_n262), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n813), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  INV_X1    g625(.A(new_n824), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n827), .A2(KEYINPUT114), .B1(G92gat), .B2(new_n812), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT115), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n806), .A2(KEYINPUT114), .A3(new_n262), .A4(new_n823), .ZN(new_n832));
  AND4_X1   g631(.A1(KEYINPUT115), .A2(new_n830), .A3(new_n813), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n826), .B1(new_n831), .B2(new_n833), .ZN(G1337gat));
  XNOR2_X1  g633(.A(KEYINPUT116), .B(G99gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n809), .B2(new_n391), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n764), .A2(new_n835), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n806), .A2(new_n262), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1338gat));
  NOR2_X1   g638(.A1(new_n809), .A2(new_n531), .ZN(new_n840));
  INV_X1    g639(.A(G106gat), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n531), .A2(G106gat), .A3(new_n263), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT117), .Z(new_n844));
  NOR3_X1   g643(.A1(new_n803), .A2(new_n805), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT53), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT53), .B1(new_n806), .B2(new_n843), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n840), .B2(new_n841), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1339gat));
  OAI22_X1  g648(.A1(new_n618), .A2(new_n604), .B1(new_n603), .B2(new_n605), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n630), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n638), .A2(new_n851), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n245), .A2(new_n250), .A3(new_n205), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(KEYINPUT54), .A3(new_n251), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n855), .B(new_n205), .C1(new_n245), .C2(new_n250), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n856), .A2(new_n857), .A3(new_n259), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n856), .B2(new_n259), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT55), .B(new_n854), .C1(new_n858), .C2(new_n859), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n852), .A2(new_n862), .A3(new_n260), .A4(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n732), .A2(new_n865), .A3(KEYINPUT119), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n862), .A2(new_n639), .A3(new_n260), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n262), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n675), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n675), .B2(new_n864), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n866), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n697), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n701), .A2(new_n263), .A3(new_n707), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n553), .A3(new_n564), .ZN(new_n877));
  INV_X1    g676(.A(new_n816), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G113gat), .B1(new_n880), .B2(new_n707), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n877), .A2(new_n566), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n272), .A3(new_n639), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1340gat));
  OAI21_X1  g683(.A(G120gat), .B1(new_n880), .B2(new_n263), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n357), .A3(new_n262), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1341gat));
  AOI21_X1  g686(.A(G127gat), .B1(new_n882), .B2(new_n698), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n698), .A2(G127gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n879), .B2(new_n889), .ZN(G1342gat));
  NOR4_X1   g689(.A1(new_n877), .A2(G134gat), .A3(new_n566), .A4(new_n675), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT56), .ZN(new_n892));
  OAI21_X1  g691(.A(G134gat), .B1(new_n880), .B2(new_n675), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1343gat));
  NOR2_X1   g693(.A1(new_n707), .A2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(new_n391), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n563), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n780), .A2(new_n263), .B1(new_n873), .B2(new_n697), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n531), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n897), .A2(new_n899), .A3(KEYINPUT121), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT121), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n564), .B(new_n895), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(new_n898), .B2(new_n531), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n876), .A2(KEYINPUT57), .A3(new_n552), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n391), .A2(new_n553), .A3(new_n564), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n639), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n902), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND4_X1   g711(.A1(new_n564), .A2(new_n897), .A3(new_n899), .A4(new_n895), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT120), .B1(new_n906), .B2(new_n908), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  AOI211_X1 g714(.A(new_n915), .B(new_n907), .C1(new_n904), .C2(new_n905), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n639), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n913), .B1(new_n917), .B2(G141gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n912), .B1(new_n918), .B2(new_n911), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT122), .B(new_n912), .C1(new_n918), .C2(new_n911), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1344gat));
  NOR2_X1   g722(.A1(new_n900), .A2(new_n901), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n538), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n438), .A3(new_n262), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n870), .B1(new_n675), .B2(new_n864), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT123), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n875), .B1(new_n929), .B2(new_n698), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT57), .B1(new_n930), .B2(new_n552), .ZN(new_n931));
  INV_X1    g730(.A(new_n905), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n262), .B(new_n908), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G148gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n927), .B1(new_n934), .B2(KEYINPUT59), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n936));
  AOI211_X1 g735(.A(KEYINPUT124), .B(new_n936), .C1(new_n933), .C2(G148gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n914), .A2(new_n916), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n939), .B2(new_n263), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(new_n438), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n926), .B1(new_n938), .B2(new_n941), .ZN(G1345gat));
  AOI21_X1  g741(.A(G155gat), .B1(new_n925), .B2(new_n698), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n939), .A2(new_n697), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(G155gat), .ZN(G1346gat));
  XNOR2_X1  g744(.A(KEYINPUT80), .B(G162gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n925), .A2(new_n732), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n939), .A2(new_n675), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n946), .ZN(G1347gat));
  NOR2_X1   g748(.A1(new_n564), .A2(new_n553), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n898), .A2(new_n878), .A3(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n707), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n898), .A2(new_n566), .A3(new_n951), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n955), .B(new_n639), .C1(new_n336), .C2(new_n335), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1348gat));
  AOI21_X1  g756(.A(G176gat), .B1(new_n955), .B2(new_n262), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n263), .A2(new_n256), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n952), .B2(new_n959), .ZN(G1349gat));
  OAI211_X1 g759(.A(new_n955), .B(new_n698), .C1(new_n288), .C2(new_n287), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT125), .Z(new_n962));
  OAI21_X1  g761(.A(G183gat), .B1(new_n953), .B2(new_n697), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g764(.A(new_n286), .B1(new_n952), .B2(new_n732), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT61), .Z(new_n967));
  NAND3_X1  g766(.A1(new_n955), .A2(new_n286), .A3(new_n732), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1351gat));
  INV_X1    g769(.A(G197gat), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n931), .A2(new_n932), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n896), .A2(new_n951), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n971), .B1(new_n974), .B2(new_n639), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n973), .A2(new_n899), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(new_n971), .A3(new_n639), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n975), .A2(new_n977), .ZN(G1352gat));
  NAND3_X1  g777(.A1(new_n976), .A2(new_n258), .A3(new_n262), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n979), .B(KEYINPUT62), .Z(new_n980));
  NAND3_X1  g779(.A1(new_n972), .A2(new_n262), .A3(new_n973), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n980), .B1(new_n982), .B2(new_n258), .ZN(G1353gat));
  NAND3_X1  g782(.A1(new_n976), .A2(new_n409), .A3(new_n698), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n698), .B(new_n973), .C1(new_n931), .C2(new_n932), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g789(.A(KEYINPUT127), .B(new_n984), .C1(new_n986), .C2(new_n987), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1354gat));
  AOI21_X1  g791(.A(G218gat), .B1(new_n976), .B2(new_n732), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n675), .A2(new_n410), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n993), .B1(new_n974), .B2(new_n994), .ZN(G1355gat));
endmodule


