//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n587, new_n588,
    new_n589, new_n590, new_n592, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n204), .B1(KEYINPUT87), .B2(new_n205), .C1(G1gat), .C2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT87), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209));
  INV_X1    g008(.A(G71gat), .ZN(new_n210));
  INV_X1    g009(.A(G78gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G57gat), .B(G64gat), .Z(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n213), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G71gat), .B(G78gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n208), .B1(KEYINPUT21), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(G183gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n219), .A2(KEYINPUT21), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G231gat), .A2(G233gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G155gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(G211gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n225), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232));
  INV_X1    g031(.A(G85gat), .ZN(new_n233));
  INV_X1    g032(.A(G92gat), .ZN(new_n234));
  AOI22_X1  g033(.A1(KEYINPUT8), .A2(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT93), .ZN(new_n236));
  NAND2_X1  g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT7), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G99gat), .B(G106gat), .Z(new_n240));
  XOR2_X1   g039(.A(new_n239), .B(new_n240), .Z(new_n241));
  INV_X1    g040(.A(KEYINPUT94), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n239), .A2(KEYINPUT94), .A3(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n246), .A2(KEYINPUT15), .ZN(new_n247));
  INV_X1    g046(.A(G29gat), .ZN(new_n248));
  INV_X1    g047(.A(G36gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT14), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT14), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(G29gat), .B2(G36gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n247), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(KEYINPUT86), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n246), .A2(KEYINPUT15), .ZN(new_n257));
  OR3_X1    g056(.A1(new_n256), .A2(new_n250), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n258), .B2(new_n247), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n245), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(KEYINPUT17), .Z(new_n261));
  OAI211_X1 g060(.A(new_n231), .B(new_n260), .C1(new_n261), .C2(new_n245), .ZN(new_n262));
  XNOR2_X1  g061(.A(G190gat), .B(G218gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n264), .B(KEYINPUT95), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n263), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G134gat), .B(G162gat), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n270), .B(KEYINPUT92), .Z(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n266), .B(KEYINPUT96), .Z(new_n273));
  NAND3_X1  g072(.A1(new_n265), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n230), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT97), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(KEYINPUT23), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n281), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n286), .A2(new_n287), .B1(KEYINPUT23), .B2(new_n279), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n283), .A2(KEYINPUT66), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT66), .B1(new_n283), .B2(new_n288), .ZN(new_n290));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT24), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n291), .A2(KEYINPUT24), .ZN(new_n293));
  OR2_X1    g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n289), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT67), .B1(new_n297), .B2(KEYINPUT25), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n288), .B(KEYINPUT68), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n283), .A4(new_n295), .ZN(new_n300));
  INV_X1    g099(.A(new_n290), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n288), .A3(KEYINPUT66), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n295), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT67), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n298), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n286), .A2(new_n287), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT26), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n279), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n291), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n313), .B(KEYINPUT70), .Z(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT27), .B(G183gat), .ZN(new_n315));
  INV_X1    g114(.A(G190gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(KEYINPUT28), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(KEYINPUT28), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n307), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n325), .B(KEYINPUT75), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n322), .A2(new_n326), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G197gat), .B(G204gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT74), .B(G218gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(KEYINPUT22), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G211gat), .ZN(new_n335));
  INV_X1    g134(.A(G211gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n332), .A2(KEYINPUT22), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(G218gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n327), .B1(new_n307), .B2(new_n321), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT76), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n328), .A2(new_n331), .A3(new_n339), .A4(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n339), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n326), .B1(new_n322), .B2(new_n323), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(KEYINPUT77), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n342), .A2(new_n345), .A3(new_n349), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n349), .B1(new_n342), .B2(new_n345), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT30), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(KEYINPUT35), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n363));
  XNOR2_X1  g162(.A(G127gat), .B(G134gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G113gat), .B(G120gat), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n365), .B1(KEYINPUT1), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n366), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT1), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n364), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n322), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n307), .A2(new_n371), .A3(new_n321), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G227gat), .ZN(new_n376));
  INV_X1    g175(.A(G233gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n363), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n307), .A2(new_n371), .A3(new_n321), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n371), .B1(new_n307), .B2(new_n321), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n363), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n362), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G15gat), .B(G43gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(G71gat), .B(G99gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n361), .B1(new_n387), .B2(new_n360), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n389), .B1(new_n379), .B2(new_n383), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT73), .B(new_n389), .C1(new_n379), .C2(new_n383), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT34), .ZN(new_n395));
  INV_X1    g194(.A(new_n375), .ZN(new_n396));
  INV_X1    g195(.A(new_n378), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n375), .A2(KEYINPUT34), .A3(new_n378), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n394), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(KEYINPUT83), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n409));
  XNOR2_X1  g208(.A(G141gat), .B(G148gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(KEYINPUT2), .ZN(new_n411));
  XNOR2_X1  g210(.A(G155gat), .B(G162gat), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT78), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n412), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT78), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n414), .B(new_n415), .C1(KEYINPUT2), .C2(new_n410), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OR2_X1    g216(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(G162gat), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n410), .B1(new_n420), .B2(KEYINPUT2), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n412), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n409), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n417), .A2(new_n408), .A3(new_n422), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n323), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n339), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G22gat), .ZN(new_n429));
  INV_X1    g228(.A(G22gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n424), .A2(new_n430), .A3(new_n427), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(G228gat), .A3(G233gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n405), .A2(KEYINPUT83), .ZN(new_n434));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n435), .A3(new_n431), .ZN(new_n436));
  AND4_X1   g235(.A1(new_n407), .A2(new_n433), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n407), .B1(new_n433), .B2(new_n436), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n388), .A2(new_n392), .A3(new_n400), .A4(new_n393), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n402), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n423), .A2(new_n372), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n417), .A2(new_n371), .A3(new_n422), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT5), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT81), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n442), .ZN(new_n448));
  INV_X1    g247(.A(new_n444), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n371), .B1(new_n417), .B2(new_n422), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT81), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n423), .A2(KEYINPUT3), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n372), .A3(new_n425), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n449), .A2(KEYINPUT4), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n458));
  NAND2_X1  g257(.A1(new_n444), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n456), .A2(new_n457), .A3(new_n442), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n456), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n444), .A2(new_n463), .A3(KEYINPUT4), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n444), .B2(KEYINPUT4), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n458), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n448), .A2(KEYINPUT5), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G1gat), .B(G29gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G85gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT0), .B(G57gat), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n473), .B(new_n474), .Z(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT84), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478));
  AOI211_X1 g277(.A(new_n478), .B(new_n475), .C1(new_n461), .C2(new_n470), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n471), .B2(new_n476), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n460), .A2(new_n454), .B1(new_n468), .B2(new_n469), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n484), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT6), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n359), .A2(new_n441), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n486), .B1(new_n485), .B2(new_n482), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n353), .A2(new_n492), .A3(new_n357), .A4(new_n354), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n491), .B(KEYINPUT35), .C1(new_n441), .C2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AND4_X1   g294(.A1(new_n492), .A2(new_n353), .A3(new_n354), .A4(new_n357), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n496), .A2(new_n439), .A3(new_n440), .A4(new_n402), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n491), .B1(new_n497), .B2(KEYINPUT35), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n490), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n437), .A2(new_n438), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n394), .A2(new_n401), .ZN(new_n504));
  INV_X1    g303(.A(new_n440), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n402), .A2(KEYINPUT36), .A3(new_n440), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n342), .A2(new_n509), .A3(new_n345), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n342), .B2(new_n345), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n349), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n355), .B1(new_n513), .B2(KEYINPUT38), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n328), .A2(new_n331), .A3(new_n343), .A4(new_n341), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n339), .B1(new_n344), .B2(new_n340), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(KEYINPUT37), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT38), .B1(new_n517), .B2(new_n510), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n349), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n488), .A3(new_n519), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n468), .A2(KEYINPUT39), .A3(new_n442), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n468), .A2(new_n442), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n449), .A2(new_n450), .A3(new_n448), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI211_X1 g323(.A(new_n476), .B(new_n521), .C1(new_n524), .C2(KEYINPUT39), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n480), .B1(KEYINPUT40), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n358), .B(new_n526), .C1(KEYINPUT40), .C2(new_n525), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n520), .A2(new_n527), .A3(new_n439), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n508), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n499), .B1(new_n502), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n277), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G113gat), .B(G141gat), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G197gat), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT11), .B(G169gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT12), .Z(new_n536));
  NOR2_X1   g335(.A1(new_n261), .A2(new_n208), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n259), .A2(new_n208), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT88), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT18), .ZN(new_n543));
  INV_X1    g342(.A(new_n539), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n259), .B2(new_n208), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n541), .B(KEYINPUT13), .Z(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n536), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n548), .A2(KEYINPUT89), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(KEYINPUT89), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n543), .A2(new_n536), .A3(new_n547), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n552), .A2(KEYINPUT90), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(KEYINPUT90), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n245), .A2(KEYINPUT10), .A3(new_n219), .ZN(new_n558));
  INV_X1    g357(.A(new_n219), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n241), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n245), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n558), .B1(new_n561), .B2(KEYINPUT10), .ZN(new_n562));
  INV_X1    g361(.A(G230gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(new_n377), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n564), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  OR3_X1    g371(.A1(new_n567), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n567), .B2(new_n569), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n557), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n531), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(new_n492), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT98), .B(G1gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(G1324gat));
  INV_X1    g379(.A(new_n358), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n583), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT42), .Z(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n205), .B2(new_n582), .ZN(G1325gat));
  INV_X1    g385(.A(G15gat), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n577), .A2(new_n587), .A3(new_n508), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n504), .A2(new_n505), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n531), .A2(new_n576), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n587), .B2(new_n590), .ZN(G1326gat));
  NOR2_X1   g390(.A1(new_n577), .A2(new_n439), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n430), .ZN(new_n593));
  XOR2_X1   g392(.A(KEYINPUT99), .B(KEYINPUT43), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(G1327gat));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n501), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT101), .B1(new_n493), .B2(new_n500), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n596), .B1(new_n529), .B2(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n598), .A2(new_n599), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n602), .A2(KEYINPUT102), .A3(new_n508), .A4(new_n528), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT103), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT35), .B1(new_n441), .B2(new_n493), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT85), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n494), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n605), .B1(new_n608), .B2(new_n490), .ZN(new_n609));
  AOI211_X1 g408(.A(KEYINPUT103), .B(new_n489), .C1(new_n607), .C2(new_n494), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT44), .B1(new_n611), .B2(new_n275), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n530), .A2(new_n275), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(KEYINPUT44), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n575), .B(KEYINPUT100), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n614), .A2(new_n556), .A3(new_n230), .A4(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(G29gat), .B1(new_n616), .B2(new_n492), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n613), .A2(new_n576), .A3(new_n230), .ZN(new_n618));
  INV_X1    g417(.A(new_n492), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n248), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT45), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(G1328gat));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n249), .A3(new_n358), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT46), .Z(new_n624));
  OAI21_X1  g423(.A(G36gat), .B1(new_n616), .B2(new_n581), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(G1329gat));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627));
  INV_X1    g426(.A(G43gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n618), .A2(new_n628), .A3(new_n589), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT105), .Z(new_n630));
  OAI21_X1  g429(.A(G43gat), .B1(new_n616), .B2(new_n508), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g432(.A(KEYINPUT48), .ZN(new_n634));
  OAI21_X1  g433(.A(G50gat), .B1(new_n616), .B2(new_n439), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT106), .ZN(new_n636));
  INV_X1    g435(.A(G50gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n618), .A2(new_n637), .A3(new_n500), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n634), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n634), .B1(new_n638), .B2(KEYINPUT107), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n635), .B(new_n641), .C1(KEYINPUT107), .C2(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(G1331gat));
  AND3_X1   g442(.A1(new_n611), .A2(new_n557), .A3(new_n277), .ZN(new_n644));
  INV_X1    g443(.A(new_n615), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n492), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT108), .B(G57gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1332gat));
  INV_X1    g448(.A(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n581), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT109), .ZN(new_n654));
  NOR2_X1   g453(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1333gat));
  INV_X1    g455(.A(new_n589), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n210), .B1(new_n646), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n508), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(G71gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n646), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1334gat));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n439), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(new_n211), .ZN(G1335gat));
  INV_X1    g464(.A(new_n230), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n556), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n614), .A2(new_n575), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n492), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT111), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n499), .A2(KEYINPUT103), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n608), .A2(new_n605), .A3(new_n490), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n671), .A2(new_n672), .B1(new_n601), .B2(new_n603), .ZN(new_n673));
  INV_X1    g472(.A(new_n275), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT112), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT112), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n611), .A2(new_n676), .A3(new_n275), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n667), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT51), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n675), .A2(new_n677), .A3(KEYINPUT51), .A4(new_n667), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n575), .A2(new_n233), .A3(new_n619), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT113), .ZN(new_n685));
  OAI22_X1  g484(.A1(new_n670), .A2(new_n233), .B1(new_n683), .B2(new_n685), .ZN(G1336gat));
  NOR2_X1   g485(.A1(new_n581), .A2(G92gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n682), .A2(new_n645), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G92gat), .B1(new_n668), .B2(new_n581), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT52), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT116), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT114), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n682), .A2(KEYINPUT114), .A3(new_n645), .A4(new_n687), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n689), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT115), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n697), .A2(new_n698), .A3(KEYINPUT52), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n697), .B2(KEYINPUT52), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n693), .B1(new_n699), .B2(new_n700), .ZN(G1337gat));
  OAI21_X1  g500(.A(G99gat), .B1(new_n668), .B2(new_n508), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n683), .A2(G99gat), .A3(new_n657), .ZN(new_n703));
  INV_X1    g502(.A(new_n575), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(G1338gat));
  INV_X1    g504(.A(G106gat), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n682), .A2(new_n706), .A3(new_n500), .A4(new_n645), .ZN(new_n707));
  OAI21_X1  g506(.A(G106gat), .B1(new_n668), .B2(new_n439), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g509(.A1(new_n540), .A2(new_n541), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n545), .A2(new_n546), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n535), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n553), .B2(new_n554), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n575), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n562), .A2(new_n565), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(KEYINPUT54), .A3(new_n566), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n718), .B(new_n572), .C1(KEYINPUT54), .C2(new_n566), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT55), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n573), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n716), .B1(new_n557), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n674), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n715), .A2(new_n573), .A3(new_n275), .A4(new_n720), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n666), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n277), .A2(new_n704), .A3(new_n557), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n581), .A2(new_n619), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n728), .A2(new_n441), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n556), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G113gat), .ZN(G1340gat));
  AOI21_X1  g531(.A(G120gat), .B1(new_n730), .B2(new_n575), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n645), .A2(G120gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n730), .B2(new_n734), .ZN(G1341gat));
  INV_X1    g534(.A(KEYINPUT118), .ZN(new_n736));
  INV_X1    g535(.A(G127gat), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT117), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(KEYINPUT117), .B2(new_n737), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n730), .A2(new_n666), .ZN(new_n740));
  MUX2_X1   g539(.A(new_n739), .B(new_n738), .S(new_n740), .Z(G1342gat));
  NAND2_X1  g540(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n730), .A2(new_n275), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n743), .B(new_n744), .Z(G1343gat));
  NOR2_X1   g544(.A1(new_n728), .A2(new_n729), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n659), .A2(new_n439), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n747), .A2(KEYINPUT122), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(KEYINPUT122), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(G141gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n752), .A3(new_n556), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT57), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n721), .A2(KEYINPUT120), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n721), .A2(KEYINPUT120), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n556), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT119), .B1(new_n715), .B2(new_n575), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n715), .A2(KEYINPUT119), .A3(new_n575), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(new_n674), .ZN(new_n762));
  INV_X1    g561(.A(new_n724), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT121), .B(new_n230), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT121), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n763), .B1(new_n761), .B2(new_n674), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n666), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n767), .A3(new_n726), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n754), .B1(new_n768), .B2(new_n500), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n728), .A2(KEYINPUT57), .A3(new_n439), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n659), .A2(new_n729), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NOR4_X1   g571(.A1(new_n769), .A2(new_n770), .A3(new_n557), .A4(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n753), .B1(new_n773), .B2(new_n752), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT58), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n776), .B(new_n753), .C1(new_n773), .C2(new_n752), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1344gat));
  INV_X1    g577(.A(G148gat), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n780));
  AOI211_X1 g579(.A(KEYINPUT59), .B(new_n779), .C1(new_n780), .C2(new_n575), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT59), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT57), .B1(new_n728), .B2(new_n439), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n726), .B1(new_n766), .B2(new_n666), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n754), .A3(new_n500), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n575), .A3(new_n771), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n782), .B1(new_n787), .B2(G148gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n575), .A2(new_n779), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n781), .A2(new_n788), .B1(new_n750), .B2(new_n789), .ZN(G1345gat));
  NAND2_X1  g589(.A1(new_n418), .A2(new_n419), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n751), .A2(new_n666), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n230), .A2(new_n791), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n791), .A2(new_n792), .B1(new_n780), .B2(new_n793), .ZN(G1346gat));
  OR2_X1    g593(.A1(new_n674), .A2(G162gat), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n750), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n768), .A2(new_n500), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT57), .ZN(new_n798));
  INV_X1    g597(.A(new_n770), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n798), .A2(new_n275), .A3(new_n799), .A4(new_n771), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n796), .B1(new_n800), .B2(G162gat), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT123), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT123), .B(new_n796), .C1(new_n800), .C2(G162gat), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(G1347gat));
  NOR2_X1   g604(.A1(new_n728), .A2(new_n619), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n441), .A2(new_n581), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(G169gat), .B1(new_n808), .B2(new_n557), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(KEYINPUT124), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n807), .A2(KEYINPUT124), .ZN(new_n811));
  NOR4_X1   g610(.A1(new_n728), .A2(new_n619), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(G169gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n556), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n814), .ZN(G1348gat));
  INV_X1    g614(.A(G176gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n808), .A2(new_n816), .A3(new_n615), .ZN(new_n817));
  AOI21_X1  g616(.A(G176gat), .B1(new_n812), .B2(new_n575), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(G1349gat));
  OAI21_X1  g618(.A(G183gat), .B1(new_n808), .B2(new_n230), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n812), .A2(new_n315), .A3(new_n666), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g622(.A(G190gat), .B1(new_n808), .B2(new_n674), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT61), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n812), .A2(new_n316), .A3(new_n275), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1351gat));
  NOR2_X1   g626(.A1(new_n659), .A2(new_n619), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n786), .A2(new_n358), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G197gat), .B1(new_n829), .B2(new_n557), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n747), .A2(new_n358), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT125), .Z(new_n832));
  NAND2_X1  g631(.A1(new_n806), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n557), .A2(G197gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(G1352gat));
  NOR3_X1   g634(.A1(new_n833), .A2(G204gat), .A3(new_n704), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT62), .ZN(new_n838));
  OAI21_X1  g637(.A(G204gat), .B1(new_n829), .B2(new_n615), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT126), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(new_n840), .A3(KEYINPUT62), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n837), .B2(KEYINPUT62), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n838), .B(new_n839), .C1(new_n842), .C2(new_n843), .ZN(G1353gat));
  NAND4_X1  g643(.A1(new_n806), .A2(new_n336), .A3(new_n666), .A4(new_n832), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n786), .A2(new_n358), .A3(new_n666), .A4(new_n828), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT63), .B1(new_n846), .B2(G211gat), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(G1354gat));
  INV_X1    g649(.A(G218gat), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n833), .B2(new_n674), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n275), .A2(new_n333), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n829), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


