

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U554 ( .A(KEYINPUT72), .B(n584), .Z(n521) );
  OR2_X1 U555 ( .A1(n771), .A2(n770), .ZN(n522) );
  AND2_X1 U556 ( .A1(n737), .A2(n736), .ZN(n523) );
  NOR2_X1 U557 ( .A1(n708), .A2(n709), .ZN(n703) );
  INV_X1 U558 ( .A(G168), .ZN(n736) );
  INV_X1 U559 ( .A(KEYINPUT100), .ZN(n731) );
  NOR2_X1 U560 ( .A1(n745), .A2(n744), .ZN(n746) );
  INV_X1 U561 ( .A(n959), .ZN(n770) );
  NAND2_X1 U562 ( .A1(G8), .A2(n752), .ZN(n779) );
  NOR2_X1 U563 ( .A1(G1384), .A2(G164), .ZN(n695) );
  XNOR2_X1 U564 ( .A(KEYINPUT15), .B(n588), .ZN(n979) );
  NOR2_X1 U565 ( .A1(n634), .A2(G651), .ZN(n664) );
  NOR2_X1 U566 ( .A1(n551), .A2(n550), .ZN(G160) );
  NOR2_X2 U567 ( .A1(G543), .A2(G651), .ZN(n655) );
  NAND2_X1 U568 ( .A1(n655), .A2(G89), .ZN(n524) );
  XNOR2_X1 U569 ( .A(n524), .B(KEYINPUT4), .ZN(n526) );
  XOR2_X1 U570 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  INV_X1 U571 ( .A(G651), .ZN(n528) );
  NOR2_X2 U572 ( .A1(n634), .A2(n528), .ZN(n659) );
  NAND2_X1 U573 ( .A1(G76), .A2(n659), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U575 ( .A(n527), .B(KEYINPUT5), .ZN(n534) );
  NOR2_X1 U576 ( .A1(G543), .A2(n528), .ZN(n529) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n529), .Z(n656) );
  NAND2_X1 U578 ( .A1(G63), .A2(n656), .ZN(n531) );
  NAND2_X1 U579 ( .A1(G51), .A2(n664), .ZN(n530) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U581 ( .A(KEYINPUT6), .B(n532), .Z(n533) );
  NAND2_X1 U582 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U583 ( .A(n535), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U584 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  OR2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  XNOR2_X2 U586 ( .A(KEYINPUT17), .B(n536), .ZN(n882) );
  AND2_X1 U587 ( .A1(G138), .A2(n882), .ZN(n544) );
  INV_X1 U588 ( .A(G2105), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n537), .A2(G2104), .ZN(n538) );
  XNOR2_X2 U590 ( .A(n538), .B(KEYINPUT65), .ZN(n883) );
  NAND2_X1 U591 ( .A1(G102), .A2(n883), .ZN(n542) );
  NOR2_X1 U592 ( .A1(G2104), .A2(n537), .ZN(n878) );
  NAND2_X1 U593 ( .A1(G126), .A2(n878), .ZN(n540) );
  AND2_X1 U594 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U595 ( .A1(G114), .A2(n879), .ZN(n539) );
  AND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U598 ( .A1(n544), .A2(n543), .ZN(G164) );
  NAND2_X1 U599 ( .A1(G125), .A2(n878), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G113), .A2(n879), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n551) );
  NAND2_X1 U602 ( .A1(G101), .A2(n883), .ZN(n547) );
  XOR2_X1 U603 ( .A(KEYINPUT23), .B(n547), .Z(n549) );
  NAND2_X1 U604 ( .A1(n882), .A2(G137), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U606 ( .A(G2446), .B(G2430), .Z(n553) );
  XNOR2_X1 U607 ( .A(G2451), .B(KEYINPUT108), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U609 ( .A(n554), .B(G2427), .Z(n556) );
  XNOR2_X1 U610 ( .A(G1341), .B(G1348), .ZN(n555) );
  XNOR2_X1 U611 ( .A(n556), .B(n555), .ZN(n560) );
  XOR2_X1 U612 ( .A(G2443), .B(G2435), .Z(n558) );
  XNOR2_X1 U613 ( .A(G2438), .B(G2454), .ZN(n557) );
  XNOR2_X1 U614 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U615 ( .A(n560), .B(n559), .Z(n561) );
  AND2_X1 U616 ( .A1(G14), .A2(n561), .ZN(G401) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G132), .ZN(G219) );
  INV_X1 U619 ( .A(G82), .ZN(G220) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  INV_X1 U621 ( .A(G120), .ZN(G236) );
  NAND2_X1 U622 ( .A1(G90), .A2(n655), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G77), .A2(n659), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U625 ( .A(KEYINPUT9), .B(n564), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G64), .A2(n656), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G52), .A2(n664), .ZN(n565) );
  AND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(G301) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n569) );
  XOR2_X1 U631 ( .A(n569), .B(KEYINPUT10), .Z(n836) );
  NAND2_X1 U632 ( .A1(n836), .A2(G567), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  INV_X1 U634 ( .A(G860), .ZN(n602) );
  NAND2_X1 U635 ( .A1(G56), .A2(n656), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n571), .Z(n578) );
  NAND2_X1 U637 ( .A1(G81), .A2(n655), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT12), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT70), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G68), .A2(n659), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U642 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n664), .A2(G43), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n974) );
  NOR2_X1 U646 ( .A1(n602), .A2(n974), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT71), .ZN(G153) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U649 ( .A1(n664), .A2(G54), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G92), .A2(n655), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G66), .A2(n656), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n659), .A2(G79), .ZN(n584) );
  NOR2_X1 U654 ( .A1(n585), .A2(n521), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  INV_X1 U656 ( .A(n979), .ZN(n708) );
  INV_X1 U657 ( .A(G868), .ZN(n599) );
  NAND2_X1 U658 ( .A1(n708), .A2(n599), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G91), .A2(n655), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G53), .A2(n664), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n598) );
  NAND2_X1 U663 ( .A1(G65), .A2(n656), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n593), .B(KEYINPUT68), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G78), .A2(n659), .ZN(n594) );
  XOR2_X1 U666 ( .A(KEYINPUT67), .B(n594), .Z(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n962) );
  XNOR2_X1 U669 ( .A(n962), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U670 ( .A1(G286), .A2(G868), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n599), .A2(G299), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U673 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n603), .A2(n979), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U676 ( .A1(n979), .A2(G868), .ZN(n605) );
  NOR2_X1 U677 ( .A1(G559), .A2(n605), .ZN(n606) );
  XOR2_X1 U678 ( .A(KEYINPUT74), .B(n606), .Z(n609) );
  NOR2_X1 U679 ( .A1(G868), .A2(n974), .ZN(n607) );
  XNOR2_X1 U680 ( .A(KEYINPUT73), .B(n607), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U682 ( .A(KEYINPUT75), .B(n610), .ZN(G282) );
  XOR2_X1 U683 ( .A(G2100), .B(KEYINPUT78), .Z(n621) );
  XOR2_X1 U684 ( .A(KEYINPUT18), .B(KEYINPUT77), .Z(n612) );
  NAND2_X1 U685 ( .A1(G123), .A2(n878), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n613), .B(KEYINPUT76), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n879), .A2(G111), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G135), .A2(n882), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G99), .A2(n883), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n1002) );
  XNOR2_X1 U694 ( .A(G2096), .B(n1002), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(G156) );
  NAND2_X1 U696 ( .A1(n664), .A2(G55), .ZN(n622) );
  XOR2_X1 U697 ( .A(KEYINPUT81), .B(n622), .Z(n624) );
  NAND2_X1 U698 ( .A1(n656), .A2(G67), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U700 ( .A(KEYINPUT82), .B(n625), .ZN(n630) );
  NAND2_X1 U701 ( .A1(G80), .A2(n659), .ZN(n626) );
  XNOR2_X1 U702 ( .A(n626), .B(KEYINPUT80), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n655), .A2(G93), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n677) );
  NAND2_X1 U706 ( .A1(n979), .A2(G559), .ZN(n675) );
  XOR2_X1 U707 ( .A(KEYINPUT79), .B(n974), .Z(n631) );
  XNOR2_X1 U708 ( .A(n675), .B(n631), .ZN(n632) );
  NOR2_X1 U709 ( .A1(G860), .A2(n632), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n677), .B(n633), .ZN(G145) );
  NAND2_X1 U711 ( .A1(G49), .A2(n664), .ZN(n636) );
  NAND2_X1 U712 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U714 ( .A1(n656), .A2(n637), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n638) );
  XOR2_X1 U716 ( .A(KEYINPUT83), .B(n638), .Z(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U718 ( .A(KEYINPUT84), .B(n641), .ZN(G288) );
  NAND2_X1 U719 ( .A1(G60), .A2(n656), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G47), .A2(n664), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U722 ( .A(KEYINPUT66), .B(n644), .Z(n648) );
  NAND2_X1 U723 ( .A1(G85), .A2(n655), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G72), .A2(n659), .ZN(n645) );
  AND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(G290) );
  NAND2_X1 U727 ( .A1(G88), .A2(n655), .ZN(n650) );
  NAND2_X1 U728 ( .A1(G75), .A2(n659), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U730 ( .A1(G62), .A2(n656), .ZN(n652) );
  NAND2_X1 U731 ( .A1(G50), .A2(n664), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U733 ( .A1(n654), .A2(n653), .ZN(G166) );
  INV_X1 U734 ( .A(G166), .ZN(G303) );
  NAND2_X1 U735 ( .A1(G86), .A2(n655), .ZN(n658) );
  NAND2_X1 U736 ( .A1(G61), .A2(n656), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n663) );
  NAND2_X1 U738 ( .A1(G73), .A2(n659), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n660), .B(KEYINPUT85), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n661), .B(KEYINPUT2), .ZN(n662) );
  NOR2_X1 U741 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n664), .A2(G48), .ZN(n665) );
  NAND2_X1 U743 ( .A1(n666), .A2(n665), .ZN(G305) );
  XOR2_X1 U744 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n667) );
  XNOR2_X1 U745 ( .A(G290), .B(n667), .ZN(n668) );
  XOR2_X1 U746 ( .A(n668), .B(KEYINPUT19), .Z(n670) );
  XOR2_X1 U747 ( .A(G303), .B(n677), .Z(n669) );
  XNOR2_X1 U748 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U749 ( .A(n671), .B(n974), .ZN(n672) );
  XNOR2_X1 U750 ( .A(n672), .B(G299), .ZN(n673) );
  XNOR2_X1 U751 ( .A(G288), .B(n673), .ZN(n674) );
  XNOR2_X1 U752 ( .A(n674), .B(G305), .ZN(n903) );
  XNOR2_X1 U753 ( .A(n675), .B(n903), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n676), .A2(G868), .ZN(n679) );
  OR2_X1 U755 ( .A1(G868), .A2(n677), .ZN(n678) );
  NAND2_X1 U756 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2084), .A2(G2078), .ZN(n681) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n680) );
  XNOR2_X1 U759 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U762 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U764 ( .A1(G236), .A2(G237), .ZN(n685) );
  NAND2_X1 U765 ( .A1(G69), .A2(n685), .ZN(n686) );
  XNOR2_X1 U766 ( .A(KEYINPUT89), .B(n686), .ZN(n687) );
  NAND2_X1 U767 ( .A1(n687), .A2(G108), .ZN(n841) );
  NAND2_X1 U768 ( .A1(G567), .A2(n841), .ZN(n692) );
  NOR2_X1 U769 ( .A1(G220), .A2(G219), .ZN(n688) );
  XOR2_X1 U770 ( .A(KEYINPUT22), .B(n688), .Z(n689) );
  NOR2_X1 U771 ( .A1(G218), .A2(n689), .ZN(n690) );
  NAND2_X1 U772 ( .A1(G96), .A2(n690), .ZN(n842) );
  NAND2_X1 U773 ( .A1(G2106), .A2(n842), .ZN(n691) );
  NAND2_X1 U774 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U775 ( .A(KEYINPUT90), .B(n693), .ZN(n840) );
  NAND2_X1 U776 ( .A1(G661), .A2(G483), .ZN(n694) );
  NOR2_X1 U777 ( .A1(n840), .A2(n694), .ZN(n839) );
  NAND2_X1 U778 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n802) );
  INV_X1 U780 ( .A(n802), .ZN(n696) );
  XNOR2_X1 U781 ( .A(n695), .B(KEYINPUT64), .ZN(n801) );
  AND2_X2 U782 ( .A1(n696), .A2(n801), .ZN(n726) );
  INV_X1 U783 ( .A(n726), .ZN(n752) );
  NOR2_X1 U784 ( .A1(G1966), .A2(n779), .ZN(n745) );
  INV_X1 U785 ( .A(KEYINPUT26), .ZN(n698) );
  AND2_X1 U786 ( .A1(G1996), .A2(n726), .ZN(n697) );
  XNOR2_X1 U787 ( .A(n698), .B(n697), .ZN(n702) );
  NAND2_X1 U788 ( .A1(G1341), .A2(n752), .ZN(n700) );
  INV_X1 U789 ( .A(n974), .ZN(n699) );
  AND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n709) );
  XNOR2_X1 U792 ( .A(n703), .B(KEYINPUT99), .ZN(n707) );
  NOR2_X1 U793 ( .A1(n726), .A2(G1348), .ZN(n705) );
  NOR2_X1 U794 ( .A1(G2067), .A2(n752), .ZN(n704) );
  NOR2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U797 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n718) );
  XOR2_X1 U799 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n713) );
  NAND2_X1 U800 ( .A1(G2072), .A2(n726), .ZN(n712) );
  XNOR2_X1 U801 ( .A(n713), .B(n712), .ZN(n716) );
  NAND2_X1 U802 ( .A1(G1956), .A2(n752), .ZN(n714) );
  XOR2_X1 U803 ( .A(KEYINPUT98), .B(n714), .Z(n715) );
  NOR2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n962), .A2(n719), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n723) );
  NOR2_X1 U807 ( .A1(n962), .A2(n719), .ZN(n721) );
  INV_X1 U808 ( .A(KEYINPUT28), .ZN(n720) );
  XNOR2_X1 U809 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U811 ( .A(n724), .B(KEYINPUT29), .ZN(n730) );
  XNOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .ZN(n915) );
  NAND2_X1 U813 ( .A1(n726), .A2(n915), .ZN(n725) );
  XOR2_X1 U814 ( .A(KEYINPUT96), .B(n725), .Z(n728) );
  NOR2_X1 U815 ( .A1(n726), .A2(G1961), .ZN(n727) );
  NOR2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n738) );
  NOR2_X1 U817 ( .A1(G301), .A2(n738), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n732) );
  XNOR2_X1 U819 ( .A(n732), .B(n731), .ZN(n743) );
  INV_X1 U820 ( .A(KEYINPUT31), .ZN(n741) );
  NOR2_X1 U821 ( .A1(G2084), .A2(n752), .ZN(n747) );
  NOR2_X1 U822 ( .A1(n745), .A2(n747), .ZN(n733) );
  NAND2_X1 U823 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U824 ( .A(KEYINPUT101), .B(n734), .ZN(n735) );
  XNOR2_X1 U825 ( .A(n735), .B(KEYINPUT30), .ZN(n737) );
  AND2_X1 U826 ( .A1(G301), .A2(n738), .ZN(n739) );
  NOR2_X1 U827 ( .A1(n523), .A2(n739), .ZN(n740) );
  XNOR2_X1 U828 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n751) );
  INV_X1 U830 ( .A(n751), .ZN(n744) );
  XNOR2_X1 U831 ( .A(n746), .B(KEYINPUT102), .ZN(n750) );
  NAND2_X1 U832 ( .A1(G8), .A2(n747), .ZN(n748) );
  XOR2_X1 U833 ( .A(KEYINPUT95), .B(n748), .Z(n749) );
  NAND2_X1 U834 ( .A1(n750), .A2(n749), .ZN(n762) );
  NAND2_X1 U835 ( .A1(n751), .A2(G286), .ZN(n757) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n779), .ZN(n754) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n752), .ZN(n753) );
  NOR2_X1 U838 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U839 ( .A1(n755), .A2(G303), .ZN(n756) );
  NAND2_X1 U840 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U841 ( .A1(n758), .A2(G8), .ZN(n760) );
  XOR2_X1 U842 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n759) );
  XNOR2_X1 U843 ( .A(n760), .B(n759), .ZN(n761) );
  NAND2_X1 U844 ( .A1(n762), .A2(n761), .ZN(n775) );
  NOR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n763) );
  XNOR2_X1 U847 ( .A(KEYINPUT104), .B(n763), .ZN(n764) );
  NOR2_X1 U848 ( .A1(n965), .A2(n764), .ZN(n765) );
  NAND2_X1 U849 ( .A1(n775), .A2(n765), .ZN(n766) );
  NAND2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n966) );
  NAND2_X1 U851 ( .A1(n766), .A2(n966), .ZN(n767) );
  NOR2_X1 U852 ( .A1(n779), .A2(n767), .ZN(n768) );
  NOR2_X1 U853 ( .A1(KEYINPUT33), .A2(n768), .ZN(n772) );
  NAND2_X1 U854 ( .A1(n965), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n769), .A2(n779), .ZN(n771) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n959) );
  NOR2_X1 U857 ( .A1(n772), .A2(n522), .ZN(n783) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U861 ( .A1(n776), .A2(n779), .ZN(n781) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U863 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  OR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U866 ( .A1(n783), .A2(n782), .ZN(n807) );
  NAND2_X1 U867 ( .A1(G129), .A2(n878), .ZN(n785) );
  NAND2_X1 U868 ( .A1(G117), .A2(n879), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U870 ( .A1(G105), .A2(n883), .ZN(n786) );
  XNOR2_X1 U871 ( .A(n786), .B(KEYINPUT93), .ZN(n787) );
  XNOR2_X1 U872 ( .A(n787), .B(KEYINPUT38), .ZN(n788) );
  NOR2_X1 U873 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U874 ( .A1(n882), .A2(G141), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n893) );
  NAND2_X1 U876 ( .A1(G1996), .A2(n893), .ZN(n800) );
  NAND2_X1 U877 ( .A1(G119), .A2(n878), .ZN(n793) );
  NAND2_X1 U878 ( .A1(G131), .A2(n882), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U880 ( .A1(n879), .A2(G107), .ZN(n794) );
  XOR2_X1 U881 ( .A(KEYINPUT92), .B(n794), .Z(n795) );
  NOR2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U883 ( .A1(n883), .A2(G95), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n889) );
  NAND2_X1 U885 ( .A1(G1991), .A2(n889), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n1005) );
  NOR2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n830) );
  NAND2_X1 U888 ( .A1(n1005), .A2(n830), .ZN(n803) );
  XOR2_X1 U889 ( .A(n803), .B(KEYINPUT94), .Z(n821) );
  INV_X1 U890 ( .A(n821), .ZN(n805) );
  XNOR2_X1 U891 ( .A(G1986), .B(G290), .ZN(n970) );
  NAND2_X1 U892 ( .A1(n830), .A2(n970), .ZN(n804) );
  NAND2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U894 ( .A1(n807), .A2(n806), .ZN(n818) );
  XOR2_X1 U895 ( .A(G2067), .B(KEYINPUT37), .Z(n808) );
  XNOR2_X1 U896 ( .A(KEYINPUT91), .B(n808), .ZN(n828) );
  NAND2_X1 U897 ( .A1(G140), .A2(n882), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G104), .A2(n883), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U900 ( .A(KEYINPUT34), .B(n811), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G128), .A2(n878), .ZN(n813) );
  NAND2_X1 U902 ( .A1(G116), .A2(n879), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U904 ( .A(KEYINPUT35), .B(n814), .Z(n815) );
  NOR2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U906 ( .A(KEYINPUT36), .B(n817), .ZN(n899) );
  NOR2_X1 U907 ( .A1(n828), .A2(n899), .ZN(n1008) );
  NAND2_X1 U908 ( .A1(n1008), .A2(n830), .ZN(n827) );
  NAND2_X1 U909 ( .A1(n818), .A2(n827), .ZN(n834) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n893), .ZN(n990) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n889), .ZN(n1003) );
  NOR2_X1 U913 ( .A1(n819), .A2(n1003), .ZN(n820) );
  NOR2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U915 ( .A(KEYINPUT105), .B(n822), .Z(n823) );
  NOR2_X1 U916 ( .A1(n990), .A2(n823), .ZN(n824) );
  XOR2_X1 U917 ( .A(KEYINPUT106), .B(n824), .Z(n825) );
  XOR2_X1 U918 ( .A(KEYINPUT39), .B(n825), .Z(n826) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n828), .A2(n899), .ZN(n993) );
  NAND2_X1 U921 ( .A1(n829), .A2(n993), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U923 ( .A(KEYINPUT107), .B(n832), .Z(n833) );
  NAND2_X1 U924 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U925 ( .A(n835), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U926 ( .A(G301), .ZN(G171) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n836), .ZN(G217) );
  INV_X1 U928 ( .A(n836), .ZN(G223) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U930 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U932 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U933 ( .A(n840), .ZN(G319) );
  INV_X1 U935 ( .A(G108), .ZN(G238) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  NOR2_X1 U937 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XOR2_X1 U939 ( .A(KEYINPUT41), .B(G1976), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n845), .B(G2474), .Z(n847) );
  XNOR2_X1 U943 ( .A(G1956), .B(G1981), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U945 ( .A(G1986), .B(G1971), .Z(n849) );
  XNOR2_X1 U946 ( .A(G1966), .B(G1961), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U948 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U949 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U951 ( .A(G2096), .B(G2100), .Z(n855) );
  XNOR2_X1 U952 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(KEYINPUT43), .B(G2090), .Z(n857) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U958 ( .A(G2084), .B(G2078), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(G227) );
  NAND2_X1 U960 ( .A1(G112), .A2(n879), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G100), .A2(n883), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(KEYINPUT112), .B(n864), .ZN(n870) );
  NAND2_X1 U964 ( .A1(n878), .A2(G124), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G136), .A2(n882), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(KEYINPUT111), .B(n868), .Z(n869) );
  NOR2_X1 U969 ( .A1(n870), .A2(n869), .ZN(G162) );
  NAND2_X1 U970 ( .A1(G139), .A2(n882), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G103), .A2(n883), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G127), .A2(n878), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G115), .A2(n879), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n995) );
  NAND2_X1 U978 ( .A1(G130), .A2(n878), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G118), .A2(n879), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U981 ( .A1(G142), .A2(n882), .ZN(n885) );
  NAND2_X1 U982 ( .A1(G106), .A2(n883), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U984 ( .A(n886), .B(KEYINPUT45), .Z(n887) );
  NOR2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n995), .B(n891), .ZN(n895) );
  XOR2_X1 U988 ( .A(G160), .B(G162), .Z(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n901) );
  XOR2_X1 U991 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n897) );
  XNOR2_X1 U992 ( .A(G164), .B(n1002), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U997 ( .A(G286), .B(n979), .Z(n904) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U999 ( .A(n905), .B(G301), .Z(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n907), .B(KEYINPUT49), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n908), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n909), .A2(G319), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(KEYINPUT113), .B(n910), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1010 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1021) );
  XNOR2_X1 U1011 ( .A(G25), .B(G1991), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n913), .B(KEYINPUT117), .ZN(n923) );
  XOR2_X1 U1013 ( .A(G2072), .B(G33), .Z(n914) );
  NAND2_X1 U1014 ( .A1(n914), .A2(G28), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(G27), .B(n915), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(G2067), .B(G26), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G1996), .B(G32), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n924), .B(KEYINPUT53), .ZN(n927) );
  XOR2_X1 U1023 ( .A(G2084), .B(G34), .Z(n925) );
  XNOR2_X1 U1024 ( .A(KEYINPUT54), .B(n925), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(G35), .B(G2090), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(n930), .B(KEYINPUT118), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(G29), .A2(n931), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT55), .B(n932), .ZN(n1019) );
  XOR2_X1 U1031 ( .A(G1961), .B(G5), .Z(n942) );
  XNOR2_X1 U1032 ( .A(G1348), .B(KEYINPUT59), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(n933), .B(G4), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(G1341), .B(G19), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(G1981), .B(G6), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(G20), .B(G1956), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT60), .B(n940), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(G21), .B(G1966), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT123), .B(n945), .ZN(n953) );
  XOR2_X1 U1045 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n951) );
  XOR2_X1 U1046 ( .A(G1986), .B(G24), .Z(n949) );
  XNOR2_X1 U1047 ( .A(G1971), .B(G22), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(G23), .B(G1976), .ZN(n946) );
  NOR2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1051 ( .A(n951), .B(n950), .Z(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1053 ( .A(KEYINPUT61), .B(n954), .Z(n956) );
  XNOR2_X1 U1054 ( .A(G16), .B(KEYINPUT122), .ZN(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(KEYINPUT125), .B(n957), .ZN(n987) );
  XNOR2_X1 U1057 ( .A(KEYINPUT56), .B(G16), .ZN(n985) );
  XOR2_X1 U1058 ( .A(G1966), .B(G168), .Z(n958) );
  XNOR2_X1 U1059 ( .A(KEYINPUT119), .B(n958), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1061 ( .A(n961), .B(KEYINPUT57), .ZN(n983) );
  XOR2_X1 U1062 ( .A(n962), .B(G1956), .Z(n964) );
  XOR2_X1 U1063 ( .A(G166), .B(G1971), .Z(n963) );
  NOR2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n972) );
  INV_X1 U1065 ( .A(n965), .ZN(n967) );
  NAND2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(KEYINPUT120), .B(n968), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(n973), .B(KEYINPUT121), .ZN(n978) );
  XOR2_X1 U1071 ( .A(G171), .B(G1961), .Z(n976) );
  XNOR2_X1 U1072 ( .A(n974), .B(G1341), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1075 ( .A(G1348), .B(n979), .Z(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(n988), .B(KEYINPUT126), .ZN(n1017) );
  XOR2_X1 U1081 ( .A(G2090), .B(G162), .Z(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1083 ( .A(KEYINPUT114), .B(n991), .Z(n992) );
  XNOR2_X1 U1084 ( .A(n992), .B(KEYINPUT51), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G2072), .B(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G164), .B(G2078), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1089 ( .A(KEYINPUT50), .B(n998), .Z(n999) );
  XNOR2_X1 U1090 ( .A(KEYINPUT115), .B(n999), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1011) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  XOR2_X1 U1093 ( .A(G160), .B(G2084), .Z(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1012), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1013), .B(KEYINPUT116), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(G29), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(G11), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(n1021), .B(n1020), .Z(G150) );
  INV_X1 U1105 ( .A(G150), .ZN(G311) );
endmodule

