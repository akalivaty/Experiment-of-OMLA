//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1134, new_n1135, new_n1136;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n454), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2106), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT66), .Z(G319));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(new_n465), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n474), .B2(new_n468), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G125), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n471), .B1(new_n475), .B2(new_n481), .ZN(G160));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n476), .A2(new_n477), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(KEYINPUT68), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n464), .A2(KEYINPUT68), .A3(new_n465), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(new_n468), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(new_n490), .B2(G124), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n489), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NOR2_X1   g070(.A1(new_n468), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n468), .A2(G138), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n503), .B2(new_n473), .ZN(new_n504));
  OAI211_X1 g079(.A(G138), .B(new_n468), .C1(new_n476), .C2(new_n477), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n501), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT70), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n513), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(new_n509), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(new_n530), .B1(new_n520), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  INV_X1    g109(.A(new_n514), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n532), .B1(new_n521), .B2(new_n533), .C1(new_n534), .C2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n512), .A2(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(G651), .B1(G90), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n514), .A2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AOI22_X1  g119(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n525), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT71), .B(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n514), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n540), .A2(G81), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n514), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n518), .A2(new_n519), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(G91), .B2(new_n540), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n540), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n514), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  AOI22_X1  g144(.A1(new_n540), .A2(G86), .B1(new_n514), .B2(G48), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT72), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n560), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n571), .B1(new_n574), .B2(G651), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR3_X1   g151(.A1(new_n576), .A2(KEYINPUT72), .A3(new_n525), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n570), .B1(new_n575), .B2(new_n577), .ZN(G305));
  NAND2_X1  g153(.A1(new_n540), .A2(G85), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n514), .A2(G47), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n525), .C2(new_n581), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT73), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n540), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n560), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(new_n592), .B2(G868), .ZN(G284));
  XOR2_X1   g168(.A(G284), .B(KEYINPUT74), .Z(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  NOR2_X1   g175(.A1(new_n551), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n592), .A2(new_n599), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT75), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n492), .A2(G135), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n490), .A2(G123), .ZN(new_n607));
  OR2_X1    g182(.A1(G99), .A2(G2105), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n608), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT77), .B(G2096), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n473), .A2(new_n469), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT76), .B(G2100), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n616), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT78), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2427), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT79), .ZN(new_n625));
  OAI21_X1  g200(.A(KEYINPUT14), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT80), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n625), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n635), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT81), .Z(new_n641));
  NOR2_X1   g216(.A1(G2072), .A2(G2078), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n444), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n639), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(KEYINPUT17), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n639), .B(new_n640), .C1(new_n444), .C2(new_n642), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT18), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n645), .A2(new_n641), .A3(new_n639), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n654));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT20), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n659), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n661), .B(new_n664), .C1(new_n656), .C2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1981), .B(G1986), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT83), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n668), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G29), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G35), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G162), .B2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT29), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2090), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT91), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G29), .B2(G32), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n492), .A2(G141), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n490), .A2(G129), .ZN(new_n682));
  NAND3_X1  g257(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT26), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  AOI22_X1  g261(.A1(new_n685), .A2(new_n686), .B1(G105), .B2(new_n469), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n681), .A2(new_n682), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(new_n674), .ZN(new_n689));
  MUX2_X1   g264(.A(new_n680), .B(new_n679), .S(new_n689), .Z(new_n690));
  XOR2_X1   g265(.A(KEYINPUT27), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(G27), .A2(G29), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G164), .B2(G29), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n611), .A2(G29), .B1(G2078), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n696), .A2(G28), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n674), .B1(new_n696), .B2(G28), .ZN(new_n698));
  AND2_X1   g273(.A1(KEYINPUT31), .A2(G11), .ZN(new_n699));
  NOR2_X1   g274(.A1(KEYINPUT31), .A2(G11), .ZN(new_n700));
  OAI22_X1  g275(.A1(new_n697), .A2(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n694), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n443), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT92), .B(G1956), .Z(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G20), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT23), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n596), .B2(new_n705), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n695), .B(new_n703), .C1(new_n704), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n704), .B2(new_n708), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n678), .A2(new_n692), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n674), .A2(G33), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n492), .A2(G139), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT25), .Z(new_n715));
  AOI22_X1  g290(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n713), .B(new_n715), .C1(new_n468), .C2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n712), .B1(new_n717), .B2(G29), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(new_n442), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT90), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT24), .ZN(new_n721));
  INV_X1    g296(.A(G34), .ZN(new_n722));
  AOI21_X1  g297(.A(G29), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n721), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G160), .B2(new_n674), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G2084), .Z(new_n726));
  XOR2_X1   g301(.A(KEYINPUT89), .B(G2067), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n674), .A2(G26), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n490), .A2(G128), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n733));
  INV_X1    g308(.A(G116), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n492), .A2(G140), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n732), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n729), .B1(new_n741), .B2(new_n674), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n720), .B(new_n726), .C1(new_n727), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n551), .A2(G16), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G16), .B2(G19), .ZN(new_n745));
  INV_X1    g320(.A(G1341), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n718), .A2(new_n442), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G168), .A2(new_n705), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n705), .B2(G21), .ZN(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n705), .A2(G5), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G171), .B2(new_n705), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G1961), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI22_X1  g334(.A1(new_n752), .A2(new_n753), .B1(G1961), .B2(new_n756), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n750), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n705), .A2(G4), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n592), .B2(new_n705), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT86), .B(G1348), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n742), .A2(new_n727), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n761), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n711), .A2(new_n743), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT93), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT85), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n674), .A2(G25), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n492), .A2(G131), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n490), .A2(G119), .ZN(new_n773));
  OR2_X1    g348(.A1(G95), .A2(G2105), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n771), .B1(new_n777), .B2(new_n674), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT35), .B(G1991), .Z(new_n779));
  XOR2_X1   g354(.A(new_n778), .B(new_n779), .Z(new_n780));
  MUX2_X1   g355(.A(G6), .B(G305), .S(G16), .Z(new_n781));
  XOR2_X1   g356(.A(KEYINPUT32), .B(G1981), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n705), .A2(G22), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G166), .B2(new_n705), .ZN(new_n785));
  INV_X1    g360(.A(G1971), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G23), .B(G288), .S(G16), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n783), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n770), .B(new_n780), .C1(new_n791), .C2(KEYINPUT34), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G24), .ZN(new_n793));
  XNOR2_X1  g368(.A(G290), .B(KEYINPUT84), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1986), .Z(new_n796));
  OAI211_X1 g371(.A(new_n792), .B(new_n796), .C1(KEYINPUT34), .C2(new_n791), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT36), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n769), .A2(new_n798), .ZN(G150));
  INV_X1    g374(.A(G150), .ZN(G311));
  INV_X1    g375(.A(G67), .ZN(new_n801));
  INV_X1    g376(.A(G80), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n560), .A2(new_n801), .B1(new_n802), .B2(new_n509), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT94), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n805), .B1(new_n802), .B2(new_n509), .C1(new_n560), .C2(new_n801), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n804), .A2(G651), .A3(new_n806), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n540), .A2(G93), .B1(new_n514), .B2(G55), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT95), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(new_n550), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n551), .A2(new_n807), .A3(new_n808), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n592), .A2(G559), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT96), .Z(new_n820));
  AOI21_X1  g395(.A(G860), .B1(new_n817), .B2(new_n818), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n811), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(G145));
  XNOR2_X1  g400(.A(new_n740), .B(new_n688), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n776), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n507), .B(KEYINPUT97), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n717), .B(new_n828), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n492), .A2(G142), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n490), .A2(G130), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n468), .A2(G118), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n616), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n829), .B(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n827), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n827), .A2(new_n836), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n494), .B(new_n610), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G160), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(G37), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n839), .A2(KEYINPUT98), .A3(new_n842), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n827), .B(new_n836), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n841), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n843), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g424(.A(G868), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n811), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(G305), .B(G303), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(G290), .B(G288), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(KEYINPUT100), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT42), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n591), .B(new_n596), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT41), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n814), .B(new_n602), .ZN(new_n865));
  MUX2_X1   g440(.A(new_n864), .B(new_n863), .S(new_n865), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n862), .B(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n851), .B1(new_n867), .B2(new_n850), .ZN(G295));
  OAI21_X1  g443(.A(new_n851), .B1(new_n867), .B2(new_n850), .ZN(G331));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n870));
  XNOR2_X1  g445(.A(G301), .B(G286), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n814), .B(new_n871), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n863), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n814), .B(new_n871), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n864), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n859), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n860), .A3(new_n875), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(KEYINPUT43), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n876), .B2(new_n859), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n879), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n870), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n880), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT102), .B1(new_n880), .B2(KEYINPUT43), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT101), .B1(new_n880), .B2(KEYINPUT43), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n883), .A2(new_n890), .A3(new_n882), .A4(new_n879), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(KEYINPUT44), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n885), .B1(new_n888), .B2(new_n892), .ZN(G397));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(G1384), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n496), .A2(new_n497), .ZN(new_n896));
  INV_X1    g471(.A(new_n499), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT4), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(KEYINPUT69), .ZN(new_n899));
  INV_X1    g474(.A(G138), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(G2105), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n897), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n896), .B1(new_n902), .B2(new_n486), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n899), .B1(new_n466), .B2(G138), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n895), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G1384), .B1(new_n504), .B2(new_n506), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(KEYINPUT45), .ZN(new_n907));
  INV_X1    g482(.A(new_n471), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT67), .B1(new_n480), .B2(G2105), .ZN(new_n909));
  AOI211_X1 g484(.A(new_n472), .B(new_n468), .C1(new_n478), .C2(new_n479), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n908), .B(G40), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT53), .B1(new_n912), .B2(new_n443), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n913), .A2(KEYINPUT122), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(KEYINPUT122), .ZN(new_n915));
  INV_X1    g490(.A(G40), .ZN(new_n916));
  AOI211_X1 g491(.A(new_n916), .B(new_n471), .C1(new_n475), .C2(new_n481), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT50), .ZN(new_n918));
  INV_X1    g493(.A(G1384), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n507), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI211_X1 g496(.A(KEYINPUT50), .B(G1384), .C1(new_n504), .C2(new_n506), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n917), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n758), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n914), .A2(new_n915), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G301), .B(KEYINPUT54), .ZN(new_n927));
  INV_X1    g502(.A(new_n907), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n443), .A2(KEYINPUT53), .A3(G40), .ZN(new_n929));
  AOI211_X1 g504(.A(new_n929), .B(new_n471), .C1(G2105), .C2(new_n480), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n919), .B1(new_n903), .B2(new_n904), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n894), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n905), .A2(KEYINPUT109), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n507), .A2(new_n935), .A3(new_n895), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(new_n911), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n914), .A2(new_n915), .A3(new_n925), .A4(new_n939), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n926), .A2(new_n931), .B1(new_n940), .B2(new_n927), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n786), .B1(new_n907), .B2(new_n911), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT103), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(new_n786), .C1(new_n907), .C2(new_n911), .ZN(new_n945));
  XOR2_X1   g520(.A(KEYINPUT104), .B(G2090), .Z(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n917), .A2(new_n921), .A3(new_n923), .A4(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n943), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G8), .ZN(new_n950));
  NOR2_X1   g525(.A1(G166), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n952), .A3(G8), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n949), .A2(new_n952), .A3(KEYINPUT105), .A4(G8), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(KEYINPUT106), .B(G8), .C1(new_n911), .C2(new_n932), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n475), .A2(new_n481), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(G40), .A3(new_n906), .A4(new_n908), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT106), .B1(new_n961), .B2(G8), .ZN(new_n962));
  INV_X1    g537(.A(G1981), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n963), .B(new_n570), .C1(new_n575), .C2(new_n577), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n514), .A2(G48), .ZN(new_n966));
  XNOR2_X1  g541(.A(KEYINPUT107), .B(G86), .ZN(new_n967));
  OAI221_X1 g542(.A(new_n966), .B1(new_n521), .B2(new_n967), .C1(new_n576), .C2(new_n525), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G1981), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n964), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n965), .B1(new_n964), .B2(new_n969), .ZN(new_n971));
  OAI22_X1  g546(.A1(new_n959), .A2(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1976), .ZN(new_n973));
  NOR2_X1   g548(.A1(G288), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT52), .B1(G288), .B2(new_n973), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n975), .B(new_n976), .C1(new_n959), .C2(new_n962), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n911), .A2(new_n932), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n978), .B1(new_n979), .B2(new_n950), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n974), .B1(new_n980), .B2(new_n958), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n972), .B(new_n977), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n948), .A2(new_n942), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n952), .B1(G8), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT123), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n957), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n987), .B1(new_n957), .B2(new_n986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n941), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n753), .B1(new_n937), .B2(new_n911), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT110), .B(G2084), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n917), .A2(new_n921), .A3(new_n923), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n950), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n995));
  NAND3_X1  g570(.A1(G286), .A2(new_n995), .A3(G8), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n995), .B1(G286), .B2(G8), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT119), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n998), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT119), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n996), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT51), .B1(new_n994), .B2(new_n1003), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n997), .A2(KEYINPUT51), .A3(new_n998), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT120), .B1(new_n994), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n917), .A2(new_n933), .A3(new_n934), .A4(new_n936), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n911), .A2(new_n920), .A3(new_n922), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1009), .A2(new_n753), .B1(new_n1010), .B2(new_n992), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1008), .B(new_n1005), .C1(new_n1011), .C2(new_n950), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1004), .A2(new_n1007), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1011), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n997), .B2(new_n998), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1013), .A2(KEYINPUT121), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT121), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT124), .B1(new_n990), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT61), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n1021));
  NOR3_X1   g596(.A1(G299), .A2(KEYINPUT114), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n596), .B2(KEYINPUT57), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n563), .A2(KEYINPUT113), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n558), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n563), .A2(KEYINPUT113), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1021), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1022), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT115), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT111), .B(G1956), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n924), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n924), .A2(KEYINPUT112), .A3(new_n1031), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT56), .B(G2072), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n912), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n912), .A2(KEYINPUT116), .A3(new_n1037), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1030), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1029), .B(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1020), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1030), .A2(new_n1043), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(KEYINPUT61), .ZN(new_n1052));
  INV_X1    g627(.A(G1996), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n912), .A2(new_n1053), .ZN(new_n1054));
  OR2_X1    g629(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1055));
  NAND2_X1  g630(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n961), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n550), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n1058), .B(new_n1059), .Z(new_n1060));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n1061));
  INV_X1    g636(.A(G2067), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n924), .A2(new_n764), .B1(new_n1062), .B2(new_n979), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1063), .A2(new_n591), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n591), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1063), .A2(new_n1061), .A3(new_n592), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1060), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1049), .A2(new_n1052), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1064), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1048), .B1(new_n1051), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n957), .A2(new_n986), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT123), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n957), .A2(new_n986), .A3(new_n987), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1013), .A2(KEYINPUT121), .A3(new_n1015), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1076), .A2(new_n1081), .A3(new_n1082), .A4(new_n941), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1019), .A2(new_n1072), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G288), .A2(G1976), .ZN(new_n1085));
  XOR2_X1   g660(.A(new_n1085), .B(KEYINPUT108), .Z(new_n1086));
  NOR3_X1   g661(.A1(new_n1086), .A2(new_n971), .A3(new_n970), .ZN(new_n1087));
  INV_X1    g662(.A(new_n964), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n958), .B2(new_n980), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n994), .A2(G168), .ZN(new_n1091));
  OR3_X1    g666(.A1(new_n1091), .A2(new_n985), .A3(KEYINPUT63), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n983), .B1(new_n1092), .B2(new_n957), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n952), .B1(new_n949), .B2(G8), .ZN(new_n1094));
  OR3_X1    g669(.A1(new_n983), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n1090), .B(new_n1093), .C1(KEYINPUT63), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1079), .A2(KEYINPUT62), .A3(new_n1080), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n940), .A2(G171), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1100), .A2(KEYINPUT125), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT125), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1084), .B(new_n1096), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n911), .A2(new_n933), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n741), .A2(new_n1062), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n740), .A2(G2067), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n688), .B(new_n1053), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n777), .A2(new_n779), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n777), .A2(new_n779), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G290), .B(G1986), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1106), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1105), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1106), .B1(new_n1117), .B2(new_n688), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1106), .A2(new_n1053), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT46), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1121), .B(KEYINPUT47), .Z(new_n1122));
  NAND2_X1  g697(.A1(new_n1113), .A2(new_n1106), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT126), .ZN(new_n1124));
  NOR2_X1   g699(.A1(G290), .A2(G1986), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1106), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n1126), .B(KEYINPUT48), .Z(new_n1127));
  NOR2_X1   g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1107), .B1(new_n1129), .B2(new_n1111), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1122), .B(new_n1128), .C1(new_n1106), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1116), .A2(new_n1131), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g707(.A1(new_n652), .A2(new_n462), .ZN(new_n1134));
  XNOR2_X1  g708(.A(new_n1134), .B(KEYINPUT127), .ZN(new_n1135));
  NOR3_X1   g709(.A1(G401), .A2(G229), .A3(new_n1135), .ZN(new_n1136));
  OAI211_X1 g710(.A(new_n848), .B(new_n1136), .C1(new_n884), .C2(new_n881), .ZN(G225));
  INV_X1    g711(.A(G225), .ZN(G308));
endmodule


