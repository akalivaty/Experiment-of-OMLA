//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n204), .B(new_n206), .C1(new_n202), .C2(new_n203), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT96), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(G50gat), .ZN(new_n211));
  INV_X1    g010(.A(G50gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT96), .A3(G43gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT95), .B(KEYINPUT15), .Z(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(G43gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(new_n217), .A3(KEYINPUT15), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n207), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n207), .A2(new_n218), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OR3_X1    g020(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT17), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT16), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n223), .A2(G1gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(G8gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT17), .B1(new_n219), .B2(new_n221), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n222), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n228), .B(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n219), .A2(new_n221), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n231), .A2(new_n235), .A3(KEYINPUT18), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT97), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n238), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n236), .B(KEYINPUT13), .Z(new_n241));
  INV_X1    g040(.A(new_n235), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n233), .A2(new_n234), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT11), .B(G169gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT12), .Z(new_n249));
  NAND4_X1  g048(.A1(new_n239), .A2(new_n240), .A3(new_n244), .A4(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n235), .A3(new_n236), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT98), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n251), .A2(new_n253), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n239), .A2(new_n240), .A3(new_n244), .A4(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n249), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT90), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT39), .ZN(new_n266));
  XNOR2_X1  g065(.A(G127gat), .B(G134gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  INV_X1    g069(.A(G113gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(G120gat), .ZN(new_n272));
  INV_X1    g071(.A(G120gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(G113gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G127gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n269), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT69), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n274), .A2(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(KEYINPUT70), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n280), .B(new_n281), .C1(new_n271), .C2(G120gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n270), .A3(new_n267), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G155gat), .B(G162gat), .ZN(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  INV_X1    g086(.A(G162gat), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT2), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G148gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G141gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT77), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n290), .A2(G141gat), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n286), .B(new_n289), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n290), .A2(G141gat), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT2), .B1(new_n295), .B2(new_n291), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n296), .A2(new_n286), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n285), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT4), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n299), .A2(KEYINPUT79), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n294), .A2(KEYINPUT79), .A3(new_n297), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n285), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n305), .A3(KEYINPUT81), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n298), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n278), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n283), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n300), .A2(new_n313), .A3(KEYINPUT4), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n306), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n316));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n317), .B(KEYINPUT78), .Z(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n316), .B1(new_n315), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n266), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT88), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n311), .A2(new_n298), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n300), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n318), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(new_n266), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n319), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G85gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT0), .B(G57gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  XOR2_X1   g132(.A(new_n333), .B(KEYINPUT87), .Z(new_n334));
  NAND3_X1  g133(.A1(new_n322), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT40), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(G169gat), .B2(G176gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT65), .ZN(new_n340));
  INV_X1    g139(.A(G183gat), .ZN(new_n341));
  INV_X1    g140(.A(G190gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT24), .ZN(new_n345));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n345), .ZN(new_n347));
  OAI221_X1 g146(.A(new_n343), .B1(new_n344), .B2(new_n345), .C1(new_n347), .C2(KEYINPUT67), .ZN(new_n348));
  OR3_X1    g147(.A1(new_n338), .A2(G169gat), .A3(G176gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n340), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n351), .B(KEYINPUT66), .Z(new_n352));
  OAI21_X1  g151(.A(KEYINPUT25), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NOR3_X1   g152(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n351), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT27), .B(G183gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT28), .A3(new_n342), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT28), .B1(new_n357), .B2(new_n342), .ZN(new_n360));
  OAI221_X1 g159(.A(new_n346), .B1(new_n354), .B2(new_n356), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n343), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT64), .B(G176gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n338), .A2(G169gat), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT25), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n340), .A2(new_n351), .A3(new_n363), .A4(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n353), .A2(new_n361), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G226gat), .ZN(new_n369));
  INV_X1    g168(.A(G233gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT75), .ZN(new_n374));
  XNOR2_X1  g173(.A(G197gat), .B(G204gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT74), .B(G218gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(KEYINPUT22), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G211gat), .ZN(new_n378));
  INV_X1    g177(.A(G211gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(KEYINPUT22), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(G218gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n371), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n374), .A2(new_n382), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT76), .B1(new_n384), .B2(new_n385), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n391));
  AOI211_X1 g190(.A(new_n391), .B(new_n371), .C1(new_n368), .C2(new_n383), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n390), .A2(new_n392), .A3(new_n373), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n389), .B1(new_n393), .B2(new_n382), .ZN(new_n394));
  XNOR2_X1  g193(.A(G8gat), .B(G36gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n389), .B(new_n397), .C1(new_n393), .C2(new_n382), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT30), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(new_n402), .A3(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n337), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n326), .A2(new_n318), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n409));
  INV_X1    g208(.A(new_n318), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n300), .B2(new_n325), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n312), .A2(KEYINPUT4), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n318), .B1(new_n414), .B2(new_n300), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n285), .B(KEYINPUT4), .C1(new_n303), .C2(new_n304), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n408), .A2(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n318), .A2(KEYINPUT5), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n306), .A2(new_n312), .A3(new_n314), .A4(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT89), .B1(new_n421), .B2(new_n334), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n408), .A2(new_n413), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n415), .A2(new_n416), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n419), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT89), .ZN(new_n427));
  INV_X1    g226(.A(new_n334), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n422), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n322), .A2(new_n329), .A3(KEYINPUT40), .A4(new_n334), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n265), .B1(new_n406), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n404), .B1(new_n335), .B2(new_n336), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n434), .A2(KEYINPUT90), .A3(new_n430), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT6), .B1(new_n421), .B2(new_n333), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n427), .B1(new_n426), .B2(new_n428), .ZN(new_n438));
  AOI211_X1 g237(.A(KEYINPUT89), .B(new_n334), .C1(new_n425), .C2(new_n419), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT91), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n430), .A2(KEYINPUT91), .A3(new_n437), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT93), .B(KEYINPUT37), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n398), .B1(new_n394), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(new_n394), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT92), .B(KEYINPUT38), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n393), .A2(new_n382), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n374), .A2(new_n386), .A3(new_n388), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n452), .B(KEYINPUT37), .C1(new_n382), .C2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n446), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n450), .A2(new_n399), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n333), .ZN(new_n457));
  OAI211_X1 g256(.A(KEYINPUT6), .B(new_n457), .C1(new_n417), .C2(new_n420), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT83), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n426), .A2(new_n460), .A3(KEYINPUT6), .A4(new_n457), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT94), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n456), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G228gat), .A2(G233gat), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n307), .B1(new_n382), .B2(KEYINPUT29), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n303), .A2(new_n304), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT84), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n383), .B1(new_n298), .B2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n382), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n468), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n468), .B1(new_n469), .B2(new_n298), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n474), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT85), .ZN(new_n479));
  XNOR2_X1  g278(.A(G78gat), .B(G106gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT31), .B(G50gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(KEYINPUT86), .A3(G22gat), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(G22gat), .B2(new_n482), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n476), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n476), .B2(new_n479), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n436), .A2(new_n467), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G227gat), .A2(G233gat), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n368), .A2(new_n311), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n368), .A2(new_n311), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n493), .A2(KEYINPUT33), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT32), .B1(new_n495), .B2(new_n490), .ZN(new_n496));
  XOR2_X1   g295(.A(G15gat), .B(G43gat), .Z(new_n497));
  XNOR2_X1  g296(.A(G71gat), .B(G99gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT71), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT32), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(KEYINPUT33), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n494), .A2(new_n496), .A3(new_n501), .A4(new_n499), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n495), .A2(new_n490), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT34), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n506), .A2(new_n514), .A3(new_n507), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n513), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n508), .A3(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(KEYINPUT36), .A3(new_n518), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n459), .A2(new_n461), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT82), .B1(new_n421), .B2(new_n333), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT82), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n426), .A2(new_n525), .A3(new_n457), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n437), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n405), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n521), .B(new_n522), .C1(new_n528), .C2(new_n488), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n489), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n444), .A2(new_n466), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT35), .ZN(new_n533));
  AOI211_X1 g332(.A(new_n487), .B(new_n405), .C1(new_n516), .C2(new_n518), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n528), .A2(new_n488), .A3(new_n519), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n264), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G127gat), .B(G155gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G211gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G64gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G57gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT100), .B(G57gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(new_n543), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n547), .A2(G71gat), .A3(G78gat), .ZN(new_n548));
  AND2_X1   g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n552));
  INV_X1    g351(.A(G57gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(G64gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n543), .A2(G57gat), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT9), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n552), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n553), .A2(G64gat), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n547), .B1(new_n544), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G71gat), .B(G78gat), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n561), .A2(KEYINPUT99), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n551), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT21), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT101), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT99), .B1(new_n561), .B2(new_n562), .ZN(new_n570));
  XNOR2_X1  g369(.A(G57gat), .B(G64gat), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n558), .B(new_n552), .C1(new_n571), .C2(new_n547), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(KEYINPUT101), .A3(new_n551), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n567), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(new_n233), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n341), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n576), .A2(new_n341), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n566), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n578), .A2(new_n579), .A3(new_n566), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n580), .A2(G231gat), .A3(G233gat), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n580), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(new_n581), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n542), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n542), .A3(new_n586), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n222), .A2(new_n230), .ZN(new_n594));
  OR2_X1    g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  INV_X1    g394(.A(G99gat), .ZN(new_n596));
  INV_X1    g395(.A(G106gat), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT8), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n599), .A2(KEYINPUT7), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(KEYINPUT7), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n595), .B(new_n598), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G99gat), .B(G106gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n599), .B(KEYINPUT7), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n606), .A2(new_n603), .A3(new_n595), .A4(new_n598), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n594), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT103), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n234), .A2(new_n607), .A3(new_n605), .ZN(new_n613));
  OR3_X1    g412(.A1(new_n594), .A2(new_n610), .A3(KEYINPUT103), .ZN(new_n614));
  AND2_X1   g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n612), .A2(new_n613), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n611), .A2(KEYINPUT103), .B1(KEYINPUT41), .B2(new_n615), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n621), .A2(new_n613), .A3(new_n614), .A4(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT104), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT105), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT104), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n626), .A3(new_n622), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n628));
  XNOR2_X1  g427(.A(G134gat), .B(G162gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n623), .A2(KEYINPUT104), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n625), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n627), .A2(new_n630), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n623), .B2(KEYINPUT104), .ZN(new_n636));
  AOI211_X1 g435(.A(new_n626), .B(KEYINPUT105), .C1(new_n620), .C2(new_n622), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n593), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT106), .Z(new_n644));
  NAND3_X1  g443(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT10), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n573), .A2(KEYINPUT101), .A3(new_n551), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT101), .B1(new_n573), .B2(new_n551), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n564), .A2(new_n608), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n573), .A2(new_n551), .A3(new_n607), .A4(new_n605), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n644), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n644), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(new_n650), .B2(new_n652), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n654), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n649), .A2(new_n653), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(new_n655), .ZN(new_n663));
  AOI211_X1 g462(.A(KEYINPUT107), .B(new_n644), .C1(new_n649), .C2(new_n653), .ZN(new_n664));
  OR3_X1    g463(.A1(new_n663), .A2(new_n664), .A3(new_n656), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n660), .B1(new_n665), .B2(new_n659), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n539), .A2(new_n642), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n523), .A2(new_n527), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n224), .ZN(G1324gat));
  NOR2_X1   g470(.A1(new_n667), .A2(new_n404), .ZN(new_n672));
  AND2_X1   g471(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n672), .A2(KEYINPUT42), .A3(new_n674), .A4(new_n676), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n679), .B(new_n680), .C1(new_n232), .C2(new_n672), .ZN(G1325gat));
  INV_X1    g480(.A(G15gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n521), .A2(new_n522), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT108), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n667), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n539), .A2(new_n519), .A3(new_n642), .A4(new_n666), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n682), .B2(new_n686), .ZN(G1326gat));
  OR3_X1    g486(.A1(new_n667), .A2(G22gat), .A3(new_n488), .ZN(new_n688));
  OAI21_X1  g487(.A(G22gat), .B1(new_n667), .B2(new_n488), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(new_n691), .A3(new_n689), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1327gat));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n489), .A2(new_n530), .B1(new_n535), .B2(new_n537), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(new_n640), .ZN(new_n698));
  INV_X1    g497(.A(new_n666), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n593), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n487), .B1(new_n433), .B2(new_n435), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n529), .B1(new_n701), .B2(new_n467), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT35), .B1(new_n444), .B2(new_n466), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n703), .A2(new_n534), .B1(KEYINPUT35), .B2(new_n536), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT44), .B(new_n639), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n263), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n258), .A2(KEYINPUT110), .A3(new_n262), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n698), .A2(new_n700), .A3(new_n705), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G29gat), .B1(new_n710), .B2(new_n669), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n263), .B(new_n700), .C1(new_n702), .C2(new_n704), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n640), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n202), .A3(new_n668), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(KEYINPUT45), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(KEYINPUT45), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(G1328gat));
  NAND3_X1  g516(.A1(new_n713), .A2(new_n203), .A3(new_n405), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n719));
  OAI21_X1  g518(.A(G36gat), .B1(new_n710), .B2(new_n404), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(G1329gat));
  AOI21_X1  g521(.A(G43gat), .B1(new_n516), .B2(new_n518), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n539), .A2(new_n639), .A3(new_n700), .A4(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n712), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n727), .A2(KEYINPUT111), .A3(new_n639), .A4(new_n723), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n726), .A2(new_n728), .B1(KEYINPUT112), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n683), .ZN(new_n731));
  OAI21_X1  g530(.A(G43gat), .B1(new_n710), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n726), .A2(new_n728), .A3(KEYINPUT112), .ZN(new_n734));
  OAI21_X1  g533(.A(G43gat), .B1(new_n710), .B2(new_n684), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n736), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g536(.A(G50gat), .B1(new_n710), .B2(new_n488), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n713), .A2(new_n212), .A3(new_n487), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1331gat));
  NOR2_X1   g544(.A1(new_n697), .A2(new_n641), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n709), .A2(new_n666), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n669), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(new_n545), .Z(G1332gat));
  NOR2_X1   g549(.A1(new_n748), .A2(new_n404), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  OAI21_X1  g554(.A(G71gat), .B1(new_n748), .B2(new_n684), .ZN(new_n756));
  INV_X1    g555(.A(G71gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n519), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n748), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1334gat));
  NOR2_X1   g560(.A1(new_n748), .A2(new_n488), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT114), .B(G78gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n593), .A2(new_n666), .A3(new_n709), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n698), .A2(new_n705), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(G85gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n766), .A2(new_n767), .A3(new_n669), .ZN(new_n768));
  INV_X1    g567(.A(new_n709), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n639), .B(new_n769), .C1(new_n702), .C2(new_n704), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n591), .A2(new_n592), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT51), .B1(new_n770), .B2(new_n593), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n699), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n776), .A2(new_n669), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n768), .B1(new_n777), .B2(new_n767), .ZN(G1336gat));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n698), .A2(new_n405), .A3(new_n705), .A4(new_n765), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n404), .A2(G92gat), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n774), .A2(new_n699), .A3(new_n775), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n781), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n785), .B(new_n781), .C1(new_n782), .C2(new_n779), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1337gat));
  OAI21_X1  g588(.A(G99gat), .B1(new_n766), .B2(new_n684), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n519), .A2(new_n596), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n776), .B2(new_n791), .ZN(G1338gat));
  NOR2_X1   g591(.A1(new_n488), .A2(G106gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n699), .A3(new_n775), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G106gat), .B1(new_n766), .B2(new_n488), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT53), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1339gat));
  INV_X1    g599(.A(new_n660), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n645), .B1(new_n569), .B2(new_n574), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n655), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n649), .A2(new_n653), .A3(new_n644), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n807), .A2(KEYINPUT116), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(KEYINPUT116), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n805), .A2(KEYINPUT107), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n654), .A2(new_n661), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT54), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n659), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n663), .B2(new_n664), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(KEYINPUT117), .A3(new_n659), .ZN(new_n818));
  AOI221_X4 g617(.A(new_n802), .B1(new_n808), .B2(new_n809), .C1(new_n815), .C2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n808), .A2(new_n809), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n817), .A2(KEYINPUT117), .A3(new_n659), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT117), .B1(new_n817), .B2(new_n659), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n802), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n709), .A2(new_n801), .A3(new_n820), .A4(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n248), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n242), .A2(new_n243), .A3(new_n241), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n236), .B1(new_n231), .B2(new_n235), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n258), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n666), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n639), .B1(new_n826), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n831), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n639), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n801), .A3(new_n825), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n773), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n593), .A2(new_n640), .A3(new_n666), .A4(new_n769), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n669), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n534), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n264), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n709), .A2(new_n271), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n842), .B2(new_n844), .ZN(G1340gat));
  NOR2_X1   g644(.A1(new_n842), .A2(new_n666), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(new_n273), .ZN(G1341gat));
  NOR2_X1   g646(.A1(new_n842), .A2(new_n773), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT118), .B1(KEYINPUT119), .B2(G127gat), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(KEYINPUT118), .B2(G127gat), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n848), .B2(new_n852), .ZN(G1342gat));
  AOI211_X1 g652(.A(new_n640), .B(new_n842), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n854));
  NOR2_X1   g653(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1343gat));
  NAND3_X1  g655(.A1(new_n731), .A2(new_n668), .A3(new_n404), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n488), .B1(new_n839), .B2(new_n840), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n815), .A2(new_n818), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT55), .B1(new_n861), .B2(new_n821), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT120), .B1(new_n819), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n260), .A2(new_n261), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n801), .B1(new_n864), .B2(new_n257), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n825), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT121), .B1(new_n868), .B2(new_n833), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n870), .B(new_n832), .C1(new_n863), .C2(new_n867), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n640), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT122), .ZN(new_n873));
  INV_X1    g672(.A(new_n838), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n875), .B(new_n640), .C1(new_n869), .C2(new_n871), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n773), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n488), .B1(new_n878), .B2(new_n840), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n263), .B(new_n860), .C1(new_n879), .C2(new_n859), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G141gat), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n839), .A2(new_n840), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n669), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n488), .B1(new_n841), .B2(KEYINPUT123), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n684), .A2(new_n404), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(G141gat), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT58), .B1(new_n888), .B2(new_n263), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n881), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n887), .A2(G141gat), .A3(new_n264), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n709), .B(new_n860), .C1(new_n879), .C2(new_n859), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(G141gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(new_n891), .B2(new_n894), .ZN(G1344gat));
  OR3_X1    g694(.A1(new_n887), .A2(G148gat), .A3(new_n666), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n699), .B(new_n860), .C1(new_n879), .C2(new_n859), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n897), .A2(new_n898), .A3(G148gat), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT57), .B1(new_n883), .B2(new_n488), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n593), .B1(new_n872), .B2(new_n874), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n641), .A2(new_n263), .A3(new_n699), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n859), .B(new_n487), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n857), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n699), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n898), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n896), .B1(new_n899), .B2(new_n907), .ZN(G1345gat));
  OAI21_X1  g707(.A(new_n860), .B1(new_n879), .B2(new_n859), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n287), .A3(new_n773), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n887), .A2(new_n773), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n287), .B2(new_n911), .ZN(G1346gat));
  NOR3_X1   g711(.A1(new_n909), .A2(new_n288), .A3(new_n640), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n887), .A2(new_n640), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n288), .B2(new_n914), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n668), .A2(new_n404), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n916), .A2(new_n519), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT124), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n487), .B1(new_n839), .B2(new_n840), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G169gat), .B1(new_n920), .B2(new_n264), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n919), .A2(new_n917), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n769), .A2(G169gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(G1348gat));
  NOR3_X1   g724(.A1(new_n920), .A2(new_n364), .A3(new_n666), .ZN(new_n926));
  AOI21_X1  g725(.A(G176gat), .B1(new_n922), .B2(new_n699), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1349gat));
  OAI21_X1  g729(.A(G183gat), .B1(new_n920), .B2(new_n773), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n922), .A2(new_n357), .A3(new_n593), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n931), .B(new_n932), .C1(KEYINPUT126), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(KEYINPUT126), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT127), .Z(new_n936));
  XNOR2_X1  g735(.A(new_n934), .B(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n342), .A3(new_n639), .ZN(new_n938));
  OAI21_X1  g737(.A(G190gat), .B1(new_n920), .B2(new_n640), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  AND2_X1   g741(.A1(new_n684), .A2(new_n916), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n904), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n264), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n858), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n769), .A2(G197gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NOR3_X1   g747(.A1(new_n946), .A2(G204gat), .A3(new_n666), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT62), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n904), .A2(new_n699), .A3(new_n943), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G204gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n904), .A2(new_n593), .A3(new_n943), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n593), .A2(new_n379), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n955), .A2(new_n956), .B1(new_n946), .B2(new_n957), .ZN(G1354gat));
  INV_X1    g757(.A(new_n944), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n639), .A2(new_n376), .ZN(new_n960));
  INV_X1    g759(.A(G218gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n639), .A3(new_n858), .ZN(new_n962));
  AOI22_X1  g761(.A1(new_n959), .A2(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G1355gat));
endmodule


