//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n809, new_n810, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917;
  AND2_X1   g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n202), .A2(new_n203), .B1(G169gat), .B2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G183gat), .B(G190gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n204), .B(new_n210), .C1(new_n203), .C2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT28), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT27), .B(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(new_n219), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n202), .B1(KEYINPUT26), .B2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n221), .A2(new_n224), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n219), .A2(G183gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n215), .A2(G190gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT24), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n232), .A2(new_n233), .A3(new_n210), .A4(new_n204), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n229), .A3(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(KEYINPUT65), .A2(G120gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(KEYINPUT65), .A2(G120gat), .ZN(new_n237));
  OAI21_X1  g036(.A(G113gat), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(G113gat), .B2(G120gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G113gat), .ZN(new_n244));
  INV_X1    g043(.A(G120gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G127gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(G134gat), .ZN(new_n248));
  INV_X1    g047(.A(G134gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(G127gat), .ZN(new_n250));
  OAI22_X1  g049(.A1(new_n240), .A2(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G227gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n214), .A2(new_n229), .A3(new_n252), .A4(new_n234), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT32), .ZN(new_n260));
  XOR2_X1   g059(.A(G71gat), .B(G99gat), .Z(new_n261));
  XNOR2_X1  g060(.A(G15gat), .B(G43gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT33), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n259), .B2(new_n264), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n260), .B(new_n263), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT34), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n258), .ZN(new_n271));
  INV_X1    g070(.A(new_n257), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI211_X1 g072(.A(KEYINPUT34), .B(new_n257), .C1(new_n254), .C2(new_n258), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n263), .A2(KEYINPUT33), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n259), .A2(KEYINPUT32), .A3(new_n276), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n269), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n269), .B2(new_n277), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G78gat), .B(G106gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G22gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G141gat), .B(G148gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT2), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(G155gat), .B2(G162gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n286), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G141gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G148gat), .ZN(new_n292));
  INV_X1    g091(.A(G148gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G141gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G155gat), .B(G162gat), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT2), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n290), .A2(new_n300), .A3(KEYINPUT73), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT73), .B1(new_n290), .B2(new_n300), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g102(.A1(G197gat), .A2(G204gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G197gat), .A2(G204gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G211gat), .A2(G218gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT22), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(KEYINPUT67), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n304), .A2(new_n305), .B1(new_n308), .B2(new_n307), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n312), .A2(new_n316), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(new_n316), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT80), .B1(new_n322), .B2(KEYINPUT29), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n303), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n290), .A2(new_n300), .A3(new_n320), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n290), .A2(new_n300), .A3(KEYINPUT74), .A4(new_n320), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(KEYINPUT69), .B(KEYINPUT29), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n329), .A2(new_n331), .B1(new_n316), .B2(new_n312), .ZN(new_n332));
  OAI211_X1 g131(.A(G228gat), .B(G233gat), .C1(new_n324), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n290), .A2(new_n300), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n314), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n330), .B1(new_n336), .B2(new_n311), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n310), .A2(KEYINPUT78), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n314), .A2(new_n335), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n313), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n320), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n337), .B2(new_n340), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n334), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n332), .ZN(new_n346));
  NAND2_X1  g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT31), .B(G50gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n333), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n333), .B2(new_n348), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n283), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n333), .A2(new_n348), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n349), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n333), .A2(new_n348), .A3(new_n350), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n282), .A3(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT35), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n280), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n361), .B(KEYINPUT68), .Z(new_n362));
  AOI21_X1  g161(.A(new_n322), .B1(new_n235), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT70), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n235), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n214), .A2(new_n229), .A3(KEYINPUT70), .A4(new_n234), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n367), .B2(new_n362), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n362), .A3(new_n366), .ZN(new_n369));
  INV_X1    g168(.A(new_n362), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n235), .A2(new_n370), .A3(new_n331), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n322), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  NAND3_X1  g174(.A1(new_n368), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT72), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT72), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n368), .A2(new_n378), .A3(new_n372), .A4(new_n375), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n368), .A2(new_n372), .ZN(new_n382));
  INV_X1    g181(.A(new_n375), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT71), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n368), .A2(KEYINPUT30), .A3(new_n372), .A4(new_n375), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n368), .A2(new_n372), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n388), .A2(KEYINPUT71), .A3(KEYINPUT30), .A4(new_n375), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n380), .A2(new_n381), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n301), .B2(new_n302), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n329), .A3(new_n252), .ZN(new_n392));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n243), .A2(new_n290), .A3(new_n300), .A4(new_n251), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT5), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n252), .B1(new_n301), .B2(new_n302), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n394), .ZN(new_n399));
  INV_X1    g198(.A(new_n393), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n392), .A2(new_n397), .A3(new_n393), .A4(new_n395), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G1gat), .B(G29gat), .Z(new_n405));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT6), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n402), .A2(new_n409), .A3(new_n403), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n404), .A2(KEYINPUT6), .A3(new_n410), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT76), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n409), .B1(new_n402), .B2(new_n403), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT76), .B1(new_n417), .B2(KEYINPUT6), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n413), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n390), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT83), .B1(new_n360), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n279), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n269), .A2(new_n275), .A3(new_n277), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n353), .A2(new_n357), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n387), .A2(new_n389), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n377), .A2(new_n381), .A3(new_n379), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n415), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n417), .A2(KEYINPUT76), .A3(KEYINPUT6), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n430), .A2(new_n431), .B1(new_n412), .B2(new_n411), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n426), .A2(new_n433), .A3(new_n434), .A4(new_n359), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n280), .A2(new_n358), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT77), .B1(new_n429), .B2(new_n432), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT77), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n419), .A2(new_n438), .A3(new_n428), .A4(new_n427), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n421), .B(new_n435), .C1(new_n440), .C2(new_n359), .ZN(new_n441));
  INV_X1    g240(.A(new_n417), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n393), .B1(new_n392), .B2(new_n395), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT39), .B1(new_n399), .B2(new_n400), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT39), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n410), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT40), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n447), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT40), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT81), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n453), .B(KEYINPUT40), .C1(new_n445), .C2(new_n447), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n449), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT82), .B1(new_n390), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(new_n451), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n453), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n451), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n429), .A2(new_n460), .A3(new_n461), .A4(new_n449), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n383), .B1(new_n382), .B2(KEYINPUT37), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n369), .A2(new_n371), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT37), .B1(new_n464), .B2(new_n322), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n235), .A2(new_n362), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n322), .ZN(new_n467));
  INV_X1    g266(.A(new_n367), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n468), .B2(new_n370), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  OR3_X1    g269(.A1(new_n463), .A2(KEYINPUT38), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n382), .A2(KEYINPUT37), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT38), .B1(new_n472), .B2(new_n463), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n432), .A2(new_n471), .A3(new_n380), .A4(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n456), .A2(new_n462), .A3(new_n358), .A4(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n437), .A2(new_n439), .A3(new_n425), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n280), .B(KEYINPUT36), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n441), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT89), .B(G64gat), .ZN(new_n480));
  INV_X1    g279(.A(G57gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(KEYINPUT88), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n480), .B(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G71gat), .A2(G78gat), .ZN(new_n484));
  OR2_X1    g283(.A1(G71gat), .A2(G78gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT9), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G64gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n481), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n484), .B(new_n485), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT21), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G127gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(G15gat), .B(G22gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT16), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(G1gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(G1gat), .B2(new_n499), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n502), .B(G8gat), .Z(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n494), .B2(new_n493), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n498), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(new_n297), .ZN(new_n507));
  XOR2_X1   g306(.A(G183gat), .B(G211gat), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n505), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT86), .B(G36gat), .Z(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(G29gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT15), .ZN(new_n514));
  INV_X1    g313(.A(G43gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(G50gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n516), .B2(KEYINPUT87), .ZN(new_n517));
  OR3_X1    g316(.A1(KEYINPUT85), .A2(G29gat), .A3(G36gat), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(KEYINPUT14), .A3(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(KEYINPUT14), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n513), .A2(new_n517), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G43gat), .B(G50gat), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n513), .A2(new_n520), .A3(new_n521), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n514), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n522), .A2(new_n523), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT17), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n528), .A2(new_n532), .A3(new_n524), .A4(new_n526), .ZN(new_n533));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  XNOR2_X1  g334(.A(G99gat), .B(G106gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537));
  INV_X1    g336(.A(G85gat), .ZN(new_n538));
  INV_X1    g337(.A(G92gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(KEYINPUT8), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT91), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n535), .A2(new_n540), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n543), .A2(new_n536), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n530), .A2(new_n531), .A3(new_n533), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n533), .A2(new_n545), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n532), .B1(new_n527), .B2(new_n528), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT92), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n527), .A2(new_n528), .A3(new_n542), .A4(new_n544), .ZN(new_n550));
  NAND3_X1  g349(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n550), .A2(KEYINPUT93), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT93), .B1(new_n550), .B2(new_n551), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n546), .B(new_n549), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n511), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT90), .B(G134gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n298), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(new_n555), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n550), .A2(new_n551), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT93), .A3(new_n551), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n555), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n549), .A4(new_n546), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n562), .A2(new_n569), .A3(KEYINPUT94), .A4(new_n560), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n533), .A2(new_n503), .ZN(new_n575));
  OAI221_X1 g374(.A(new_n574), .B1(new_n529), .B2(new_n503), .C1(new_n575), .C2(new_n548), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT18), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n530), .A2(new_n503), .A3(new_n533), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n529), .A2(new_n503), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n579), .A2(KEYINPUT18), .A3(new_n574), .A4(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n529), .B(new_n503), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n574), .B(KEYINPUT13), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n578), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT12), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n581), .A3(new_n584), .A4(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n493), .B1(new_n542), .B2(KEYINPUT95), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n545), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n542), .B(new_n544), .C1(new_n493), .C2(KEYINPUT95), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT10), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n545), .A2(new_n602), .A3(new_n493), .ZN(new_n603));
  INV_X1    g402(.A(G230gat), .ZN(new_n604));
  OAI22_X1  g403(.A1(new_n601), .A2(new_n603), .B1(new_n604), .B2(new_n256), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n256), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n599), .A2(new_n606), .A3(new_n600), .ZN(new_n607));
  XOR2_X1   g406(.A(G120gat), .B(G148gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT96), .ZN(new_n609));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n605), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n605), .B2(new_n607), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n597), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n605), .A2(new_n607), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n611), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n605), .A2(new_n607), .A3(new_n612), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(KEYINPUT97), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NOR4_X1   g419(.A1(new_n510), .A2(new_n573), .A3(new_n596), .A4(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n479), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n432), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT98), .B(G1gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(G1324gat));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n626));
  INV_X1    g425(.A(new_n622), .ZN(new_n627));
  OAI21_X1  g426(.A(G8gat), .B1(new_n627), .B2(new_n390), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT16), .B(G8gat), .Z(new_n629));
  NAND3_X1  g428(.A1(new_n622), .A2(new_n429), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n626), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n626), .B2(new_n630), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT99), .Z(G1325gat));
  OR3_X1    g432(.A1(new_n627), .A2(G15gat), .A3(new_n424), .ZN(new_n634));
  OAI21_X1  g433(.A(G15gat), .B1(new_n627), .B2(new_n477), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(G1326gat));
  NAND2_X1  g435(.A1(new_n622), .A2(new_n425), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT100), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT43), .B(G22gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(G1327gat));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n479), .A2(new_n641), .A3(new_n573), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n572), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n556), .A2(new_n560), .B1(new_n562), .B2(new_n569), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n441), .B2(new_n478), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n641), .A3(KEYINPUT44), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n510), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n651), .A2(new_n596), .A3(new_n620), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G29gat), .B1(new_n653), .B2(new_n419), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n648), .A2(new_n652), .ZN(new_n655));
  INV_X1    g454(.A(G29gat), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n656), .A3(new_n432), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT45), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(G1328gat));
  NOR2_X1   g458(.A1(new_n390), .A2(new_n512), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT102), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(KEYINPUT46), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n662), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(KEYINPUT46), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n512), .B1(new_n653), .B2(new_n390), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(G1329gat));
  NAND3_X1  g467(.A1(new_n655), .A2(new_n515), .A3(new_n280), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT104), .ZN(new_n670));
  INV_X1    g469(.A(new_n477), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n650), .A2(new_n671), .A3(new_n652), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n670), .B1(new_n673), .B2(new_n515), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g474(.A(G50gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n650), .A2(new_n425), .A3(new_n652), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(KEYINPUT106), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(KEYINPUT106), .B2(new_n677), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n655), .A2(new_n676), .A3(new_n425), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(KEYINPUT48), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(G50gat), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT48), .B1(new_n682), .B2(new_n680), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(G1331gat));
  NOR2_X1   g486(.A1(new_n510), .A2(new_n573), .ZN(new_n688));
  INV_X1    g487(.A(new_n620), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n595), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n479), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT107), .Z(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n432), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G57gat), .ZN(G1332gat));
  INV_X1    g493(.A(KEYINPUT49), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n692), .B(new_n429), .C1(new_n695), .C2(new_n489), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n698), .A2(new_n699), .B1(new_n695), .B2(new_n489), .ZN(new_n700));
  INV_X1    g499(.A(new_n699), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(new_n489), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n700), .A2(new_n703), .ZN(G1333gat));
  XNOR2_X1  g503(.A(new_n280), .B(KEYINPUT109), .ZN(new_n705));
  AOI21_X1  g504(.A(G71gat), .B1(new_n692), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n671), .A2(G71gat), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n692), .B2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n425), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n651), .A2(new_n595), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n479), .A2(new_n573), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n648), .A2(KEYINPUT51), .A3(new_n712), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n689), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n538), .A3(new_n432), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n651), .A2(new_n595), .A3(new_n689), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n650), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G85gat), .B1(new_n722), .B2(new_n419), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(G1336gat));
  NOR2_X1   g523(.A1(new_n390), .A2(G92gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n644), .A2(new_n429), .A3(new_n649), .A4(new_n721), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G92gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n731), .A3(new_n716), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n713), .A2(KEYINPUT110), .A3(new_n714), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n725), .A2(new_n620), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n729), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT111), .B1(new_n736), .B2(KEYINPUT52), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738));
  AOI211_X1 g537(.A(new_n738), .B(new_n727), .C1(new_n735), .C2(new_n729), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n730), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g541(.A(KEYINPUT112), .B(new_n730), .C1(new_n737), .C2(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1337gat));
  XOR2_X1   g543(.A(KEYINPUT113), .B(G99gat), .Z(new_n745));
  NAND3_X1  g544(.A1(new_n719), .A2(new_n280), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n722), .A2(new_n477), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(new_n745), .ZN(G1338gat));
  OAI21_X1  g547(.A(G106gat), .B1(new_n722), .B2(new_n358), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n689), .A2(G106gat), .A3(new_n358), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT114), .Z(new_n751));
  NAND3_X1  g550(.A1(new_n732), .A2(new_n733), .A3(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754));
  INV_X1    g553(.A(new_n749), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n718), .B2(new_n750), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(G1339gat));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n599), .A2(new_n600), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n602), .ZN(new_n760));
  INV_X1    g559(.A(new_n603), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n606), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n762), .A2(new_n605), .A3(KEYINPUT54), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  OAI221_X1 g563(.A(new_n764), .B1(new_n604), .B2(new_n256), .C1(new_n601), .C2(new_n603), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n611), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n758), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n582), .A2(new_n583), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n574), .B1(new_n579), .B2(new_n580), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n590), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n594), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n762), .A2(new_n605), .A3(KEYINPUT54), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(KEYINPUT55), .A3(new_n611), .A4(new_n765), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n767), .A2(new_n771), .A3(new_n618), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT115), .B1(new_n774), .B2(new_n647), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n594), .A2(new_n770), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n772), .A2(new_n611), .A3(new_n765), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n758), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n773), .A2(new_n618), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n573), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n777), .A2(new_n758), .B1(new_n593), .B2(new_n594), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n782), .A2(new_n779), .B1(new_n620), .B2(new_n771), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n775), .B(new_n781), .C1(new_n783), .C2(new_n573), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n510), .ZN(new_n785));
  NOR4_X1   g584(.A1(new_n510), .A2(new_n573), .A3(new_n595), .A4(new_n620), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n432), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n436), .A2(new_n429), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(G113gat), .B1(new_n793), .B2(new_n595), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n788), .A2(KEYINPUT116), .A3(new_n358), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n786), .B1(new_n784), .B2(new_n510), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n425), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n429), .A2(new_n419), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n280), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n596), .A2(new_n244), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n794), .B1(new_n802), .B2(new_n803), .ZN(G1340gat));
  NOR4_X1   g603(.A1(new_n792), .A2(new_n237), .A3(new_n236), .A4(new_n689), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n620), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(G120gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT117), .ZN(G1341gat));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n247), .A3(new_n651), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n799), .A2(new_n510), .A3(new_n801), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n247), .ZN(G1342gat));
  NOR3_X1   g610(.A1(new_n792), .A2(G134gat), .A3(new_n647), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT56), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n799), .A2(new_n647), .A3(new_n801), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n249), .B2(new_n814), .ZN(G1343gat));
  AND2_X1   g614(.A1(new_n477), .A2(new_n800), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n425), .A2(KEYINPUT57), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n786), .B1(new_n785), .B2(KEYINPUT118), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n784), .A2(new_n819), .A3(new_n510), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n817), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT57), .B1(new_n788), .B2(new_n425), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n595), .B(new_n816), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G141gat), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n477), .A2(new_n425), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n390), .ZN(new_n827));
  NOR4_X1   g626(.A1(new_n789), .A2(G141gat), .A3(new_n596), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT120), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n823), .B2(G141gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n824), .A2(new_n836), .A3(new_n829), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n831), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n824), .B2(new_n829), .ZN(new_n839));
  AOI211_X1 g638(.A(KEYINPUT120), .B(new_n828), .C1(new_n823), .C2(G141gat), .ZN(new_n840));
  OAI22_X1  g639(.A1(new_n839), .A2(new_n840), .B1(new_n834), .B2(new_n833), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n838), .A2(new_n841), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n783), .A2(new_n573), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n774), .A2(new_n647), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n510), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n787), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n846), .B2(new_n425), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n797), .A2(new_n817), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n816), .A2(new_n620), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT59), .B(G148gat), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n689), .A2(KEYINPUT59), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n789), .A2(new_n827), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n620), .ZN(new_n856));
  OAI221_X1 g655(.A(new_n851), .B1(new_n852), .B2(new_n853), .C1(G148gat), .C2(new_n856), .ZN(G1345gat));
  INV_X1    g656(.A(new_n855), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n858), .A2(KEYINPUT121), .A3(new_n510), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT121), .B1(new_n858), .B2(new_n510), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n297), .A3(new_n860), .ZN(new_n861));
  OR3_X1    g660(.A1(new_n852), .A2(new_n297), .A3(new_n510), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(G1346gat));
  OAI21_X1  g662(.A(new_n298), .B1(new_n858), .B2(new_n647), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n573), .A2(G162gat), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n852), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g666(.A1(new_n797), .A2(new_n432), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n429), .A3(new_n426), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(G169gat), .B1(new_n870), .B2(new_n595), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n705), .A2(new_n419), .A3(new_n429), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT123), .Z(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n795), .B2(new_n798), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n596), .A2(new_n206), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(G1348gat));
  NAND3_X1  g675(.A1(new_n870), .A2(new_n207), .A3(new_n620), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n874), .A2(new_n620), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n207), .ZN(G1349gat));
  AOI21_X1  g678(.A(new_n215), .B1(new_n874), .B2(new_n651), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n651), .A2(new_n222), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n870), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT60), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n882), .B(new_n884), .ZN(G1350gat));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n874), .A2(new_n573), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(G190gat), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT125), .B(new_n219), .C1(new_n874), .C2(new_n573), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT126), .B(new_n886), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n870), .A2(new_n219), .A3(new_n573), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT126), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT61), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT126), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n891), .B(new_n892), .C1(new_n894), .C2(new_n895), .ZN(G1351gat));
  NOR2_X1   g695(.A1(new_n825), .A2(new_n390), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n868), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(G197gat), .B1(new_n899), .B2(new_n595), .ZN(new_n900));
  NOR4_X1   g699(.A1(new_n849), .A2(new_n432), .A3(new_n390), .A4(new_n671), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n595), .A2(G197gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(G1352gat));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n620), .ZN(new_n904));
  XOR2_X1   g703(.A(KEYINPUT127), .B(G204gat), .Z(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n898), .A2(new_n689), .A3(new_n905), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT62), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1353gat));
  OR3_X1    g708(.A1(new_n898), .A2(G211gat), .A3(new_n510), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n901), .A2(new_n651), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n911), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT63), .B1(new_n911), .B2(G211gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1354gat));
  INV_X1    g713(.A(G218gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n915), .A3(new_n573), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n901), .A2(new_n573), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n915), .ZN(G1355gat));
endmodule


