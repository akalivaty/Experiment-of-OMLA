//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n527,
    new_n528, new_n531, new_n532, new_n533, new_n534, new_n535, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1116, new_n1117, new_n1118;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT66), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  INV_X1    g052(.A(new_n474), .ZN(new_n478));
  OR2_X1    g053(.A1(new_n478), .A2(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(KEYINPUT67), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT68), .Z(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n460), .B1(new_n466), .B2(new_n468), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT69), .Z(new_n488));
  AND3_X1   g063(.A1(new_n483), .A2(new_n485), .A3(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(G114), .B2(new_n460), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n463), .A2(new_n469), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT70), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n502), .B(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n503), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(new_n501), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(G166));
  INV_X1    g090(.A(new_n508), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G89), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n503), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G51), .ZN(new_n519));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n507), .A2(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n517), .A2(new_n519), .A3(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  AOI22_X1  g101(.A1(new_n516), .A2(G90), .B1(new_n518), .B2(G52), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n501), .B2(new_n528), .ZN(G301));
  INV_X1    g104(.A(G301), .ZN(G171));
  NAND2_X1  g105(.A1(new_n516), .A2(G81), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT72), .B(G43), .ZN(new_n533));
  OAI221_X1 g108(.A(new_n531), .B1(new_n501), .B2(new_n532), .C1(new_n510), .C2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND4_X1  g114(.A1(G319), .A2(G483), .A3(G661), .A4(new_n539), .ZN(G188));
  NAND2_X1  g115(.A1(new_n518), .A2(G53), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT9), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n503), .A2(new_n544), .A3(new_n507), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G91), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n542), .B(new_n547), .C1(new_n501), .C2(new_n548), .ZN(G299));
  INV_X1    g124(.A(G166), .ZN(G303));
  NAND3_X1  g125(.A1(new_n543), .A2(G87), .A3(new_n545), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n505), .A2(new_n506), .ZN(new_n552));
  AOI21_X1  g127(.A(KEYINPUT5), .B1(new_n504), .B2(G543), .ZN(new_n553));
  OR3_X1    g128(.A1(new_n552), .A2(G74), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n518), .A2(G49), .B1(G651), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G288));
  NOR2_X1   g131(.A1(new_n552), .A2(new_n553), .ZN(new_n557));
  INV_X1    g132(.A(G61), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT74), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G73), .ZN(new_n560));
  INV_X1    g135(.A(G543), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR3_X1   g137(.A1(new_n557), .A2(KEYINPUT74), .A3(new_n558), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n518), .A2(G48), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n546), .A2(G86), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(G305));
  INV_X1    g143(.A(G85), .ZN(new_n569));
  INV_X1    g144(.A(G47), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n508), .A2(new_n569), .B1(new_n510), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n501), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n546), .A2(G92), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT10), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n577), .B(KEYINPUT75), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n518), .A2(KEYINPUT76), .ZN(new_n584));
  INV_X1    g159(.A(G54), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n585), .B1(new_n510), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G79), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT77), .B1(new_n588), .B2(new_n561), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n588), .A2(new_n561), .A3(KEYINPUT77), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n557), .C2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n584), .A2(new_n587), .B1(G651), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n580), .A2(new_n583), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n576), .B1(new_n595), .B2(G868), .ZN(G321));
  XNOR2_X1  g171(.A(G321), .B(KEYINPUT78), .ZN(G284));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G299), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(G168), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(new_n598), .B2(G168), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n535), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g182(.A1(new_n463), .A2(new_n469), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n608), .A2(G2104), .A3(new_n460), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT13), .Z(new_n612));
  INV_X1    g187(.A(G2100), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n481), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n486), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n460), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND3_X1  g196(.A1(new_n614), .A2(new_n615), .A3(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(G2427), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n628), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G14), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n632), .A2(new_n635), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  INV_X1    g222(.A(new_n640), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n647), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1956), .B(G2474), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n657), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT20), .Z(new_n661));
  AOI211_X1 g236(.A(new_n659), .B(new_n661), .C1(new_n654), .C2(new_n658), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1991), .B(G1996), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT82), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G229));
  INV_X1    g244(.A(G16), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G22), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(G166), .B2(new_n670), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1971), .ZN(new_n673));
  NOR2_X1   g248(.A1(G16), .A2(G23), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT85), .ZN(new_n675));
  AND3_X1   g250(.A1(new_n551), .A2(new_n555), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n675), .B1(new_n551), .B2(new_n555), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n674), .B1(new_n678), .B2(G16), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT33), .B(G1976), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g256(.A(G6), .B(G305), .S(G16), .Z(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT32), .B(G1981), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI211_X1 g261(.A(new_n673), .B(new_n686), .C1(new_n682), .C2(new_n683), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT86), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n670), .A2(G24), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n574), .B2(new_n670), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT84), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1986), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G25), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n481), .A2(G131), .ZN(new_n698));
  OAI21_X1  g273(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n699));
  INV_X1    g274(.A(G107), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G2105), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n486), .B2(G119), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n697), .B1(new_n704), .B2(new_n696), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT35), .B(G1991), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT83), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n695), .A2(KEYINPUT87), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n690), .A2(new_n691), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n481), .A2(G141), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n486), .A2(G129), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT26), .Z(new_n717));
  NAND3_X1  g292(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n714), .A2(new_n715), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G32), .B(new_n719), .S(G29), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT27), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1996), .ZN(new_n722));
  NOR2_X1   g297(.A1(G171), .A2(new_n670), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G5), .B2(new_n670), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT93), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n696), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n696), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G2090), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n722), .B(new_n727), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n595), .A2(new_n670), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G4), .B2(new_n670), .ZN(new_n734));
  INV_X1    g309(.A(G1348), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n620), .A2(new_n696), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT92), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(KEYINPUT92), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  INV_X1    g316(.A(G28), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n742), .B2(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n739), .A2(new_n740), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G19), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n535), .B2(G16), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n724), .A2(new_n725), .B1(G1341), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(G1341), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n696), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n696), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n746), .A2(new_n749), .A3(new_n750), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n696), .A2(G33), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n608), .A2(G127), .ZN(new_n757));
  NAND2_X1  g332(.A1(G115), .A2(G2104), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n460), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT89), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  AOI211_X1 g337(.A(new_n759), .B(new_n762), .C1(G139), .C2(new_n481), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n756), .B1(new_n763), .B2(new_n696), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2072), .ZN(new_n765));
  INV_X1    g340(.A(G34), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(KEYINPUT24), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n696), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G160), .B2(new_n696), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2084), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n755), .A2(new_n765), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n734), .A2(new_n735), .ZN(new_n773));
  NAND2_X1  g348(.A1(G299), .A2(G16), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n670), .A2(G20), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT23), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT90), .B1(G16), .B2(G21), .ZN(new_n779));
  NAND2_X1  g354(.A1(G168), .A2(G16), .ZN(new_n780));
  MUX2_X1   g355(.A(KEYINPUT90), .B(new_n779), .S(new_n780), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT91), .B(G1966), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n696), .A2(G26), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT28), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n481), .A2(G140), .ZN(new_n787));
  NOR2_X1   g362(.A1(G104), .A2(G2105), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT88), .ZN(new_n789));
  INV_X1    g364(.A(G116), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n465), .B1(new_n790), .B2(G2105), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n789), .A2(new_n791), .B1(G128), .B2(new_n486), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n786), .B1(new_n793), .B2(G29), .ZN(new_n794));
  INV_X1    g369(.A(G2067), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n778), .A2(new_n783), .A3(new_n784), .A4(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n736), .A2(new_n772), .A3(new_n773), .A4(new_n797), .ZN(new_n798));
  AOI211_X1 g373(.A(new_n732), .B(new_n798), .C1(new_n731), .C2(new_n730), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n712), .A2(new_n713), .A3(new_n799), .ZN(G150));
  INV_X1    g375(.A(G150), .ZN(G311));
  NAND2_X1  g376(.A1(new_n595), .A2(G559), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT38), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n516), .A2(G93), .B1(new_n518), .B2(G55), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n501), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n534), .B(new_n806), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n803), .B(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n809), .A2(new_n810), .A3(G860), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n806), .A2(G860), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n811), .A2(new_n813), .ZN(G145));
  INV_X1    g389(.A(KEYINPUT97), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n763), .B2(KEYINPUT96), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n815), .B2(new_n763), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n719), .B(new_n793), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n499), .A2(new_n496), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n820));
  INV_X1    g395(.A(G114), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n490), .B1(new_n821), .B2(G2105), .ZN(new_n822));
  NAND2_X1  g397(.A1(G126), .A2(G2105), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n466), .B2(new_n468), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT95), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n819), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n818), .B(new_n827), .ZN(new_n828));
  MUX2_X1   g403(.A(new_n817), .B(new_n816), .S(new_n828), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n703), .B(KEYINPUT99), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n486), .A2(G130), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT98), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G118), .B2(new_n460), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n832), .A2(KEYINPUT98), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n481), .B2(G142), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n830), .B(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(new_n611), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n829), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n620), .B(G160), .ZN(new_n841));
  XNOR2_X1  g416(.A(G162), .B(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(G37), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n840), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT100), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g421(.A1(new_n806), .A2(new_n598), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n678), .B(new_n574), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(G305), .B(G303), .ZN(new_n850));
  OR3_X1    g425(.A1(new_n849), .A2(KEYINPUT102), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n849), .A2(KEYINPUT102), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT42), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n594), .B(G299), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(KEYINPUT41), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n595), .A2(G299), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT101), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n857), .B2(KEYINPUT101), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n859), .B1(new_n862), .B2(KEYINPUT41), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n604), .B(new_n807), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n862), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n856), .B1(new_n867), .B2(KEYINPUT103), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(KEYINPUT103), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n868), .B(new_n869), .Z(new_n870));
  OAI21_X1  g445(.A(new_n847), .B1(new_n870), .B2(new_n598), .ZN(G295));
  OAI21_X1  g446(.A(new_n847), .B1(new_n870), .B2(new_n598), .ZN(G331));
  XNOR2_X1  g447(.A(new_n807), .B(G301), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G168), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n866), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n863), .B2(new_n875), .ZN(new_n877));
  INV_X1    g452(.A(new_n855), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n880), .B2(new_n858), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n862), .B2(new_n880), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT104), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(new_n885), .A3(new_n882), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(KEYINPUT43), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n876), .B(new_n855), .C1(new_n863), .C2(new_n875), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n879), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n890), .A2(KEYINPUT44), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n887), .A2(KEYINPUT105), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT105), .B1(new_n887), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n883), .A2(KEYINPUT43), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n888), .B1(new_n879), .B2(new_n889), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI22_X1  g471(.A1(new_n892), .A2(new_n893), .B1(KEYINPUT44), .B2(new_n896), .ZN(G397));
  INV_X1    g472(.A(G1384), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n827), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G40), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n472), .A2(new_n900), .A3(new_n476), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(KEYINPUT106), .Z(new_n904));
  INV_X1    g479(.A(G1996), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n719), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n793), .B(new_n795), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n703), .B(new_n706), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(KEYINPUT108), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(KEYINPUT108), .B2(new_n910), .ZN(new_n912));
  INV_X1    g487(.A(G1986), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n574), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT107), .Z(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n913), .B2(new_n574), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n904), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT49), .ZN(new_n919));
  INV_X1    g494(.A(G1981), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n516), .A2(G86), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n566), .B2(new_n921), .ZN(new_n922));
  AND4_X1   g497(.A1(new_n920), .A2(new_n567), .A3(new_n565), .A4(new_n564), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n566), .A2(new_n920), .A3(new_n567), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n564), .A2(new_n565), .ZN(new_n926));
  INV_X1    g501(.A(new_n921), .ZN(new_n927));
  OAI21_X1  g502(.A(G1981), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(KEYINPUT49), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n899), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n930), .A2(new_n901), .ZN(new_n931));
  INV_X1    g506(.A(G8), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n924), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(G288), .A2(KEYINPUT85), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n551), .A2(new_n555), .A3(new_n675), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(G1976), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(new_n937), .B2(KEYINPUT113), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT113), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n678), .B2(G1976), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT52), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n678), .A2(new_n939), .A3(G1976), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(KEYINPUT113), .ZN(new_n943));
  INV_X1    g518(.A(G1976), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT52), .B1(G288), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n933), .A4(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n934), .A2(new_n941), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n902), .A2(G1384), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n827), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n827), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n902), .B1(G164), .B2(G1384), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n901), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n948), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1971), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n827), .A2(new_n950), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT109), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n827), .A2(new_n949), .A3(new_n950), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n954), .A2(new_n901), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT110), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n956), .A2(new_n957), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n819), .A2(new_n493), .A3(new_n492), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n898), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n901), .C1(KEYINPUT50), .C2(new_n899), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(G2090), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(G166), .A2(new_n932), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n971), .B1(new_n974), .B2(KEYINPUT55), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(G8), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n932), .B1(new_n964), .B2(new_n969), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(KEYINPUT112), .A3(new_n976), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n947), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n899), .A2(KEYINPUT50), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n983), .B(new_n901), .C1(KEYINPUT50), .C2(new_n966), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(G2090), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n964), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G8), .ZN(new_n987));
  INV_X1    g562(.A(new_n976), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(KEYINPUT114), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n932), .B1(new_n964), .B2(new_n985), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(new_n976), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n982), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT126), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n968), .A2(new_n725), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n966), .A2(new_n902), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n899), .A2(new_n902), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n998), .A2(KEYINPUT53), .A3(new_n753), .A4(new_n901), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n1000), .B(KEYINPUT124), .Z(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT125), .B(KEYINPUT53), .Z(new_n1002));
  NAND2_X1  g577(.A1(new_n956), .A2(new_n963), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n753), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G171), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(new_n901), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G164), .A2(G1384), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1007), .B1(KEYINPUT45), .B2(new_n1008), .ZN(new_n1009));
  OAI22_X1  g584(.A1(new_n1009), .A2(G1966), .B1(G2084), .B2(new_n968), .ZN(new_n1010));
  OAI21_X1  g585(.A(G8), .B1(new_n1010), .B2(G286), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(KEYINPUT51), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1010), .A2(G286), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n1013), .B2(new_n1011), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1006), .B1(new_n1015), .B2(KEYINPUT62), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n995), .B(new_n1016), .C1(KEYINPUT62), .C2(new_n1015), .ZN(new_n1017));
  XNOR2_X1  g592(.A(G299), .B(KEYINPUT57), .ZN(new_n1018));
  INV_X1    g593(.A(G1956), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n984), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n961), .A2(new_n962), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(G2072), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1020), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1027));
  OR3_X1    g602(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT121), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1026), .B2(KEYINPUT121), .ZN(new_n1029));
  NAND2_X1  g604(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT61), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n968), .A2(new_n735), .B1(new_n931), .B2(new_n795), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n594), .B1(KEYINPUT60), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT123), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n594), .A2(KEYINPUT60), .A3(new_n1034), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT122), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n1035), .A2(new_n1036), .B1(new_n1038), .B2(KEYINPUT122), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n1040), .A2(new_n1041), .B1(KEYINPUT60), .B2(new_n1034), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT58), .B(G1341), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n1021), .A2(G1996), .B1(new_n931), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n535), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT59), .Z(new_n1046));
  INV_X1    g621(.A(new_n1031), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(KEYINPUT120), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1033), .A2(new_n1042), .A3(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1027), .A2(new_n594), .A3(new_n1034), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(new_n1026), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n996), .B1(new_n999), .B2(new_n953), .ZN(new_n1053));
  OR3_X1    g628(.A1(new_n1004), .A2(G171), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT54), .B1(new_n1006), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1005), .A2(G171), .ZN(new_n1056));
  OAI21_X1  g631(.A(G171), .B1(new_n1004), .B2(new_n1053), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT54), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1015), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1055), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1052), .A2(new_n1061), .A3(new_n995), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n979), .A2(new_n981), .ZN(new_n1065));
  INV_X1    g640(.A(new_n947), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1010), .A2(G8), .A3(G168), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1010), .A2(KEYINPUT115), .A3(G8), .A4(G168), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1065), .A2(new_n993), .A3(new_n1066), .A4(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1072), .A2(KEYINPUT116), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n982), .A2(new_n1074), .A3(new_n993), .A4(new_n1071), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT63), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1064), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1072), .A2(KEYINPUT116), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(KEYINPUT117), .A3(new_n1076), .A4(new_n1075), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n980), .A2(new_n976), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n982), .A2(KEYINPUT63), .A3(new_n1071), .A4(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1065), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n934), .A2(new_n944), .A3(new_n551), .A4(new_n555), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n925), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1084), .A2(new_n1066), .B1(new_n933), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT118), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1083), .A2(new_n1090), .A3(new_n1087), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1063), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1017), .B1(new_n1092), .B2(KEYINPUT127), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1091), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1090), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1095));
  OAI211_X1 g670(.A(KEYINPUT127), .B(new_n1062), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n918), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n904), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n916), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(KEYINPUT48), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1100), .A2(KEYINPUT48), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n1101), .B(new_n1102), .C1(new_n904), .C2(new_n912), .ZN(new_n1103));
  INV_X1    g678(.A(new_n907), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n904), .B1(new_n1104), .B2(new_n719), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1099), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT46), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n904), .B2(new_n905), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1105), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(new_n1109), .B(KEYINPUT47), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n704), .A2(new_n706), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n908), .A2(new_n1111), .B1(G2067), .B2(new_n793), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n1103), .B(new_n1110), .C1(new_n904), .C2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1098), .A2(new_n1113), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g689(.A(G227), .ZN(new_n1116));
  NAND2_X1  g690(.A1(new_n1116), .A2(G319), .ZN(new_n1117));
  OR3_X1    g691(.A1(G229), .A2(G401), .A3(new_n1117), .ZN(new_n1118));
  NOR3_X1   g692(.A1(new_n896), .A2(new_n845), .A3(new_n1118), .ZN(G308));
  INV_X1    g693(.A(G308), .ZN(G225));
endmodule


