//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n576, new_n577, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT64), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G101), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT68), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n464), .A2(new_n466), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT67), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n464), .A2(new_n466), .A3(new_n479), .A4(G125), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n474), .A2(new_n482), .ZN(G160));
  XNOR2_X1  g058(.A(new_n466), .B(new_n467), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT69), .A3(new_n464), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n470), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n487), .A3(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n485), .A2(new_n487), .A3(KEYINPUT70), .A4(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n485), .A2(new_n487), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(new_n473), .ZN(new_n495));
  INV_X1    g070(.A(G136), .ZN(new_n496));
  NOR2_X1   g071(.A1(G100), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(new_n473), .B2(G112), .ZN(new_n498));
  OAI22_X1  g073(.A1(new_n495), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n493), .A2(new_n499), .ZN(G162));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n473), .A2(G138), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n484), .A2(new_n464), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n503), .B1(new_n475), .B2(new_n502), .ZN(new_n506));
  OR3_X1    g081(.A1(new_n473), .A2(KEYINPUT71), .A3(G114), .ZN(new_n507));
  OR2_X1    g082(.A1(G102), .A2(G2105), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT71), .B1(new_n473), .B2(G114), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n507), .A2(G2104), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n505), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n505), .A2(KEYINPUT72), .A3(new_n506), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(G164));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n517), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT5), .B(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT73), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  NAND2_X1  g104(.A1(G75), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(new_n526), .ZN(new_n531));
  INV_X1    g106(.A(G62), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n525), .A2(G543), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n533), .A2(G651), .B1(new_n534), .B2(G50), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n529), .A2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  NAND3_X1  g112(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n534), .A2(G51), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT74), .B(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n524), .A2(new_n527), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n542), .B1(new_n541), .B2(new_n544), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n538), .B(new_n539), .C1(new_n545), .C2(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  XNOR2_X1  g123(.A(KEYINPUT77), .B(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n528), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  INV_X1    g126(.A(new_n534), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G64), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n531), .B2(new_n554), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n555), .A2(KEYINPUT76), .A3(G651), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT76), .B1(new_n555), .B2(G651), .ZN(new_n557));
  OAI221_X1 g132(.A(new_n550), .B1(new_n551), .B2(new_n552), .C1(new_n556), .C2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  AOI22_X1  g134(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G651), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n524), .A2(G81), .A3(new_n527), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n534), .A2(G43), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(KEYINPUT78), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT79), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n569), .B(new_n562), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  AND3_X1   g147(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G36), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT80), .Z(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G188));
  NAND2_X1  g153(.A1(new_n534), .A2(G53), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n528), .A2(G91), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n526), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n561), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(G299));
  OAI21_X1  g159(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n534), .A2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n524), .A2(new_n527), .ZN(new_n587));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n528), .A2(G86), .B1(G48), .B2(new_n534), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n531), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(KEYINPUT81), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n593), .B2(G651), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n595), .B2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n528), .A2(G85), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n531), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n534), .B2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G290));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n531), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(new_n534), .B2(G54), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT10), .B1(new_n587), .B2(new_n605), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G171), .B2(new_n613), .ZN(G284));
  OAI21_X1  g190(.A(new_n614), .B1(G171), .B2(new_n613), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT82), .Z(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(G868), .B2(new_n619), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(G868), .B2(new_n619), .ZN(G280));
  AND3_X1   g196(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n571), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g204(.A(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(new_n473), .B2(G111), .ZN(new_n632));
  OAI22_X1  g207(.A1(new_n495), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(G123), .B2(new_n492), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n473), .A2(G2104), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n475), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT85), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(G2100), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT85), .B(G2100), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n635), .B(new_n642), .C1(new_n643), .C2(new_n640), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT86), .Z(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2435), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2443), .B(G2446), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G14), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT87), .Z(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT17), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT89), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n676), .A2(new_n679), .A3(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT91), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G25), .ZN(new_n694));
  OAI21_X1  g269(.A(KEYINPUT92), .B1(new_n694), .B2(G29), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n694), .A2(KEYINPUT92), .A3(G29), .ZN(new_n696));
  INV_X1    g271(.A(G107), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n465), .B1(new_n697), .B2(G2105), .ZN(new_n698));
  OR2_X1    g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G131), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n495), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G119), .B2(new_n492), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n695), .B(new_n696), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT35), .B(G1991), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT93), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n705), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G6), .ZN(new_n711));
  INV_X1    g286(.A(G305), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n710), .A2(G22), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G303), .B2(G16), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1971), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n714), .B(new_n711), .C1(new_n712), .C2(new_n710), .ZN(new_n720));
  OAI21_X1  g295(.A(KEYINPUT94), .B1(G16), .B2(G23), .ZN(new_n721));
  OR3_X1    g296(.A1(KEYINPUT94), .A2(G16), .A3(G23), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n721), .B(new_n722), .C1(G288), .C2(new_n710), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT33), .B(G1976), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT95), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n716), .A2(new_n719), .A3(new_n720), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT96), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n727), .A2(new_n728), .A3(KEYINPUT34), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n728), .B1(new_n727), .B2(KEYINPUT34), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n709), .B1(KEYINPUT34), .B2(new_n727), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G24), .B(G290), .S(G16), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1986), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT97), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n732), .A2(KEYINPUT97), .A3(new_n734), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g313(.A(KEYINPUT97), .B(KEYINPUT36), .C1(new_n732), .C2(new_n734), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G16), .A2(G21), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G168), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT99), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G29), .B2(G33), .ZN(new_n746));
  OR3_X1    g321(.A1(new_n745), .A2(G29), .A3(G33), .ZN(new_n747));
  NAND2_X1  g322(.A1(G115), .A2(G2104), .ZN(new_n748));
  INV_X1    g323(.A(G127), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n475), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2105), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT100), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n485), .A2(new_n487), .A3(G139), .A4(new_n473), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT101), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n753), .A2(KEYINPUT101), .A3(new_n754), .A4(new_n756), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n746), .B(new_n747), .C1(new_n761), .C2(new_n704), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2072), .ZN(new_n763));
  OR2_X1    g338(.A1(G29), .A2(G32), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n485), .A2(new_n487), .A3(G141), .A4(new_n473), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT103), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT105), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT26), .ZN(new_n772));
  INV_X1    g347(.A(G105), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n636), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n492), .A2(KEYINPUT104), .A3(G129), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(KEYINPUT104), .B1(new_n492), .B2(G129), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n764), .B1(new_n779), .B2(new_n704), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT27), .B(G1996), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT106), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(KEYINPUT24), .A2(G34), .ZN(new_n784));
  NAND2_X1  g359(.A1(KEYINPUT24), .A2(G34), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n784), .A2(new_n704), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G160), .B2(new_n704), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT102), .ZN(new_n788));
  INV_X1    g363(.A(G2084), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n763), .A2(new_n783), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT107), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n763), .A2(new_n793), .A3(new_n783), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n780), .A2(new_n782), .ZN(new_n796));
  OAI21_X1  g371(.A(G29), .B1(new_n493), .B2(new_n499), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT29), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n704), .A2(G35), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n798), .B1(new_n797), .B2(new_n799), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n800), .A2(new_n801), .A3(G2090), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n710), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n571), .B2(new_n710), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n796), .B(new_n802), .C1(G1341), .C2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT31), .B(G11), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT30), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n807), .A2(G28), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(G28), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n808), .A2(new_n809), .A3(G29), .ZN(new_n810));
  NOR2_X1   g385(.A1(G164), .A2(new_n704), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G27), .B2(new_n704), .ZN(new_n812));
  INV_X1    g387(.A(G2078), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G4), .A2(G16), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n622), .B2(G16), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(G1348), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G29), .B2(new_n634), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT108), .B1(G5), .B2(G16), .ZN(new_n819));
  OR3_X1    g394(.A1(KEYINPUT108), .A2(G5), .A3(G16), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n819), .B(new_n820), .C1(G301), .C2(new_n710), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1961), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n816), .A2(G1348), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n814), .A2(new_n818), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n704), .A2(G26), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT98), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT28), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n494), .A2(G140), .A3(new_n473), .ZN(new_n828));
  OR2_X1    g403(.A1(G104), .A2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G128), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n490), .B2(new_n491), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n827), .B1(new_n834), .B2(new_n704), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2067), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n788), .A2(new_n789), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n813), .B2(new_n812), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n824), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n795), .A2(new_n805), .A3(new_n806), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(G2090), .B1(new_n800), .B2(new_n801), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT109), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n710), .A2(KEYINPUT23), .A3(G20), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT23), .ZN(new_n845));
  INV_X1    g420(.A(G20), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(G16), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n844), .B(new_n847), .C1(new_n619), .C2(new_n710), .ZN(new_n848));
  INV_X1    g423(.A(G1956), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OAI211_X1 g425(.A(KEYINPUT109), .B(G2090), .C1(new_n800), .C2(new_n801), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n843), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT110), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT110), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n843), .A2(new_n854), .A3(new_n850), .A4(new_n851), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n804), .A2(G1341), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n840), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n740), .A2(new_n744), .A3(new_n858), .ZN(G311));
  NAND3_X1  g434(.A1(new_n740), .A2(new_n744), .A3(new_n858), .ZN(G150));
  INV_X1    g435(.A(G55), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n552), .A2(new_n861), .B1(new_n561), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G93), .B2(new_n528), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G860), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT37), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n563), .A2(new_n564), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT78), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n564), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n569), .B1(new_n872), .B2(new_n562), .ZN(new_n873));
  INV_X1    g448(.A(new_n570), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n865), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT111), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n567), .A2(new_n864), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT111), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n571), .A2(new_n878), .A3(new_n865), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n612), .A2(new_n623), .ZN(new_n881));
  XOR2_X1   g456(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n880), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n867), .B1(new_n884), .B2(G860), .ZN(G145));
  XNOR2_X1  g460(.A(new_n634), .B(G160), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G162), .ZN(new_n887));
  INV_X1    g462(.A(new_n639), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n703), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n492), .A2(G119), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n639), .B1(new_n891), .B2(new_n702), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n893));
  INV_X1    g468(.A(G106), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n473), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(new_n492), .B2(G130), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n494), .A2(G142), .A3(new_n473), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT113), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n889), .A2(new_n892), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n896), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n891), .A2(new_n639), .A3(new_n702), .ZN(new_n901));
  INV_X1    g476(.A(new_n702), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n888), .B1(new_n902), .B2(new_n890), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n900), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n759), .A2(KEYINPUT112), .A3(new_n760), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n492), .A2(G128), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n908), .A2(new_n511), .A3(new_n828), .A4(new_n830), .ZN(new_n909));
  INV_X1    g484(.A(new_n511), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n831), .B2(new_n833), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(new_n779), .ZN(new_n913));
  OAI221_X1 g488(.A(new_n772), .B1(new_n773), .B2(new_n636), .C1(new_n767), .C2(new_n768), .ZN(new_n914));
  INV_X1    g489(.A(new_n778), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n915), .B2(new_n776), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n909), .A2(new_n911), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n907), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n779), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n761), .B(KEYINPUT112), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n917), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n905), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n887), .B1(new_n924), .B2(KEYINPUT114), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n899), .A2(new_n904), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n906), .B1(new_n920), .B2(new_n922), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n919), .A2(new_n905), .A3(new_n923), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT114), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n925), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n930), .A3(new_n887), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g511(.A1(new_n865), .A2(new_n613), .ZN(new_n937));
  NAND2_X1  g512(.A1(G299), .A2(KEYINPUT115), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT115), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n580), .A2(new_n939), .A3(new_n581), .A4(new_n583), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n622), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(G299), .A2(new_n612), .A3(KEYINPUT115), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n941), .A2(KEYINPUT41), .A3(new_n942), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT41), .B1(new_n941), .B2(new_n942), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n880), .B(new_n625), .ZN(new_n948));
  MUX2_X1   g523(.A(new_n943), .B(new_n947), .S(new_n948), .Z(new_n949));
  XNOR2_X1  g524(.A(G303), .B(G288), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(G305), .ZN(new_n951));
  XNOR2_X1  g526(.A(G290), .B(KEYINPUT116), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT117), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(new_n955), .A3(KEYINPUT42), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n949), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n937), .B1(new_n961), .B2(new_n613), .ZN(G295));
  OAI21_X1  g537(.A(new_n937), .B1(new_n961), .B2(new_n613), .ZN(G331));
  XNOR2_X1  g538(.A(G286), .B(G301), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n880), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n876), .A2(new_n877), .A3(new_n879), .A4(new_n964), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n966), .A2(new_n943), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n946), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n954), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G37), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n878), .B1(new_n571), .B2(new_n865), .ZN(new_n972));
  AOI211_X1 g547(.A(KEYINPUT111), .B(new_n864), .C1(new_n568), .C2(new_n570), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n964), .B1(new_n974), .B2(new_n877), .ZN(new_n975));
  INV_X1    g550(.A(new_n967), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n947), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n966), .A2(new_n943), .A3(new_n967), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n953), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n970), .A2(new_n971), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT118), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n970), .A2(new_n979), .A3(new_n983), .A4(new_n971), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n970), .A2(new_n979), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(KEYINPUT118), .A3(new_n983), .A4(new_n971), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n981), .A2(KEYINPUT44), .A3(new_n984), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(G397));
  INV_X1    g566(.A(G1996), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n916), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n834), .B(G2067), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n779), .A2(G1996), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n703), .A2(new_n708), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n707), .B1(new_n891), .B2(new_n702), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(G1986), .B2(G290), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(G1986), .B2(G290), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n511), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n474), .A2(new_n482), .A3(G40), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n513), .A2(new_n1003), .A3(new_n514), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1007), .B1(new_n1010), .B2(new_n1005), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n511), .A2(new_n1003), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT56), .B(G2072), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1007), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1016), .B(new_n1017), .C1(new_n1010), .C2(KEYINPUT50), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n849), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n1021));
  XNOR2_X1  g596(.A(G299), .B(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1010), .A2(KEYINPUT50), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1007), .B1(new_n1012), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1348), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1016), .A2(new_n1012), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G2067), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1024), .B1(new_n1031), .B2(new_n612), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1015), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT121), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT121), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1019), .A2(new_n1015), .A3(new_n1022), .A4(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT60), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1040), .B2(new_n622), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n1038), .A3(new_n622), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(KEYINPUT60), .A3(new_n1031), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1031), .A2(KEYINPUT60), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1043), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(new_n1041), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1034), .A2(new_n1024), .A3(new_n1036), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT61), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1011), .A2(new_n992), .A3(new_n1013), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT58), .B(G1341), .Z(new_n1053));
  NAND2_X1  g628(.A1(new_n1029), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(KEYINPUT122), .A3(new_n571), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT59), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1055), .A2(KEYINPUT122), .A3(new_n1058), .A4(new_n571), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1024), .A2(KEYINPUT61), .A3(new_n1033), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1051), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1037), .B1(new_n1048), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT125), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1007), .B1(new_n1005), .B2(new_n1004), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n1003), .A4(new_n514), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n813), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1067), .A2(KEYINPUT124), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(KEYINPUT124), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(KEYINPUT53), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1011), .A2(new_n813), .A3(new_n1013), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1073));
  INV_X1    g648(.A(G1961), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1071), .A2(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g651(.A(G301), .B(KEYINPUT54), .Z(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1066), .A2(new_n1006), .A3(new_n1016), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n743), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1025), .A2(new_n1027), .A3(new_n789), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(G168), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1079), .B1(new_n1083), .B2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(G168), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1086));
  OAI211_X1 g661(.A(G8), .B(new_n1083), .C1(new_n1086), .C2(new_n1079), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1076), .A2(new_n1078), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1976), .ZN(new_n1090));
  OAI221_X1 g665(.A(G8), .B1(new_n1090), .B2(G288), .C1(new_n1007), .C2(new_n1004), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n1092));
  INV_X1    g667(.A(G288), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(G1976), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1091), .A2(KEYINPUT52), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1029), .A2(G8), .ZN(new_n1097));
  INV_X1    g672(.A(G1981), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n590), .B2(new_n594), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT120), .B1(G305), .B2(G1981), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n1099), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1097), .B1(new_n1103), .B2(KEYINPUT49), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT49), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1105), .B(new_n1101), .C1(new_n1102), .C2(new_n1099), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1095), .B(new_n1096), .C1(new_n1104), .C2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1971), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1018), .A2(G2090), .ZN(new_n1109));
  OAI21_X1  g684(.A(G8), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AND2_X1   g685(.A1(G303), .A2(G8), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(KEYINPUT119), .A2(KEYINPUT55), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1116), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1073), .A2(G2090), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1118), .B(G8), .C1(new_n1108), .C2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1065), .A2(KEYINPUT53), .A3(new_n813), .A4(new_n1013), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1075), .A2(new_n1077), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1107), .A2(new_n1117), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1064), .B1(new_n1089), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1096), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1095), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1117), .A3(new_n1120), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1128), .A2(new_n1088), .A3(KEYINPUT125), .A4(new_n1122), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1063), .A2(new_n1124), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1087), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n1084), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1085), .A2(new_n1087), .A3(KEYINPUT62), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1127), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(G171), .A3(new_n1076), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1120), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1107), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1139), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n712), .A2(new_n1098), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1097), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1083), .A2(G8), .A3(G168), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1127), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(G8), .B1(new_n1119), .B2(new_n1108), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1143), .B1(new_n1146), .B2(new_n1116), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1144), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1107), .A2(new_n1147), .A3(new_n1120), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1142), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1136), .A2(new_n1138), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1009), .B1(new_n1130), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n994), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1008), .B1(new_n1153), .B2(new_n779), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1008), .A2(new_n992), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT46), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT47), .ZN(new_n1158));
  INV_X1    g733(.A(G2067), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n834), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n996), .B2(new_n998), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n1008), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT126), .Z(new_n1163));
  NAND2_X1  g738(.A1(new_n1000), .A2(new_n1008), .ZN(new_n1164));
  NOR4_X1   g739(.A1(new_n1006), .A2(new_n1007), .A3(G290), .A4(G1986), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT48), .Z(new_n1166));
  AOI21_X1  g741(.A(new_n1163), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1152), .A2(new_n1158), .A3(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g743(.A(G227), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n658), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1171), .B1(new_n933), .B2(new_n934), .ZN(new_n1172));
  NOR2_X1   g746(.A1(G229), .A2(new_n460), .ZN(new_n1173));
  AND4_X1   g747(.A1(new_n988), .A2(new_n985), .A3(new_n1172), .A4(new_n1173), .ZN(G308));
  NAND4_X1  g748(.A1(new_n985), .A2(new_n1172), .A3(new_n988), .A4(new_n1173), .ZN(G225));
endmodule


