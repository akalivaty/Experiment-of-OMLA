

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748;

  INV_X1 U371 ( .A(n376), .ZN(n350) );
  INV_X1 U372 ( .A(n570), .ZN(n353) );
  INV_X1 U373 ( .A(n385), .ZN(n352) );
  XNOR2_X1 U374 ( .A(n652), .B(KEYINPUT6), .ZN(n592) );
  BUF_X1 U375 ( .A(n538), .Z(n652) );
  XNOR2_X1 U376 ( .A(n486), .B(n485), .ZN(n527) );
  OR2_X1 U377 ( .A1(n711), .A2(G902), .ZN(n486) );
  INV_X1 U378 ( .A(KEYINPUT64), .ZN(n398) );
  XNOR2_X2 U379 ( .A(n462), .B(G134), .ZN(n443) );
  INV_X1 U380 ( .A(n347), .ZN(n567) );
  NAND2_X1 U381 ( .A1(n557), .A2(n348), .ZN(n347) );
  NOR2_X1 U382 ( .A1(n349), .A2(n558), .ZN(n348) );
  INV_X1 U383 ( .A(n556), .ZN(n349) );
  NAND2_X1 U384 ( .A1(n351), .A2(n350), .ZN(n375) );
  NAND2_X1 U385 ( .A1(n353), .A2(n352), .ZN(n351) );
  NOR2_X1 U386 ( .A1(n526), .A2(n667), .ZN(n490) );
  BUF_X1 U387 ( .A(n607), .Z(n723) );
  XNOR2_X2 U388 ( .A(n528), .B(KEYINPUT93), .ZN(n562) );
  XNOR2_X2 U389 ( .A(n737), .B(n459), .ZN(n483) );
  NAND2_X1 U390 ( .A1(n655), .A2(n541), .ZN(n528) );
  NOR2_X2 U391 ( .A1(n372), .A2(n371), .ZN(n605) );
  NAND2_X1 U392 ( .A1(n374), .A2(n373), .ZN(n372) );
  AND2_X1 U393 ( .A1(n375), .A2(n578), .ZN(n374) );
  OR2_X1 U394 ( .A1(n385), .A2(KEYINPUT48), .ZN(n354) );
  NOR2_X1 U395 ( .A1(n550), .A2(n549), .ZN(n632) );
  NOR2_X1 U396 ( .A1(n572), .A2(n575), .ZN(n477) );
  NOR2_X1 U397 ( .A1(n648), .A2(n501), .ZN(n502) );
  XNOR2_X1 U398 ( .A(n490), .B(n489), .ZN(n548) );
  XNOR2_X1 U399 ( .A(n440), .B(n439), .ZN(n511) );
  NOR2_X2 U400 ( .A1(n506), .A2(n503), .ZN(n504) );
  XNOR2_X1 U401 ( .A(n369), .B(n368), .ZN(n520) );
  OR2_X2 U402 ( .A1(n610), .A2(G902), .ZN(n451) );
  XNOR2_X2 U403 ( .A(n443), .B(n442), .ZN(n737) );
  XNOR2_X1 U404 ( .A(n547), .B(n546), .ZN(n378) );
  XNOR2_X1 U405 ( .A(KEYINPUT46), .B(KEYINPUT65), .ZN(n546) );
  XNOR2_X1 U406 ( .A(KEYINPUT3), .B(G119), .ZN(n444) );
  AND2_X1 U407 ( .A1(n380), .A2(n379), .ZN(n560) );
  INV_X1 U408 ( .A(n524), .ZN(n379) );
  XNOR2_X1 U409 ( .A(n381), .B(n523), .ZN(n380) );
  AND2_X1 U410 ( .A1(n511), .A2(n647), .ZN(n655) );
  BUF_X1 U411 ( .A(n527), .Z(n541) );
  NAND2_X1 U412 ( .A1(n548), .A2(n494), .ZN(n496) );
  XNOR2_X1 U413 ( .A(n536), .B(n535), .ZN(n692) );
  NAND2_X1 U414 ( .A1(n507), .A2(n501), .ZN(n594) );
  BUF_X1 U415 ( .A(n454), .Z(n740) );
  XNOR2_X1 U416 ( .A(n400), .B(n399), .ZN(n426) );
  XNOR2_X1 U417 ( .A(G131), .B(G143), .ZN(n387) );
  NOR2_X1 U418 ( .A1(n378), .A2(n376), .ZN(n371) );
  XNOR2_X1 U419 ( .A(n527), .B(KEYINPUT1), .ZN(n512) );
  AND2_X1 U420 ( .A1(n592), .A2(n367), .ZN(n366) );
  NAND2_X1 U421 ( .A1(n361), .A2(n360), .ZN(n363) );
  NAND2_X1 U422 ( .A1(n365), .A2(n364), .ZN(n361) );
  OR2_X1 U423 ( .A1(n592), .A2(n367), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n483), .B(n450), .ZN(n610) );
  NOR2_X1 U425 ( .A1(n529), .A2(n586), .ZN(n530) );
  NAND2_X1 U426 ( .A1(n363), .A2(n359), .ZN(n369) );
  NOR2_X1 U427 ( .A1(n366), .A2(n587), .ZN(n359) );
  INV_X1 U428 ( .A(KEYINPUT34), .ZN(n368) );
  BUF_X1 U429 ( .A(n526), .Z(n575) );
  INV_X1 U430 ( .A(KEYINPUT19), .ZN(n489) );
  XNOR2_X1 U431 ( .A(n483), .B(n482), .ZN(n711) );
  XNOR2_X1 U432 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n544) );
  INV_X1 U433 ( .A(KEYINPUT100), .ZN(n508) );
  OR2_X1 U434 ( .A1(n594), .A2(n593), .ZN(n623) );
  INV_X1 U435 ( .A(n667), .ZN(n382) );
  XNOR2_X1 U436 ( .A(KEYINPUT83), .B(KEYINPUT45), .ZN(n355) );
  INV_X1 U437 ( .A(KEYINPUT48), .ZN(n376) );
  NOR2_X1 U438 ( .A1(n511), .A2(n592), .ZN(n452) );
  NOR2_X2 U439 ( .A1(n596), .A2(n607), .ZN(n597) );
  XNOR2_X2 U440 ( .A(n496), .B(n495), .ZN(n516) );
  XNOR2_X2 U441 ( .A(n356), .B(n355), .ZN(n607) );
  NAND2_X1 U442 ( .A1(n357), .A2(n384), .ZN(n356) );
  XNOR2_X1 U443 ( .A(n358), .B(KEYINPUT44), .ZN(n357) );
  NOR2_X2 U444 ( .A1(n582), .A2(n581), .ZN(n358) );
  NAND2_X1 U445 ( .A1(n514), .A2(n515), .ZN(n360) );
  NAND2_X1 U446 ( .A1(n363), .A2(n362), .ZN(n665) );
  INV_X1 U447 ( .A(n366), .ZN(n362) );
  INV_X1 U448 ( .A(n514), .ZN(n365) );
  INV_X1 U449 ( .A(n515), .ZN(n367) );
  NAND2_X1 U450 ( .A1(n370), .A2(n378), .ZN(n373) );
  NOR2_X1 U451 ( .A1(n570), .A2(n354), .ZN(n370) );
  INV_X1 U452 ( .A(n538), .ZN(n589) );
  NAND2_X1 U453 ( .A1(n538), .A2(n382), .ZN(n381) );
  INV_X1 U454 ( .A(n506), .ZN(n507) );
  BUF_X1 U455 ( .A(n708), .Z(n718) );
  BUF_X1 U456 ( .A(n582), .Z(n522) );
  XOR2_X1 U457 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n383) );
  AND2_X1 U458 ( .A1(n595), .A2(n623), .ZN(n384) );
  AND2_X1 U459 ( .A1(n569), .A2(KEYINPUT47), .ZN(n385) );
  INV_X1 U460 ( .A(KEYINPUT101), .ZN(n513) );
  INV_X1 U461 ( .A(KEYINPUT30), .ZN(n523) );
  BUF_X1 U462 ( .A(n605), .Z(n738) );
  XNOR2_X1 U463 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U464 ( .A(n434), .B(n433), .ZN(n720) );
  OR2_X1 U465 ( .A1(n740), .A2(G952), .ZN(n699) );
  XNOR2_X1 U466 ( .A(n594), .B(n508), .ZN(n510) );
  XNOR2_X1 U467 ( .A(n545), .B(n544), .ZN(n747) );
  XNOR2_X1 U468 ( .A(KEYINPUT13), .B(G475), .ZN(n397) );
  XNOR2_X1 U469 ( .A(G125), .B(KEYINPUT10), .ZN(n386) );
  XNOR2_X1 U470 ( .A(n386), .B(G140), .ZN(n736) );
  XNOR2_X1 U471 ( .A(G146), .B(n736), .ZN(n432) );
  INV_X1 U472 ( .A(n432), .ZN(n390) );
  NOR2_X1 U473 ( .A1(G953), .A2(G237), .ZN(n446) );
  NAND2_X1 U474 ( .A1(G214), .A2(n446), .ZN(n388) );
  XNOR2_X1 U475 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U476 ( .A(n390), .B(n389), .ZN(n395) );
  XOR2_X1 U477 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n392) );
  XNOR2_X1 U478 ( .A(G113), .B(KEYINPUT12), .ZN(n391) );
  XNOR2_X1 U479 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U480 ( .A(G122), .B(G104), .ZN(n470) );
  XOR2_X1 U481 ( .A(n393), .B(n470), .Z(n394) );
  XNOR2_X1 U482 ( .A(n395), .B(n394), .ZN(n616) );
  NOR2_X1 U483 ( .A1(G902), .A2(n616), .ZN(n396) );
  XNOR2_X1 U484 ( .A(n397), .B(n396), .ZN(n517) );
  INV_X1 U485 ( .A(n517), .ZN(n551) );
  XOR2_X1 U486 ( .A(KEYINPUT97), .B(KEYINPUT7), .Z(n402) );
  XNOR2_X2 U487 ( .A(n398), .B(G953), .ZN(n454) );
  NAND2_X1 U488 ( .A1(n454), .A2(G234), .ZN(n400) );
  XOR2_X1 U489 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n399) );
  NAND2_X1 U490 ( .A1(G217), .A2(n426), .ZN(n401) );
  XNOR2_X1 U491 ( .A(n402), .B(n401), .ZN(n409) );
  XNOR2_X2 U492 ( .A(G143), .B(KEYINPUT78), .ZN(n404) );
  INV_X1 U493 ( .A(G128), .ZN(n403) );
  XNOR2_X2 U494 ( .A(n404), .B(n403), .ZN(n462) );
  XOR2_X1 U495 ( .A(KEYINPUT9), .B(G107), .Z(n406) );
  XNOR2_X1 U496 ( .A(G116), .B(G122), .ZN(n405) );
  XNOR2_X1 U497 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U498 ( .A(n443), .B(n407), .ZN(n408) );
  XNOR2_X1 U499 ( .A(n409), .B(n408), .ZN(n715) );
  NOR2_X1 U500 ( .A1(G902), .A2(n715), .ZN(n410) );
  XOR2_X1 U501 ( .A(G478), .B(n410), .Z(n552) );
  OR2_X1 U502 ( .A1(n551), .A2(n552), .ZN(n638) );
  XNOR2_X1 U503 ( .A(G902), .B(KEYINPUT15), .ZN(n598) );
  NAND2_X1 U504 ( .A1(n598), .A2(G234), .ZN(n411) );
  XNOR2_X1 U505 ( .A(n411), .B(KEYINPUT20), .ZN(n435) );
  AND2_X1 U506 ( .A1(n435), .A2(G221), .ZN(n412) );
  XNOR2_X1 U507 ( .A(n412), .B(KEYINPUT21), .ZN(n647) );
  INV_X1 U508 ( .A(n647), .ZN(n419) );
  NAND2_X1 U509 ( .A1(G234), .A2(G237), .ZN(n413) );
  XNOR2_X1 U510 ( .A(n413), .B(KEYINPUT14), .ZN(n414) );
  XNOR2_X1 U511 ( .A(KEYINPUT72), .B(n414), .ZN(n415) );
  NAND2_X1 U512 ( .A1(G952), .A2(n415), .ZN(n683) );
  NOR2_X1 U513 ( .A1(n683), .A2(G953), .ZN(n493) );
  NAND2_X1 U514 ( .A1(G902), .A2(n415), .ZN(n491) );
  NOR2_X1 U515 ( .A1(n740), .A2(n491), .ZN(n416) );
  XNOR2_X1 U516 ( .A(n416), .B(KEYINPUT103), .ZN(n417) );
  NOR2_X1 U517 ( .A1(G900), .A2(n417), .ZN(n418) );
  NOR2_X1 U518 ( .A1(n493), .A2(n418), .ZN(n524) );
  NOR2_X1 U519 ( .A1(n419), .A2(n524), .ZN(n537) );
  INV_X1 U520 ( .A(G902), .ZN(n421) );
  INV_X1 U521 ( .A(G237), .ZN(n420) );
  NAND2_X1 U522 ( .A1(n421), .A2(n420), .ZN(n474) );
  NAND2_X1 U523 ( .A1(n474), .A2(G214), .ZN(n422) );
  XNOR2_X1 U524 ( .A(n422), .B(KEYINPUT89), .ZN(n667) );
  NAND2_X1 U525 ( .A1(n537), .A2(n382), .ZN(n423) );
  NOR2_X1 U526 ( .A1(n638), .A2(n423), .ZN(n453) );
  XNOR2_X1 U527 ( .A(G119), .B(G128), .ZN(n424) );
  XNOR2_X1 U528 ( .A(n383), .B(n424), .ZN(n425) );
  XOR2_X1 U529 ( .A(G137), .B(n425), .Z(n428) );
  NAND2_X1 U530 ( .A1(n426), .A2(G221), .ZN(n427) );
  XNOR2_X1 U531 ( .A(n428), .B(n427), .ZN(n434) );
  XOR2_X1 U532 ( .A(KEYINPUT90), .B(KEYINPUT74), .Z(n430) );
  XNOR2_X1 U533 ( .A(G110), .B(KEYINPUT91), .ZN(n429) );
  XNOR2_X1 U534 ( .A(n430), .B(n429), .ZN(n431) );
  NOR2_X1 U535 ( .A1(n720), .A2(G902), .ZN(n440) );
  XOR2_X1 U536 ( .A(KEYINPUT92), .B(KEYINPUT73), .Z(n437) );
  NAND2_X1 U537 ( .A1(n435), .A2(G217), .ZN(n436) );
  XNOR2_X1 U538 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U539 ( .A(n438), .B(KEYINPUT25), .ZN(n439) );
  XNOR2_X1 U540 ( .A(KEYINPUT4), .B(G146), .ZN(n458) );
  XNOR2_X1 U541 ( .A(G137), .B(G131), .ZN(n441) );
  XNOR2_X1 U542 ( .A(n458), .B(n441), .ZN(n442) );
  XNOR2_X1 U543 ( .A(KEYINPUT68), .B(G101), .ZN(n459) );
  XNOR2_X1 U544 ( .A(G116), .B(G113), .ZN(n445) );
  XNOR2_X1 U545 ( .A(n445), .B(n444), .ZN(n469) );
  NAND2_X1 U546 ( .A1(n446), .A2(G210), .ZN(n448) );
  INV_X1 U547 ( .A(KEYINPUT5), .ZN(n447) );
  XNOR2_X1 U548 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U549 ( .A(n469), .B(n449), .ZN(n450) );
  XNOR2_X2 U550 ( .A(n451), .B(G472), .ZN(n538) );
  NAND2_X1 U551 ( .A1(n453), .A2(n452), .ZN(n572) );
  NAND2_X1 U552 ( .A1(n454), .A2(G224), .ZN(n457) );
  XNOR2_X2 U553 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n455) );
  XNOR2_X1 U554 ( .A(n455), .B(KEYINPUT88), .ZN(n456) );
  XNOR2_X1 U555 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U556 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U557 ( .A(n461), .B(n460), .ZN(n468) );
  INV_X1 U558 ( .A(n462), .ZN(n466) );
  XNOR2_X1 U559 ( .A(G125), .B(KEYINPUT17), .ZN(n464) );
  XNOR2_X1 U560 ( .A(KEYINPUT18), .B(KEYINPUT87), .ZN(n463) );
  XNOR2_X1 U561 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U562 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U563 ( .A(n468), .B(n467), .ZN(n473) );
  XNOR2_X1 U564 ( .A(G110), .B(G107), .ZN(n479) );
  XNOR2_X1 U565 ( .A(n469), .B(n479), .ZN(n472) );
  XNOR2_X1 U566 ( .A(n470), .B(KEYINPUT16), .ZN(n471) );
  XNOR2_X1 U567 ( .A(n472), .B(n471), .ZN(n730) );
  XNOR2_X1 U568 ( .A(n473), .B(n730), .ZN(n700) );
  INV_X1 U569 ( .A(n598), .ZN(n600) );
  OR2_X2 U570 ( .A1(n700), .A2(n600), .ZN(n476) );
  NAND2_X1 U571 ( .A1(n474), .A2(G210), .ZN(n475) );
  XNOR2_X2 U572 ( .A(n476), .B(n475), .ZN(n526) );
  XNOR2_X1 U573 ( .A(n477), .B(KEYINPUT36), .ZN(n487) );
  XNOR2_X1 U574 ( .A(G104), .B(G140), .ZN(n478) );
  XNOR2_X1 U575 ( .A(n479), .B(n478), .ZN(n481) );
  NAND2_X1 U576 ( .A1(n740), .A2(G227), .ZN(n480) );
  XNOR2_X1 U577 ( .A(n481), .B(n480), .ZN(n482) );
  INV_X1 U578 ( .A(KEYINPUT71), .ZN(n484) );
  XNOR2_X1 U579 ( .A(n484), .B(G469), .ZN(n485) );
  BUF_X2 U580 ( .A(n512), .Z(n654) );
  NAND2_X1 U581 ( .A1(n487), .A2(n654), .ZN(n557) );
  XOR2_X1 U582 ( .A(G125), .B(KEYINPUT37), .Z(n488) );
  XNOR2_X1 U583 ( .A(n557), .B(n488), .ZN(G27) );
  INV_X1 U584 ( .A(G898), .ZN(n726) );
  NAND2_X1 U585 ( .A1(G953), .A2(n726), .ZN(n731) );
  NOR2_X1 U586 ( .A1(n491), .A2(n731), .ZN(n492) );
  OR2_X1 U587 ( .A1(n493), .A2(n492), .ZN(n494) );
  INV_X1 U588 ( .A(KEYINPUT0), .ZN(n495) );
  NOR2_X1 U589 ( .A1(n552), .A2(n517), .ZN(n497) );
  XNOR2_X1 U590 ( .A(n497), .B(KEYINPUT98), .ZN(n669) );
  AND2_X1 U591 ( .A1(n669), .A2(n647), .ZN(n498) );
  NAND2_X1 U592 ( .A1(n516), .A2(n498), .ZN(n500) );
  XNOR2_X1 U593 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n499) );
  XNOR2_X1 U594 ( .A(n500), .B(n499), .ZN(n506) );
  XOR2_X1 U595 ( .A(KEYINPUT99), .B(n511), .Z(n648) );
  INV_X1 U596 ( .A(n654), .ZN(n501) );
  NAND2_X1 U597 ( .A1(n502), .A2(n592), .ZN(n503) );
  XOR2_X1 U598 ( .A(KEYINPUT32), .B(n504), .Z(n579) );
  XNOR2_X1 U599 ( .A(G119), .B(KEYINPUT126), .ZN(n505) );
  XNOR2_X1 U600 ( .A(n579), .B(n505), .ZN(G21) );
  NOR2_X1 U601 ( .A1(n511), .A2(n652), .ZN(n509) );
  NAND2_X1 U602 ( .A1(n510), .A2(n509), .ZN(n580) );
  XNOR2_X1 U603 ( .A(n580), .B(G110), .ZN(G12) );
  NAND2_X1 U604 ( .A1(n655), .A2(n512), .ZN(n583) );
  XNOR2_X1 U605 ( .A(n583), .B(n513), .ZN(n514) );
  XNOR2_X1 U606 ( .A(KEYINPUT86), .B(KEYINPUT33), .ZN(n515) );
  INV_X1 U607 ( .A(n516), .ZN(n587) );
  NAND2_X1 U608 ( .A1(n517), .A2(n552), .ZN(n518) );
  XOR2_X1 U609 ( .A(n518), .B(KEYINPUT102), .Z(n565) );
  XOR2_X1 U610 ( .A(KEYINPUT77), .B(n565), .Z(n519) );
  NAND2_X1 U611 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U612 ( .A(n521), .B(KEYINPUT35), .ZN(n582) );
  XOR2_X1 U613 ( .A(n522), .B(G122), .Z(G24) );
  INV_X1 U614 ( .A(KEYINPUT38), .ZN(n525) );
  XNOR2_X1 U615 ( .A(n526), .B(n525), .ZN(n533) );
  INV_X1 U616 ( .A(n533), .ZN(n666) );
  NAND2_X1 U617 ( .A1(n560), .A2(n666), .ZN(n529) );
  INV_X1 U618 ( .A(n562), .ZN(n586) );
  XNOR2_X1 U619 ( .A(n530), .B(KEYINPUT39), .ZN(n571) );
  NOR2_X1 U620 ( .A1(n571), .A2(n638), .ZN(n532) );
  XNOR2_X1 U621 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n531) );
  XNOR2_X1 U622 ( .A(n532), .B(n531), .ZN(n748) );
  NOR2_X1 U623 ( .A1(n533), .A2(n667), .ZN(n534) );
  XNOR2_X1 U624 ( .A(n534), .B(KEYINPUT106), .ZN(n673) );
  NAND2_X1 U625 ( .A1(n673), .A2(n669), .ZN(n536) );
  XOR2_X1 U626 ( .A(KEYINPUT41), .B(KEYINPUT107), .Z(n535) );
  NAND2_X1 U627 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U628 ( .A1(n511), .A2(n539), .ZN(n540) );
  XNOR2_X1 U629 ( .A(KEYINPUT28), .B(n540), .ZN(n542) );
  NAND2_X1 U630 ( .A1(n542), .A2(n541), .ZN(n550) );
  INV_X1 U631 ( .A(n550), .ZN(n543) );
  NAND2_X1 U632 ( .A1(n692), .A2(n543), .ZN(n545) );
  NAND2_X1 U633 ( .A1(n748), .A2(n747), .ZN(n547) );
  INV_X1 U634 ( .A(n548), .ZN(n549) );
  XNOR2_X1 U635 ( .A(KEYINPUT69), .B(KEYINPUT47), .ZN(n553) );
  NAND2_X1 U636 ( .A1(n552), .A2(n551), .ZN(n642) );
  NAND2_X1 U637 ( .A1(n638), .A2(n642), .ZN(n672) );
  NAND2_X1 U638 ( .A1(n553), .A2(n672), .ZN(n554) );
  NAND2_X1 U639 ( .A1(n554), .A2(KEYINPUT80), .ZN(n555) );
  NAND2_X1 U640 ( .A1(n632), .A2(n555), .ZN(n556) );
  NOR2_X1 U641 ( .A1(KEYINPUT80), .A2(KEYINPUT47), .ZN(n558) );
  INV_X1 U642 ( .A(n560), .ZN(n561) );
  NOR2_X1 U643 ( .A1(n561), .A2(n575), .ZN(n563) );
  NAND2_X1 U644 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U645 ( .A(KEYINPUT104), .B(n564), .Z(n566) );
  NAND2_X1 U646 ( .A1(n566), .A2(n565), .ZN(n635) );
  NAND2_X1 U647 ( .A1(n567), .A2(n635), .ZN(n570) );
  INV_X1 U648 ( .A(n632), .ZN(n636) );
  NAND2_X1 U649 ( .A1(n636), .A2(KEYINPUT80), .ZN(n568) );
  NAND2_X1 U650 ( .A1(n568), .A2(n672), .ZN(n569) );
  OR2_X1 U651 ( .A1(n642), .A2(n571), .ZN(n646) );
  INV_X1 U652 ( .A(n646), .ZN(n577) );
  NOR2_X1 U653 ( .A1(n572), .A2(n654), .ZN(n574) );
  INV_X1 U654 ( .A(KEYINPUT43), .ZN(n573) );
  XNOR2_X1 U655 ( .A(n574), .B(n573), .ZN(n576) );
  AND2_X1 U656 ( .A1(n576), .A2(n575), .ZN(n622) );
  NOR2_X1 U657 ( .A1(n577), .A2(n622), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n605), .A2(KEYINPUT82), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U660 ( .A1(n583), .A2(n589), .ZN(n584) );
  XNOR2_X1 U661 ( .A(n584), .B(KEYINPUT95), .ZN(n660) );
  NOR2_X1 U662 ( .A1(n660), .A2(n587), .ZN(n585) );
  XNOR2_X1 U663 ( .A(n585), .B(KEYINPUT31), .ZN(n641) );
  NOR2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U665 ( .A(KEYINPUT94), .B(n588), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n625) );
  NAND2_X1 U667 ( .A1(n641), .A2(n625), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n591), .A2(n672), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n648), .A2(n592), .ZN(n593) );
  NOR2_X1 U670 ( .A1(n597), .A2(KEYINPUT2), .ZN(n599) );
  NOR2_X2 U671 ( .A1(n599), .A2(n598), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n600), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n607), .A2(n601), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n602), .A2(KEYINPUT82), .ZN(n603) );
  NOR2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n605), .A2(KEYINPUT2), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT84), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n608), .A2(n723), .ZN(n690) );
  NOR2_X2 U679 ( .A1(n609), .A2(n690), .ZN(n708) );
  NAND2_X1 U680 ( .A1(n708), .A2(G472), .ZN(n612) );
  XOR2_X1 U681 ( .A(KEYINPUT62), .B(n610), .Z(n611) );
  XNOR2_X1 U682 ( .A(n612), .B(n611), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n613), .A2(n699), .ZN(n615) );
  XOR2_X1 U684 ( .A(KEYINPUT109), .B(KEYINPUT63), .Z(n614) );
  XNOR2_X1 U685 ( .A(n615), .B(n614), .ZN(G57) );
  NAND2_X1 U686 ( .A1(n708), .A2(G475), .ZN(n618) );
  XNOR2_X1 U687 ( .A(n616), .B(KEYINPUT59), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(n619) );
  NAND2_X1 U689 ( .A1(n619), .A2(n699), .ZN(n621) );
  XNOR2_X1 U690 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(G60) );
  XOR2_X1 U692 ( .A(G140), .B(n622), .Z(G42) );
  XNOR2_X1 U693 ( .A(G101), .B(n623), .ZN(G3) );
  NOR2_X1 U694 ( .A1(n638), .A2(n625), .ZN(n624) );
  XOR2_X1 U695 ( .A(G104), .B(n624), .Z(G6) );
  NOR2_X1 U696 ( .A1(n642), .A2(n625), .ZN(n630) );
  XOR2_X1 U697 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n627) );
  XNOR2_X1 U698 ( .A(G107), .B(KEYINPUT26), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U700 ( .A(KEYINPUT110), .B(n628), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(n629), .ZN(G9) );
  XOR2_X1 U702 ( .A(G128), .B(KEYINPUT29), .Z(n634) );
  INV_X1 U703 ( .A(n642), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n634), .B(n633), .ZN(G30) );
  XNOR2_X1 U706 ( .A(G143), .B(n635), .ZN(G45) );
  NOR2_X1 U707 ( .A1(n636), .A2(n638), .ZN(n637) );
  XOR2_X1 U708 ( .A(G146), .B(n637), .Z(G48) );
  NOR2_X1 U709 ( .A1(n638), .A2(n641), .ZN(n639) );
  XOR2_X1 U710 ( .A(KEYINPUT112), .B(n639), .Z(n640) );
  XNOR2_X1 U711 ( .A(G113), .B(n640), .ZN(G15) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n644) );
  XNOR2_X1 U713 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U715 ( .A(G116), .B(n645), .ZN(G18) );
  XNOR2_X1 U716 ( .A(G134), .B(n646), .ZN(G36) );
  XNOR2_X1 U717 ( .A(KEYINPUT121), .B(KEYINPUT52), .ZN(n681) );
  NOR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U719 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT116), .ZN(n659) );
  XOR2_X1 U723 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n657) );
  NOR2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U725 ( .A(n657), .B(n656), .Z(n658) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n661) );
  NAND2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n663) );
  XOR2_X1 U728 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n662) );
  XNOR2_X1 U729 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n664), .A2(n692), .ZN(n679) );
  INV_X1 U731 ( .A(n665), .ZN(n677) );
  NAND2_X1 U732 ( .A1(n533), .A2(n667), .ZN(n668) );
  XOR2_X1 U733 ( .A(KEYINPUT119), .B(n668), .Z(n670) );
  NAND2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U735 ( .A(n671), .B(KEYINPUT120), .ZN(n675) );
  NAND2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U739 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U742 ( .A1(G953), .A2(n684), .ZN(n697) );
  XOR2_X1 U743 ( .A(KEYINPUT2), .B(KEYINPUT79), .Z(n686) );
  NOR2_X1 U744 ( .A1(n738), .A2(n686), .ZN(n685) );
  XNOR2_X1 U745 ( .A(n685), .B(KEYINPUT81), .ZN(n689) );
  INV_X1 U746 ( .A(n686), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n723), .A2(n687), .ZN(n688) );
  NAND2_X1 U748 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n695) );
  INV_X1 U750 ( .A(n692), .ZN(n693) );
  NOR2_X1 U751 ( .A1(n693), .A2(n665), .ZN(n694) );
  NOR2_X1 U752 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U754 ( .A(KEYINPUT53), .B(n698), .Z(G75) );
  INV_X1 U755 ( .A(n699), .ZN(n722) );
  NAND2_X1 U756 ( .A1(n708), .A2(G210), .ZN(n705) );
  BUF_X1 U757 ( .A(n700), .Z(n703) );
  XOR2_X1 U758 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n701) );
  XOR2_X1 U759 ( .A(n701), .B(KEYINPUT85), .Z(n702) );
  XNOR2_X1 U760 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U761 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X2 U762 ( .A1(n722), .A2(n706), .ZN(n707) );
  XNOR2_X1 U763 ( .A(KEYINPUT56), .B(n707), .ZN(G51) );
  NAND2_X1 U764 ( .A1(n718), .A2(G469), .ZN(n713) );
  XOR2_X1 U765 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n709) );
  XNOR2_X1 U766 ( .A(n709), .B(KEYINPUT122), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U768 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U769 ( .A1(n722), .A2(n714), .ZN(G54) );
  NAND2_X1 U770 ( .A1(n718), .A2(G478), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U772 ( .A1(n722), .A2(n717), .ZN(G63) );
  NAND2_X1 U773 ( .A1(n718), .A2(G217), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U775 ( .A1(n722), .A2(n721), .ZN(G66) );
  NOR2_X1 U776 ( .A1(n723), .A2(G953), .ZN(n728) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n724) );
  XOR2_X1 U778 ( .A(KEYINPUT61), .B(n724), .Z(n725) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n734) );
  XNOR2_X1 U781 ( .A(G101), .B(KEYINPUT123), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n730), .B(n729), .ZN(n732) );
  NAND2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U785 ( .A(KEYINPUT124), .B(n735), .ZN(G69) );
  XOR2_X1 U786 ( .A(n737), .B(n736), .Z(n741) );
  XNOR2_X1 U787 ( .A(n738), .B(n741), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n740), .A2(n739), .ZN(n745) );
  XOR2_X1 U789 ( .A(G227), .B(n741), .Z(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(G900), .ZN(n743) );
  NAND2_X1 U791 ( .A1(G953), .A2(n743), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U793 ( .A(KEYINPUT125), .B(n746), .Z(G72) );
  XNOR2_X1 U794 ( .A(n747), .B(G137), .ZN(G39) );
  XNOR2_X1 U795 ( .A(n748), .B(G131), .ZN(G33) );
endmodule

