//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n632, new_n635, new_n637, new_n638, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n464), .A2(G2105), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n470), .A2(new_n474), .B1(G101), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(new_n465), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n473), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n480), .B2(new_n481), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n476), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n466), .A2(new_n469), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n473), .C2(G112), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n488), .A2(new_n473), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G124), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n490), .B(new_n491), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  XNOR2_X1  g074(.A(new_n499), .B(KEYINPUT70), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n466), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n473), .A2(G138), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n470), .A2(KEYINPUT71), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(new_n488), .B2(new_n503), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n505), .A2(KEYINPUT4), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n478), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n504), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n502), .B1(new_n508), .B2(new_n513), .ZN(G164));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G62), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(KEYINPUT74), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(KEYINPUT74), .B1(G75), .B2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n515), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n517), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(new_n526), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(new_n520), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT73), .B(G88), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n524), .A2(new_n532), .ZN(G166));
  NAND2_X1  g108(.A1(new_n527), .A2(G51), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT75), .B(G89), .Z(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n536), .A2(new_n540), .ZN(G168));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n518), .B2(new_n519), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT76), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n547));
  AND2_X1   g122(.A1(KEYINPUT5), .A2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(KEYINPUT5), .A2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n547), .B(new_n544), .C1(new_n550), .C2(new_n542), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(G651), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n525), .A2(new_n526), .B1(new_n518), .B2(new_n519), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT77), .B(G90), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n553), .A2(new_n554), .B1(new_n527), .B2(G52), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  NAND2_X1  g132(.A1(new_n527), .A2(G43), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n530), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(new_n515), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n518), .B2(new_n519), .ZN(new_n570));
  AND2_X1   g145(.A1(G78), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n553), .A2(G91), .ZN(new_n573));
  AND2_X1   g148(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n574));
  NOR2_X1   g149(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n527), .B2(G53), .ZN(new_n577));
  INV_X1    g152(.A(new_n526), .ZN(new_n578));
  NOR2_X1   g153(.A1(KEYINPUT6), .A2(G651), .ZN(new_n579));
  OAI211_X1 g154(.A(G53), .B(G543), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n574), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n572), .B(new_n573), .C1(new_n577), .C2(new_n581), .ZN(G299));
  OR2_X1    g157(.A1(new_n536), .A2(new_n540), .ZN(G286));
  INV_X1    g158(.A(G166), .ZN(G303));
  OAI21_X1  g159(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n529), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n553), .A2(G87), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n553), .A2(G86), .B1(new_n527), .B2(G48), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n520), .A2(G61), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n515), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n594), .A2(KEYINPUT79), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(KEYINPUT79), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(G305));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  INV_X1    g173(.A(G72), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n550), .A2(new_n598), .B1(new_n599), .B2(new_n517), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n515), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n601), .B2(new_n600), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n553), .A2(G85), .B1(new_n527), .B2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(KEYINPUT81), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n518), .B2(new_n519), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(KEYINPUT82), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n615), .A2(G79), .A3(G543), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(G651), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n527), .A2(G54), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n618), .A2(KEYINPUT83), .A3(new_n619), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n624));
  INV_X1    g199(.A(G92), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n530), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n553), .A2(KEYINPUT10), .A3(G92), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n622), .A2(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n610), .B1(new_n628), .B2(G868), .ZN(G284));
  OAI21_X1  g204(.A(new_n610), .B1(new_n628), .B2(G868), .ZN(G321));
  NAND2_X1  g205(.A1(G286), .A2(G868), .ZN(new_n631));
  INV_X1    g206(.A(G299), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G868), .ZN(G297));
  OAI21_X1  g208(.A(new_n631), .B1(new_n632), .B2(G868), .ZN(G280));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n628), .B1(new_n635), .B2(G860), .ZN(G148));
  NAND2_X1  g211(.A1(new_n628), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g214(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n640));
  XNOR2_X1  g215(.A(G323), .B(new_n640), .ZN(G282));
  NAND2_X1  g216(.A1(new_n509), .A2(new_n475), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT13), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n489), .A2(G135), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n492), .A2(G123), .ZN(new_n647));
  OAI221_X1 g222(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n473), .C2(G111), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT85), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n645), .A2(new_n651), .ZN(G156));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(KEYINPUT14), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT87), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G1341), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(KEYINPUT87), .ZN(new_n667));
  INV_X1    g242(.A(G1341), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(KEYINPUT87), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(G1348), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n671), .B1(new_n666), .B2(new_n670), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n658), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n674), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n676), .A2(new_n657), .A3(new_n672), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n677), .A3(G14), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT88), .ZN(G401));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(new_n683), .B2(KEYINPUT18), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT89), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT90), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT18), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(KEYINPUT17), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n681), .A2(new_n682), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2096), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n687), .B(new_n692), .ZN(G227));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1956), .B(G2474), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1961), .B(G1966), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n697), .A2(KEYINPUT92), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n703), .B(new_n704), .Z(new_n705));
  NOR3_X1   g280(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT20), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n708), .B1(new_n705), .B2(new_n707), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n694), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(new_n694), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n713), .A2(new_n714), .A3(new_n709), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n712), .A2(new_n715), .A3(new_n717), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(G229));
  NAND2_X1  g297(.A1(G166), .A2(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G16), .B2(G22), .ZN(new_n724));
  INV_X1    g299(.A(G1971), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n727), .A2(G6), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G305), .B2(G16), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT32), .B(G1981), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n724), .A2(new_n725), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n726), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n727), .A2(G23), .ZN(new_n734));
  INV_X1    g309(.A(G288), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n727), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT33), .B(G1976), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n730), .B2(new_n729), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT34), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT94), .Z(new_n743));
  NOR3_X1   g318(.A1(new_n733), .A2(new_n739), .A3(KEYINPUT34), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n745));
  INV_X1    g320(.A(new_n489), .ZN(new_n746));
  INV_X1    g321(.A(G131), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n489), .A2(KEYINPUT93), .A3(G131), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n751));
  INV_X1    g326(.A(G107), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n751), .B1(new_n481), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n492), .B2(G119), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  MUX2_X1   g330(.A(G25), .B(new_n755), .S(G29), .Z(new_n756));
  XOR2_X1   g331(.A(KEYINPUT35), .B(G1991), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G1986), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n727), .A2(G24), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G290), .B2(G16), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n744), .B(new_n762), .C1(new_n759), .C2(new_n761), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n743), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT36), .ZN(new_n765));
  INV_X1    g340(.A(G29), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G32), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT99), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n493), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n492), .A2(KEYINPUT99), .A3(G129), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT26), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n475), .A2(G105), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n489), .B2(G141), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n767), .B1(new_n779), .B2(new_n766), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT27), .ZN(new_n781));
  INV_X1    g356(.A(G1996), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n766), .A2(G33), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n509), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(new_n473), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n489), .A2(G139), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n784), .B1(new_n792), .B2(new_n766), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2072), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n727), .A2(G19), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n563), .B2(new_n727), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1341), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n727), .A2(G21), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G168), .B2(new_n727), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1966), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n794), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G27), .A2(G29), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G164), .B2(G29), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G2078), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(G2078), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n727), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT23), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n632), .B2(new_n727), .ZN(new_n808));
  INV_X1    g383(.A(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n801), .A2(new_n804), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  AND2_X1   g386(.A1(KEYINPUT24), .A2(G34), .ZN(new_n812));
  NOR2_X1   g387(.A1(KEYINPUT24), .A2(G34), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n766), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT98), .Z(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G160), .B2(G29), .ZN(new_n816));
  INV_X1    g391(.A(G2084), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n727), .A2(G5), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G171), .B2(new_n727), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(G1961), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n628), .A2(new_n727), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G4), .B2(new_n727), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n818), .B(new_n821), .C1(new_n671), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n766), .A2(G35), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G162), .B2(new_n766), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT29), .B(G2090), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n766), .A2(G26), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT28), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n489), .A2(G140), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n492), .A2(G128), .ZN(new_n832));
  NOR2_X1   g407(.A1(G104), .A2(G2105), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT95), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n834), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n830), .B1(new_n837), .B2(new_n766), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT96), .B(G2067), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n823), .A2(new_n671), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT30), .B(G28), .ZN(new_n842));
  OR2_X1    g417(.A1(KEYINPUT31), .A2(G11), .ZN(new_n843));
  NAND2_X1  g418(.A1(KEYINPUT31), .A2(G11), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n842), .A2(new_n766), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n649), .B2(new_n766), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT100), .Z(new_n847));
  NAND4_X1  g422(.A1(new_n828), .A2(new_n840), .A3(new_n841), .A4(new_n847), .ZN(new_n848));
  NOR4_X1   g423(.A1(new_n783), .A2(new_n811), .A3(new_n824), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n765), .A2(new_n849), .ZN(G150));
  INV_X1    g425(.A(G150), .ZN(G311));
  XNOR2_X1  g426(.A(KEYINPUT101), .B(G93), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n553), .A2(new_n852), .B1(new_n527), .B2(G55), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n515), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G860), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n628), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  INV_X1    g437(.A(new_n856), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n563), .A2(new_n863), .A3(new_n853), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n854), .A2(new_n856), .B1(new_n562), .B2(new_n560), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n862), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT102), .Z(new_n869));
  OAI21_X1  g444(.A(new_n858), .B1(new_n867), .B2(KEYINPUT39), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n860), .B1(new_n869), .B2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(KEYINPUT105), .B(G37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n489), .A2(G142), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  INV_X1    g449(.A(G118), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n481), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n492), .B2(G130), .ZN(new_n877));
  INV_X1    g452(.A(new_n643), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n750), .A2(new_n878), .A3(new_n754), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n750), .B2(new_n754), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n873), .B(new_n877), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n877), .A2(new_n873), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n884), .A3(new_n879), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT4), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n488), .A2(new_n503), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(KEYINPUT71), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n890), .A2(new_n507), .B1(new_n504), .B2(new_n512), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n891), .A2(new_n502), .A3(new_n836), .ZN(new_n892));
  NOR2_X1   g467(.A1(G164), .A2(new_n837), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n779), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n508), .A2(new_n513), .ZN(new_n895));
  INV_X1    g470(.A(new_n502), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n836), .ZN(new_n898));
  NAND2_X1  g473(.A1(G164), .A2(new_n837), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n778), .A3(new_n899), .ZN(new_n900));
  AOI211_X1 g475(.A(new_n887), .B(new_n792), .C1(new_n894), .C2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n792), .A2(new_n887), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n792), .A2(new_n887), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n894), .A2(new_n900), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n886), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n495), .A2(new_n649), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n495), .A2(new_n649), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n486), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(G160), .A3(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n894), .A2(new_n900), .A3(new_n904), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n902), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n919), .A2(new_n882), .A3(new_n885), .A4(new_n905), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n907), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n917), .B1(new_n907), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n872), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n925));
  XNOR2_X1  g500(.A(G166), .B(new_n735), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n607), .A2(G305), .A3(new_n608), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(G305), .B1(new_n607), .B2(new_n608), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n930), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n926), .A3(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n925), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n936), .B(KEYINPUT42), .C1(new_n925), .C2(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(KEYINPUT42), .B2(new_n936), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n866), .B(new_n637), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n626), .A2(new_n627), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n618), .A2(KEYINPUT83), .A3(new_n619), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT83), .B1(new_n618), .B2(new_n619), .ZN(new_n943));
  OAI211_X1 g518(.A(G299), .B(new_n941), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n622), .A2(new_n623), .ZN(new_n946));
  AOI21_X1  g521(.A(G299), .B1(new_n946), .B2(new_n941), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n628), .A2(KEYINPUT106), .A3(G299), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n940), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n944), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT41), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n939), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n952), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n939), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n938), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(G868), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(G868), .B2(new_n857), .ZN(G295));
  OAI21_X1  g534(.A(new_n958), .B1(G868), .B2(new_n857), .ZN(G331));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n552), .A2(new_n555), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n552), .B2(new_n555), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n964), .A2(new_n965), .A3(G286), .ZN(new_n966));
  NAND2_X1  g541(.A1(G301), .A2(KEYINPUT109), .ZN(new_n967));
  AOI21_X1  g542(.A(G168), .B1(new_n967), .B2(new_n963), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n866), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(G286), .B1(new_n964), .B2(new_n965), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(G168), .A3(new_n963), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n864), .A2(new_n865), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(KEYINPUT110), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n970), .A2(new_n972), .A3(new_n971), .A4(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n974), .A2(new_n953), .A3(new_n950), .A4(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n969), .A2(new_n973), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n952), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n934), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n977), .A2(new_n979), .ZN(new_n982));
  INV_X1    g557(.A(new_n934), .ZN(new_n983));
  AOI21_X1  g558(.A(G37), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n934), .B1(new_n977), .B2(new_n979), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT111), .B1(new_n987), .B2(G37), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n961), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n978), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n948), .A2(new_n949), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(KEYINPUT41), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n991), .B(KEYINPUT41), .C1(new_n948), .C2(new_n949), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(KEYINPUT41), .B2(new_n955), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n990), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n974), .A2(new_n976), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n952), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n934), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n980), .A2(new_n872), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n999), .A2(KEYINPUT43), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT112), .B1(new_n989), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n982), .A2(new_n983), .ZN(new_n1003));
  INV_X1    g578(.A(G37), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n985), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n988), .A2(new_n1005), .A3(new_n980), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n999), .A2(new_n961), .A3(new_n1000), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n961), .B2(new_n1006), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1011), .B2(new_n1014), .ZN(G397));
  AOI21_X1  g590(.A(KEYINPUT122), .B1(new_n632), .B2(KEYINPUT57), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n573), .A2(new_n572), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT121), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n577), .B2(new_n581), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1017), .A2(KEYINPUT121), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1016), .B1(new_n1021), .B2(KEYINPUT57), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n632), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT45), .B(new_n1026), .C1(new_n891), .C2(new_n502), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(G164), .B2(G1384), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1029), .A3(KEYINPUT115), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n897), .A2(new_n1031), .A3(KEYINPUT45), .A4(new_n1026), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n476), .B(G40), .C1(new_n483), .C2(new_n485), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT56), .B(G2072), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n897), .A2(new_n1038), .A3(new_n1026), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1035), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n809), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1025), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1348), .B1(new_n1044), .B2(new_n1039), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n897), .A2(new_n1026), .A3(new_n1035), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(G2067), .ZN(new_n1048));
  NOR3_X1   g623(.A1(G164), .A2(G1384), .A3(new_n1034), .ZN(new_n1049));
  INV_X1    g624(.A(G2067), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(KEYINPUT123), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1045), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n628), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1037), .A2(new_n1025), .A3(new_n1042), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1043), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT61), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1036), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n1034), .B(new_n1059), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1956), .B1(new_n1044), .B2(new_n1039), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1060), .A2(new_n1024), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1058), .B1(new_n1062), .B2(new_n1043), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1024), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(new_n1056), .A3(KEYINPUT61), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1034), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1067), .A2(new_n782), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT58), .B(G1341), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1049), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT59), .B(new_n563), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1070), .B1(new_n1067), .B2(new_n782), .ZN(new_n1073));
  INV_X1    g648(.A(new_n563), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1054), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1041), .A2(new_n671), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1077), .A2(new_n628), .A3(new_n1051), .A4(new_n1048), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1078), .A2(KEYINPUT60), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1071), .A2(new_n1075), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1057), .B1(new_n1066), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n1084));
  INV_X1    g659(.A(G8), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1049), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1047), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT118), .B(G1981), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n591), .B(new_n1090), .C1(new_n595), .C2(new_n596), .ZN(new_n1091));
  INV_X1    g666(.A(new_n591), .ZN(new_n1092));
  OAI21_X1  g667(.A(G1981), .B1(new_n1092), .B2(new_n594), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT49), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1083), .B1(new_n1088), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g675(.A(KEYINPUT119), .B(new_n1098), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n735), .A2(G1976), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT117), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n735), .B2(G1976), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1088), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1104), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1102), .A2(new_n1111), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1067), .A2(G1971), .B1(G2090), .B2(new_n1041), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G8), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G166), .A2(new_n1085), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT55), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1113), .A2(G8), .A3(new_n1116), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1112), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1027), .A2(new_n1029), .A3(new_n1035), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(G2078), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT124), .B(G1961), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1122), .A2(new_n1124), .B1(new_n1041), .B2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g701(.A(G2078), .B(new_n1034), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1127));
  OAI211_X1 g702(.A(G301), .B(new_n1126), .C1(new_n1127), .C2(KEYINPUT53), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT54), .ZN(new_n1129));
  INV_X1    g704(.A(G2078), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1067), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1123), .ZN(new_n1132));
  AND4_X1   g707(.A1(G40), .A2(new_n476), .A3(new_n482), .A4(new_n1124), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1033), .A2(new_n1133), .B1(new_n1041), .B2(new_n1125), .ZN(new_n1134));
  AOI21_X1  g709(.A(G301), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1120), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1044), .A2(new_n1138), .A3(new_n817), .A4(new_n1039), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT120), .B1(new_n1041), .B2(G2084), .ZN(new_n1140));
  INV_X1    g715(.A(G1966), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1121), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G286), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1139), .A2(new_n1140), .A3(G168), .A4(new_n1142), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(G8), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT51), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(KEYINPUT51), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1132), .A2(new_n1126), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1132), .A2(G301), .A3(new_n1134), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1082), .A2(new_n1137), .A3(new_n1151), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1091), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1049), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT116), .B1(new_n1047), .B2(G8), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1099), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT119), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1088), .A2(new_n1083), .A3(new_n1099), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(G288), .A2(G1976), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1088), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1110), .A2(new_n1106), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1107), .B(new_n1104), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1165), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n1167), .A2(new_n1168), .B1(new_n1172), .B2(new_n1119), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1143), .A2(G8), .A3(G168), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1112), .A2(new_n1118), .A3(new_n1119), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1119), .A2(new_n1171), .A3(new_n1165), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1178), .A2(KEYINPUT63), .A3(new_n1118), .A4(new_n1174), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1173), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT51), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1147), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n1182), .B2(new_n1144), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT62), .B1(new_n1183), .B2(new_n1149), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1120), .A2(new_n1153), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1148), .A2(new_n1150), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1158), .A2(new_n1180), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1029), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1035), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n836), .B(new_n1050), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1193), .A2(KEYINPUT114), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(KEYINPUT114), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1191), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n778), .B(G1996), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1194), .A2(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n750), .A2(new_n757), .A3(new_n754), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n757), .B1(new_n750), .B2(new_n754), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1196), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(G290), .B(G1986), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1202), .B1(new_n1196), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1189), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1191), .B1(new_n779), .B2(new_n1192), .ZN(new_n1206));
  OR3_X1    g781(.A1(new_n1191), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1207));
  OAI21_X1  g782(.A(KEYINPUT46), .B1(new_n1191), .B2(G1996), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT47), .Z(new_n1210));
  NOR3_X1   g785(.A1(new_n1191), .A2(G1986), .A3(G290), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT48), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1210), .B1(new_n1202), .B2(new_n1212), .ZN(new_n1213));
  AOI22_X1  g788(.A1(new_n1198), .A2(new_n1199), .B1(new_n1050), .B2(new_n837), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1214), .A2(KEYINPUT125), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1191), .B1(new_n1214), .B2(KEYINPUT125), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1213), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1205), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n1220));
  NOR2_X1   g794(.A1(G227), .A2(new_n460), .ZN(new_n1221));
  XNOR2_X1  g795(.A(new_n1221), .B(KEYINPUT126), .ZN(new_n1222));
  AND3_X1   g796(.A1(new_n721), .A2(new_n1222), .A3(new_n678), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n923), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g798(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n1220), .B1(new_n1010), .B2(new_n1225), .ZN(new_n1226));
  AOI211_X1 g800(.A(KEYINPUT127), .B(new_n1224), .C1(new_n1002), .C2(new_n1009), .ZN(new_n1227));
  NOR2_X1   g801(.A1(new_n1226), .A2(new_n1227), .ZN(G308));
  NAND2_X1  g802(.A1(new_n1010), .A2(new_n1225), .ZN(G225));
endmodule


