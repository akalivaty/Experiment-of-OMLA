//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265, new_n1266;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT64), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(KEYINPUT64), .B1(new_n207), .B2(new_n208), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n206), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(new_n217), .A2(new_n218), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(new_n218), .B2(new_n217), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n215), .A2(new_n226), .ZN(G361));
  XOR2_X1   g0027(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G226), .B(G232), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n202), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n239), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n251));
  INV_X1    g0051(.A(new_n222), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n255), .B(new_n247), .C1(G41), .C2(G45), .ZN(new_n256));
  AND3_X1   g0056(.A1(new_n251), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n257), .A2(G226), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G222), .ZN(new_n262));
  OR3_X1    g0062(.A1(new_n261), .A2(KEYINPUT67), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT67), .B1(new_n261), .B2(new_n262), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n260), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n270), .A2(G223), .B1(G77), .B2(new_n269), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n263), .A2(new_n264), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n273));
  AOI211_X1 g0073(.A(new_n250), .B(new_n258), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G179), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G50), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n222), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n247), .B2(G20), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n278), .B1(new_n281), .B2(G50), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n265), .A2(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n283), .A2(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(G20), .B2(new_n203), .ZN(new_n290));
  INV_X1    g0090(.A(new_n280), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n282), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n274), .B2(G169), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n276), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n274), .A2(G190), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n292), .B(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT70), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT70), .A2(G200), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n295), .B(new_n296), .C1(new_n274), .C2(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n294), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n277), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n241), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT12), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n284), .A2(G77), .B1(G20), .B2(new_n241), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n202), .B2(new_n288), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(KEYINPUT11), .A3(new_n280), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n281), .A2(G68), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n307), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n309), .A2(new_n280), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(KEYINPUT11), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n250), .B1(new_n257), .B2(G238), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n266), .A2(new_n268), .A3(G226), .A4(new_n260), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G97), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n273), .ZN(new_n320));
  XOR2_X1   g0120(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n315), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n315), .B2(new_n320), .ZN(new_n324));
  OAI21_X1  g0124(.A(G169), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT73), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n315), .A2(new_n320), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n321), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n315), .A2(new_n320), .A3(new_n322), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G169), .A3(new_n327), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n330), .A2(KEYINPUT13), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(KEYINPUT72), .A3(new_n332), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT72), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n330), .A2(new_n339), .A3(KEYINPUT13), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n275), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n314), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n340), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G190), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n314), .B1(new_n333), .B2(G200), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n270), .A2(G238), .B1(G107), .B2(new_n269), .ZN(new_n347));
  INV_X1    g0147(.A(G232), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n261), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n273), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n250), .B1(new_n257), .B2(G244), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n300), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n281), .A2(G77), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT15), .B(G87), .Z(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n356));
  INV_X1    g0156(.A(new_n283), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(KEYINPUT68), .B2(new_n287), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n287), .A2(KEYINPUT68), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n360), .A2(KEYINPUT69), .A3(new_n280), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT69), .B1(new_n360), .B2(new_n280), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n354), .B1(G77), .B2(new_n277), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n350), .A2(new_n351), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n353), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n352), .A2(new_n275), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n368), .A2(new_n363), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n304), .A2(new_n342), .A3(new_n346), .A4(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT7), .B1(new_n269), .B2(new_n223), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n375), .B(G20), .C1(new_n266), .C2(new_n268), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G58), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n241), .ZN(new_n379));
  OAI21_X1  g0179(.A(G20), .B1(new_n379), .B2(new_n201), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n287), .A2(G159), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT16), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n375), .B1(new_n259), .B2(G20), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n267), .A2(G33), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n388));
  OAI211_X1 g0188(.A(KEYINPUT7), .B(new_n223), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n241), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n385), .B1(new_n390), .B2(new_n382), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n384), .A2(new_n391), .A3(new_n280), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n357), .A2(new_n277), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n281), .B2(new_n357), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n266), .A2(new_n268), .A3(G226), .A4(G1698), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n266), .A2(new_n268), .A3(G223), .A4(new_n260), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT74), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT74), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n396), .A2(new_n397), .A3(new_n401), .A4(new_n398), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n402), .A3(new_n273), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n250), .B1(new_n257), .B2(G232), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n275), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n369), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n395), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n395), .A2(KEYINPUT18), .A3(new_n405), .A4(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n392), .A2(new_n394), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n406), .A2(G200), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n403), .A2(G190), .A3(new_n404), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n413), .A2(new_n414), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n415), .A2(new_n392), .A3(new_n394), .A4(new_n416), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n373), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n266), .A2(new_n268), .A3(G257), .A4(new_n260), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n266), .A2(new_n268), .A3(G264), .A4(G1698), .ZN(new_n424));
  INV_X1    g0224(.A(G303), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n423), .B(new_n424), .C1(new_n425), .C2(new_n259), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n273), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n247), .A2(G45), .A3(G274), .ZN(new_n428));
  OR2_X1    g0228(.A1(KEYINPUT5), .A2(G41), .ZN(new_n429));
  NAND2_X1  g0229(.A1(KEYINPUT5), .A2(G41), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT5), .B(G41), .ZN(new_n432));
  INV_X1    g0232(.A(G45), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(G1), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n432), .A2(new_n434), .B1(new_n252), .B2(new_n253), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n431), .B1(new_n435), .B2(G270), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n369), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n277), .A2(G116), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n247), .A2(G33), .ZN(new_n439));
  AND4_X1   g0239(.A1(new_n222), .A2(new_n277), .A3(new_n279), .A4(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n440), .B2(G116), .ZN(new_n441));
  OR2_X1    g0241(.A1(KEYINPUT75), .A2(G97), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT75), .A2(G97), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n265), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(G20), .B1(G33), .B2(G283), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G116), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n279), .A2(new_n222), .B1(G20), .B2(new_n447), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n446), .A2(KEYINPUT20), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT20), .B1(new_n446), .B2(new_n448), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n441), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n437), .A2(new_n451), .A3(KEYINPUT21), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT80), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n437), .A2(new_n451), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT21), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT80), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n437), .A2(new_n451), .A3(new_n457), .A4(KEYINPUT21), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n427), .A2(new_n436), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n275), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n451), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n453), .A2(new_n456), .A3(new_n458), .A4(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n459), .A2(new_n365), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n451), .B(new_n463), .C1(G200), .C2(new_n459), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT6), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT75), .A2(G97), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT75), .A2(G97), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G107), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G97), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n470), .ZN(new_n473));
  NOR2_X1   g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n473), .A2(KEYINPUT6), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT76), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n442), .A2(new_n443), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT6), .B1(new_n477), .B2(G107), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT76), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n474), .A2(KEYINPUT6), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n472), .B2(new_n470), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n476), .A2(new_n482), .A3(G20), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n386), .A2(new_n389), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(G107), .B1(G77), .B2(new_n287), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n291), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n305), .A2(new_n472), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n291), .A2(new_n277), .A3(new_n439), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(new_n472), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT78), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(KEYINPUT77), .B2(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n266), .A2(new_n268), .A3(G244), .A4(new_n260), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n266), .A2(new_n268), .A3(G250), .A4(G1698), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n498), .C1(new_n493), .C2(new_n492), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n273), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n431), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n435), .A2(G257), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n500), .A2(G190), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT79), .ZN(new_n504));
  INV_X1    g0304(.A(new_n492), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(new_n259), .A3(G244), .A4(new_n260), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n495), .A2(new_n497), .A3(new_n506), .A4(new_n498), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n273), .B1(G257), .B2(new_n435), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT79), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(G190), .A4(new_n501), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n490), .A2(new_n504), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n369), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n508), .A2(new_n275), .A3(new_n501), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n514), .B(new_n515), .C1(new_n486), .C2(new_n489), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n259), .A2(G250), .A3(new_n260), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n259), .A2(G257), .A3(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G294), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n273), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n431), .B1(new_n435), .B2(G264), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(G179), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT83), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n522), .A2(KEYINPUT83), .A3(G179), .A4(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n523), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G169), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n470), .A2(G20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n531), .A2(KEYINPUT23), .B1(G20), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g0333(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n534));
  NAND2_X1  g0334(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n534), .A2(new_n531), .A3(KEYINPUT82), .A4(new_n535), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n266), .A2(new_n268), .A3(new_n223), .A4(G87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT22), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT22), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n259), .A2(new_n543), .A3(new_n223), .A4(G87), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n540), .A2(KEYINPUT24), .A3(new_n545), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n280), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n305), .A2(KEYINPUT25), .A3(new_n470), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT25), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n277), .B2(G107), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n440), .A2(G107), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n530), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G250), .B1(new_n433), .B2(G1), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n428), .B1(new_n273), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n266), .A2(new_n268), .A3(G238), .A4(new_n260), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n266), .A2(new_n268), .A3(G244), .A4(G1698), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(new_n532), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n558), .B1(new_n561), .B2(new_n273), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(G169), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n275), .B2(new_n562), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n355), .A2(new_n277), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n477), .B2(new_n285), .ZN(new_n567));
  INV_X1    g0367(.A(G87), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n568), .B(new_n470), .C1(new_n467), .C2(new_n468), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n223), .B1(new_n318), .B2(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n259), .A2(new_n223), .A3(G68), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n565), .B1(new_n573), .B2(new_n280), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n440), .A2(new_n355), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n365), .B(new_n558), .C1(new_n561), .C2(new_n273), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n561), .A2(new_n273), .ZN(new_n578));
  INV_X1    g0378(.A(new_n558), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n300), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n488), .A2(new_n568), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n565), .B(new_n582), .C1(new_n573), .C2(new_n280), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n564), .A2(new_n576), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n528), .A2(G190), .ZN(new_n585));
  AOI21_X1  g0385(.A(G200), .B1(new_n522), .B2(new_n523), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n550), .B(new_n554), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n556), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n422), .A2(new_n465), .A3(new_n517), .A4(new_n588), .ZN(G372));
  NAND2_X1  g0389(.A1(new_n346), .A2(new_n371), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n342), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT86), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n420), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n591), .A2(KEYINPUT86), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n412), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n302), .A2(new_n303), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n294), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT84), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n524), .A2(new_n525), .B1(new_n528), .B2(G169), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n527), .B1(new_n550), .B2(new_n554), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n516), .B(new_n513), .C1(new_n462), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n584), .A2(new_n587), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n602), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n454), .A2(new_n455), .B1(new_n460), .B2(new_n451), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n556), .A2(new_n458), .A3(new_n453), .A4(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n517), .A2(new_n604), .A3(KEYINPUT84), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n563), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n562), .A2(new_n275), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n576), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n490), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n584), .A2(new_n515), .A3(new_n613), .A4(new_n514), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n614), .B2(KEYINPUT26), .ZN(new_n615));
  INV_X1    g0415(.A(new_n580), .ZN(new_n616));
  INV_X1    g0416(.A(new_n582), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n562), .A2(G190), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n616), .A2(new_n574), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT85), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n620), .B1(new_n516), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n613), .A2(KEYINPUT85), .A3(new_n515), .A4(new_n514), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n608), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n422), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n597), .A2(new_n628), .ZN(G369));
  AND2_X1   g0429(.A1(new_n223), .A2(G13), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n247), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G213), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G343), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n451), .ZN(new_n637));
  MUX2_X1   g0437(.A(new_n462), .B(new_n465), .S(new_n637), .Z(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(G330), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n555), .A2(new_n636), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n556), .A2(new_n640), .A3(new_n587), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n600), .A2(new_n636), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n636), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n462), .A2(new_n556), .A3(new_n587), .A4(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n600), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(G399));
  INV_X1    g0448(.A(new_n569), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n447), .ZN(new_n650));
  INV_X1    g0450(.A(new_n216), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(G41), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n650), .A2(new_n247), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n221), .B2(new_n652), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT87), .Z(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT29), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n517), .A2(new_n604), .A3(new_n606), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n516), .A2(new_n620), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n612), .B1(new_n659), .B2(new_n623), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n622), .A2(new_n624), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n658), .B(new_n660), .C1(new_n661), .C2(new_n623), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n657), .B1(new_n662), .B2(new_n645), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n636), .B1(new_n608), .B2(new_n626), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n657), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n578), .A2(new_n579), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n528), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n460), .A3(new_n508), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT30), .ZN(new_n669));
  AND4_X1   g0469(.A1(new_n275), .A2(new_n528), .A3(new_n459), .A4(new_n666), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n668), .A2(new_n669), .B1(new_n670), .B2(new_n511), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  AOI211_X1 g0472(.A(KEYINPUT31), .B(new_n645), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n517), .A2(new_n588), .A3(new_n465), .A4(new_n645), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT31), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n636), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n673), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n665), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n656), .B1(new_n680), .B2(G1), .ZN(G364));
  NOR2_X1   g0481(.A1(new_n223), .A2(G179), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n365), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n300), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G283), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n223), .A2(new_n275), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n365), .A3(G200), .ZN(new_n688));
  XOR2_X1   g0488(.A(KEYINPUT33), .B(G317), .Z(new_n689));
  OAI22_X1  g0489(.A1(new_n685), .A2(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n365), .A2(G200), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n223), .B1(new_n691), .B2(new_n275), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(G294), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(G190), .A2(G200), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n682), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n259), .B1(new_n697), .B2(G329), .ZN(new_n698));
  INV_X1    g0498(.A(G326), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n687), .A2(G190), .A3(G200), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT90), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n687), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT90), .B1(new_n223), .B2(new_n275), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(new_n691), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(G322), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n300), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(G190), .A3(new_n682), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT94), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT94), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n694), .B(new_n707), .C1(new_n713), .C2(new_n425), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n703), .A2(new_n695), .A3(new_n704), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n714), .B1(G311), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n718), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(KEYINPUT92), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n717), .A2(KEYINPUT92), .A3(new_n716), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G77), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n684), .A2(G107), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n726), .B(new_n259), .C1(new_n378), .C2(new_n705), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n697), .A2(G159), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT93), .B(KEYINPUT32), .Z(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n241), .B2(new_n688), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n728), .A2(new_n729), .B1(new_n202), .B2(new_n700), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n727), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n713), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G87), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n692), .A2(KEYINPUT95), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n692), .A2(KEYINPUT95), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G97), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n725), .A2(new_n733), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT96), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n719), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n742), .B2(new_n741), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n222), .B1(G20), .B2(new_n369), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n630), .B(KEYINPUT88), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G45), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G1), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n652), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n651), .A2(new_n269), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n752), .A2(G355), .B1(new_n447), .B2(new_n651), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n245), .A2(new_n433), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n651), .A2(new_n259), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G45), .B2(new_n220), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n745), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n751), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT89), .Z(new_n763));
  NAND2_X1  g0563(.A1(new_n746), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT97), .ZN(new_n765));
  INV_X1    g0565(.A(new_n760), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n638), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n639), .A2(new_n750), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n638), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(G396));
  INV_X1    g0571(.A(new_n371), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n363), .A2(new_n636), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n367), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n371), .A2(new_n645), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n664), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n679), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n664), .A2(new_n776), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(KEYINPUT99), .B1(new_n780), .B2(new_n751), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(KEYINPUT99), .A3(new_n751), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n745), .A2(new_n758), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n688), .ZN(new_n788));
  INV_X1    g0588(.A(new_n700), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n788), .A2(G283), .B1(new_n789), .B2(G303), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n706), .A2(G294), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n684), .A2(G87), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n259), .B1(new_n697), .B2(G311), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n740), .B1(new_n713), .B2(new_n470), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n794), .B(new_n795), .C1(new_n724), .C2(G116), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n706), .A2(G143), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n788), .A2(G150), .B1(new_n789), .B2(G137), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n797), .B(new_n798), .C1(new_n723), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT34), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n259), .B1(new_n696), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G58), .B2(new_n693), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n805), .B1(new_n241), .B2(new_n685), .C1(new_n713), .C2(new_n202), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n800), .B2(new_n801), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n796), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n745), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n750), .B1(G77), .B2(new_n787), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT98), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(new_n759), .C2(new_n776), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n785), .A2(new_n814), .ZN(G384));
  NAND2_X1  g0615(.A1(new_n476), .A2(new_n482), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT35), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n476), .A2(new_n482), .A3(KEYINPUT35), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n818), .A2(G116), .A3(new_n224), .A4(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT36), .Z(new_n821));
  INV_X1    g0621(.A(G77), .ZN(new_n822));
  OR3_X1    g0622(.A1(new_n220), .A2(new_n822), .A3(new_n379), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n247), .B(G13), .C1(new_n823), .C2(new_n240), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT40), .ZN(new_n826));
  INV_X1    g0626(.A(new_n634), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n395), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(KEYINPUT101), .A2(KEYINPUT37), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n408), .A2(new_n828), .A3(new_n418), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(KEYINPUT101), .A2(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n395), .A2(new_n827), .B1(KEYINPUT101), .B2(KEYINPUT37), .ZN(new_n833));
  INV_X1    g0633(.A(new_n831), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n833), .A2(new_n408), .A3(new_n418), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n828), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n421), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT38), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n828), .B1(new_n412), .B2(new_n420), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n832), .A2(new_n835), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n314), .A2(new_n636), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n346), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT100), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n342), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(KEYINPUT100), .B(new_n314), .C1(new_n336), .C2(new_n341), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n343), .A2(G179), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n851), .A2(new_n329), .A3(new_n334), .A4(new_n335), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(new_n314), .A3(new_n636), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n678), .B(new_n776), .C1(new_n850), .C2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n826), .B1(new_n844), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n774), .A2(new_n775), .ZN(new_n857));
  INV_X1    g0657(.A(new_n846), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT100), .B1(new_n852), .B2(new_n314), .ZN(new_n859));
  INV_X1    g0659(.A(new_n849), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n857), .B1(new_n861), .B2(new_n853), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n836), .B(new_n838), .C1(KEYINPUT103), .C2(KEYINPUT38), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n832), .A2(KEYINPUT103), .A3(new_n835), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n842), .B(new_n864), .C1(new_n840), .C2(new_n841), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n862), .A2(new_n866), .A3(KEYINPUT40), .A4(new_n678), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n856), .A2(new_n867), .A3(new_n422), .A4(new_n678), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n856), .A2(G330), .A3(new_n867), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n422), .A2(new_n778), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n868), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n597), .ZN(new_n874));
  INV_X1    g0674(.A(new_n422), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n665), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n873), .B(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n859), .A2(new_n860), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n645), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n863), .A2(new_n881), .A3(new_n865), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n836), .A2(new_n838), .A3(KEYINPUT38), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n842), .B1(new_n840), .B2(new_n841), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT102), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT102), .B1(new_n887), .B2(KEYINPUT39), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n880), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n779), .A2(new_n775), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n850), .A2(new_n854), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n412), .A2(new_n827), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n878), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n247), .B2(new_n747), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n878), .A2(new_n898), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n825), .B1(new_n900), .B2(new_n901), .ZN(G367));
  NOR2_X1   g0702(.A1(new_n583), .A2(new_n645), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n612), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n620), .B2(new_n903), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n517), .B1(new_n490), .B2(new_n645), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n516), .B1(new_n907), .B2(new_n556), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n645), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n646), .A2(new_n517), .A3(new_n606), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT42), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n906), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT104), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n913), .B(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n516), .A2(new_n645), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n907), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n644), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n915), .A2(new_n919), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n652), .B(KEYINPUT41), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n644), .ZN(new_n924));
  INV_X1    g0724(.A(new_n643), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n462), .A2(new_n645), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n646), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n639), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n680), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT105), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n644), .B2(KEYINPUT106), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(KEYINPUT106), .B2(new_n644), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n917), .A2(new_n647), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT45), .Z(new_n936));
  NOR2_X1   g0736(.A1(new_n917), .A2(new_n647), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n931), .A2(new_n934), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n923), .B1(new_n940), .B2(new_n680), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n920), .B(new_n921), .C1(new_n749), .C2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n755), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n235), .A2(new_n943), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n745), .B(new_n760), .C1(new_n651), .C2(new_n355), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n751), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT107), .B1(new_n713), .B2(new_n447), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT46), .Z(new_n948));
  INV_X1    g0748(.A(G317), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n269), .B1(new_n696), .B2(new_n949), .C1(new_n692), .C2(new_n470), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n684), .A2(new_n469), .B1(G294), .B2(new_n788), .ZN(new_n951));
  INV_X1    g0751(.A(G311), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n951), .B1(new_n952), .B2(new_n700), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n950), .B(new_n953), .C1(G303), .C2(new_n706), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n948), .B(new_n954), .C1(new_n686), .C2(new_n723), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT108), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n738), .A2(new_n241), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n734), .B2(G58), .ZN(new_n958));
  INV_X1    g0758(.A(G137), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n259), .B1(new_n696), .B2(new_n959), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n685), .A2(new_n822), .B1(new_n799), .B2(new_n688), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(G143), .C2(new_n789), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n958), .B(new_n962), .C1(new_n286), .C2(new_n705), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G50), .B2(new_n724), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(KEYINPUT47), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n745), .B1(new_n965), .B2(KEYINPUT47), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n946), .B1(new_n766), .B2(new_n905), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n942), .A2(new_n968), .ZN(G387));
  INV_X1    g0769(.A(KEYINPUT112), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n925), .A2(new_n760), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n232), .A2(new_n433), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n972), .A2(new_n755), .B1(new_n650), .B2(new_n752), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT50), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n357), .B2(new_n202), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n283), .A2(KEYINPUT50), .A3(G50), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n433), .B1(new_n241), .B2(new_n822), .ZN(new_n977));
  NOR4_X1   g0777(.A1(new_n650), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n973), .A2(new_n978), .B1(G107), .B2(new_n216), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n751), .B1(new_n979), .B2(new_n761), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n971), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT109), .B(G322), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n952), .A2(new_n688), .B1(new_n700), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G317), .B2(new_n706), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n723), .B2(new_n425), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT110), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT48), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(G294), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n713), .A2(new_n991), .B1(new_n686), .B2(new_n692), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT111), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n988), .A2(new_n989), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT49), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n994), .A2(KEYINPUT49), .A3(new_n995), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n269), .B1(new_n699), .B2(new_n696), .C1(new_n685), .C2(new_n447), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n734), .A2(G77), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n718), .A2(G68), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n259), .B1(new_n696), .B2(new_n286), .C1(new_n700), .C2(new_n799), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n685), .A2(new_n472), .B1(new_n283), .B2(new_n688), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G50), .C2(new_n706), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n739), .A2(new_n355), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n970), .B(new_n982), .C1(new_n1010), .C2(new_n809), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n809), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT112), .B1(new_n1012), .B2(new_n981), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1011), .A2(new_n1013), .B1(new_n749), .B2(new_n929), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n652), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n931), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n680), .B2(new_n929), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1014), .A2(new_n1017), .ZN(G393));
  NOR2_X1   g0818(.A1(new_n239), .A2(new_n943), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n761), .B1(new_n216), .B2(new_n477), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n750), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT113), .Z(new_n1022));
  NOR2_X1   g0822(.A1(new_n738), .A2(new_n822), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n269), .B1(new_n697), .B2(G143), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n792), .B(new_n1024), .C1(new_n202), .C2(new_n688), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(new_n734), .C2(G68), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n705), .A2(new_n799), .B1(new_n286), .B2(new_n700), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT51), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1026), .B(new_n1028), .C1(new_n283), .C2(new_n723), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n447), .A2(new_n692), .B1(new_n688), .B2(new_n425), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n718), .B2(G294), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(KEYINPUT114), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n726), .B(new_n269), .C1(new_n696), .C2(new_n983), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n734), .B2(G283), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(KEYINPUT114), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n705), .A2(new_n952), .B1(new_n949), .B2(new_n700), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT52), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1029), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1022), .B1(new_n1040), .B2(new_n745), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n917), .B2(new_n766), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n939), .B(new_n924), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n749), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n940), .A2(new_n652), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(new_n930), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(G390));
  INV_X1    g0849(.A(new_n775), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n664), .B2(new_n776), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n880), .B1(new_n1051), .B2(new_n892), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n886), .A3(new_n889), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n662), .A2(new_n645), .A3(new_n774), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1054), .A2(new_n775), .B1(new_n861), .B2(new_n853), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n866), .A2(new_n880), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n862), .A2(new_n778), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1053), .A2(new_n1060), .A3(new_n1058), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n597), .B(new_n871), .C1(new_n875), .C2(new_n665), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1054), .A2(new_n775), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT115), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n892), .B1(new_n1067), .B2(new_n857), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n679), .A2(new_n857), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1069), .A2(new_n893), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n891), .B1(new_n1061), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1065), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1015), .B1(new_n1064), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1062), .A2(new_n1074), .A3(new_n1063), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT39), .B1(new_n839), .B2(new_n843), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n863), .A2(new_n881), .A3(new_n865), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n888), .B1(new_n1081), .B2(KEYINPUT102), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1061), .B(new_n1057), .C1(new_n1082), .C2(new_n1052), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1060), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n749), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1082), .A2(new_n758), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n751), .B1(new_n283), .B2(new_n786), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1023), .B1(new_n734), .B2(G87), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n269), .B1(new_n991), .B2(new_n696), .C1(new_n685), .C2(new_n241), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G283), .B2(new_n789), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(new_n447), .C2(new_n705), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n723), .A2(new_n477), .B1(new_n470), .B2(new_n688), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(KEYINPUT116), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(KEYINPUT116), .B2(new_n1093), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n713), .A2(new_n286), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT53), .ZN(new_n1097));
  XOR2_X1   g0897(.A(KEYINPUT54), .B(G143), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n724), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n738), .A2(new_n799), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n685), .A2(new_n202), .B1(new_n1101), .B2(new_n700), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n705), .A2(new_n803), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n269), .B1(new_n697), .B2(G125), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n959), .B2(new_n688), .ZN(new_n1105));
  NOR4_X1   g0905(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1097), .A2(new_n1099), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1095), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1109), .A2(KEYINPUT117), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n745), .B1(new_n1109), .B2(KEYINPUT117), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1087), .B(new_n1088), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1078), .A2(new_n1086), .A3(new_n1112), .ZN(G378));
  INV_X1    g0913(.A(KEYINPUT57), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1065), .B1(new_n1085), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n292), .A2(new_n827), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n304), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n304), .A2(new_n1117), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n870), .B2(KEYINPUT120), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n880), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT102), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1128), .B2(new_n888), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n892), .B1(new_n779), .B2(new_n775), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n895), .B1(new_n1130), .B2(new_n887), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n856), .A2(new_n867), .A3(KEYINPUT120), .A4(G330), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1125), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1132), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n890), .B2(new_n897), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT120), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n869), .A2(new_n1138), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1114), .B1(new_n1116), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1065), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1077), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(KEYINPUT57), .A3(new_n1141), .A4(new_n1135), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n1146), .A3(new_n652), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1135), .A2(new_n1141), .A3(new_n749), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n750), .B1(G50), .B2(new_n787), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n259), .A2(G41), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n685), .A2(new_n378), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G283), .C2(new_n697), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1003), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n788), .A2(G97), .B1(new_n789), .B2(G116), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n470), .B2(new_n705), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n957), .B(new_n1156), .C1(new_n355), .C2(new_n718), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(G41), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G50), .B1(new_n265), .B2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1158), .A2(KEYINPUT58), .B1(new_n1150), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n734), .A2(new_n1098), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT119), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n720), .A2(new_n959), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n738), .A2(new_n286), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n788), .A2(G132), .B1(new_n789), .B2(G125), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n1101), .B2(new_n705), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n684), .A2(G159), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n697), .C2(G124), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1161), .B1(KEYINPUT58), .B2(new_n1158), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1149), .B1(new_n1175), .B2(new_n745), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1124), .B2(new_n759), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1148), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1147), .A2(new_n1179), .ZN(G375));
  NAND2_X1  g0980(.A1(new_n892), .A2(new_n758), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n750), .B1(G68), .B2(new_n787), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n734), .A2(G97), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n269), .B1(new_n696), .B2(new_n425), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n688), .A2(new_n447), .B1(new_n700), .B2(new_n991), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(G77), .C2(new_n684), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n706), .A2(G283), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1183), .A2(new_n1186), .A3(new_n1008), .A4(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n723), .A2(new_n470), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G132), .A2(new_n789), .B1(new_n788), .B2(new_n1098), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n959), .B2(new_n705), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT121), .Z(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n286), .B2(new_n720), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n269), .B(new_n1151), .C1(G128), .C2(new_n697), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n202), .B2(new_n738), .C1(new_n799), .C2(new_n713), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n1188), .A2(new_n1189), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1182), .B1(new_n1196), .B2(new_n745), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1115), .A2(new_n749), .B1(new_n1181), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1075), .A2(new_n922), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1115), .A2(new_n1144), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(G381));
  AND3_X1   g1001(.A1(new_n1147), .A2(KEYINPUT122), .A3(new_n1179), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT122), .B1(new_n1147), .B2(new_n1179), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1202), .A2(new_n1203), .A3(G378), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1014), .A2(new_n770), .A3(new_n1017), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1048), .A2(new_n814), .A3(new_n785), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1205), .A2(G387), .A3(G381), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT123), .ZN(G407));
  INV_X1    g1009(.A(G213), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(G343), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT124), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1210), .B1(new_n1204), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(G407), .A2(new_n1214), .ZN(G409));
  NAND2_X1  g1015(.A1(G387), .A2(new_n1048), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n942), .A2(G390), .A3(new_n968), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1205), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT61), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1216), .A3(new_n1205), .A4(new_n1217), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n785), .A2(KEYINPUT125), .A3(new_n814), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT60), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1115), .B2(new_n1144), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1071), .A2(new_n1065), .A3(new_n1073), .A4(KEYINPUT60), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1227), .A2(new_n652), .A3(new_n1075), .A4(new_n1228), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1225), .A2(new_n1229), .A3(new_n1198), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1198), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(G384), .B(KEYINPUT125), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1230), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1147), .A2(G378), .A3(new_n1179), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1086), .A2(new_n1112), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1116), .A2(new_n1142), .A3(new_n923), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1078), .B(new_n1235), .C1(new_n1236), .C2(new_n1178), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1213), .B(new_n1233), .C1(new_n1234), .C2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1224), .B1(KEYINPUT63), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1233), .A2(G2897), .A3(new_n1213), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1211), .A2(G2897), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(new_n1233), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1211), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT63), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1211), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1233), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1244), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1239), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1213), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1222), .B1(new_n1242), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT62), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1248), .A2(new_n1253), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1254), .A2(KEYINPUT126), .B1(KEYINPUT62), .B2(new_n1238), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1248), .A2(new_n1256), .A3(new_n1253), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1252), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1221), .A2(KEYINPUT127), .A3(new_n1223), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT127), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1250), .B1(new_n1258), .B2(new_n1261), .ZN(G405));
  INV_X1    g1062(.A(new_n1234), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G378), .B1(new_n1147), .B2(new_n1179), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(new_n1247), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1261), .B(new_n1266), .ZN(G402));
endmodule


