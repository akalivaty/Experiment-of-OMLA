

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742;

  INV_X1 U374 ( .A(G953), .ZN(n460) );
  XOR2_X1 U375 ( .A(KEYINPUT67), .B(G101), .Z(n446) );
  XNOR2_X1 U376 ( .A(n535), .B(KEYINPUT33), .ZN(n361) );
  XNOR2_X1 U377 ( .A(n604), .B(n603), .ZN(n610) );
  NOR2_X2 U378 ( .A1(n610), .A2(n609), .ZN(n736) );
  XNOR2_X1 U379 ( .A(n541), .B(KEYINPUT35), .ZN(n640) );
  XOR2_X1 U380 ( .A(G104), .B(G107), .Z(n351) );
  NAND2_X1 U381 ( .A1(n651), .A2(n736), .ZN(n654) );
  XNOR2_X1 U382 ( .A(n508), .B(KEYINPUT1), .ZN(n670) );
  NOR2_X2 U383 ( .A1(n524), .A2(n523), .ZN(n526) );
  XNOR2_X2 U384 ( .A(n494), .B(n493), .ZN(n524) );
  XNOR2_X1 U385 ( .A(n487), .B(n486), .ZN(n533) );
  NAND2_X1 U386 ( .A1(n360), .A2(n368), .ZN(n487) );
  AND2_X1 U387 ( .A1(n367), .A2(n354), .ZN(n360) );
  NOR2_X1 U388 ( .A1(n689), .A2(G953), .ZN(n417) );
  NOR2_X1 U389 ( .A1(G953), .A2(G237), .ZN(n426) );
  XNOR2_X1 U390 ( .A(n456), .B(n455), .ZN(n508) );
  XNOR2_X1 U391 ( .A(n507), .B(KEYINPUT68), .ZN(n671) );
  XNOR2_X1 U392 ( .A(n527), .B(n439), .ZN(n534) );
  XNOR2_X1 U393 ( .A(n434), .B(n362), .ZN(n621) );
  XNOR2_X1 U394 ( .A(n365), .B(n363), .ZN(n362) );
  XNOR2_X1 U395 ( .A(n446), .B(n364), .ZN(n363) );
  AND2_X2 U396 ( .A1(n613), .A2(n612), .ZN(n641) );
  XNOR2_X1 U397 ( .A(n654), .B(KEYINPUT2), .ZN(n613) );
  NAND2_X1 U398 ( .A1(n515), .A2(n353), .ZN(n594) );
  NOR2_X1 U399 ( .A1(n549), .A2(n512), .ZN(n515) );
  NOR2_X1 U400 ( .A1(n449), .A2(G952), .ZN(n649) );
  NOR2_X1 U401 ( .A1(n577), .A2(n742), .ZN(n579) );
  NAND2_X1 U402 ( .A1(n419), .A2(G953), .ZN(n420) );
  INV_X1 U403 ( .A(KEYINPUT5), .ZN(n364) );
  XNOR2_X1 U404 ( .A(n428), .B(n427), .ZN(n365) );
  XOR2_X1 U405 ( .A(n391), .B(KEYINPUT8), .Z(n397) );
  NAND2_X1 U406 ( .A1(n460), .A2(G234), .ZN(n391) );
  XNOR2_X1 U407 ( .A(G113), .B(G104), .ZN(n379) );
  XNOR2_X1 U408 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n462) );
  XNOR2_X1 U409 ( .A(n568), .B(n567), .ZN(n651) );
  XNOR2_X1 U410 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n567) );
  XNOR2_X1 U411 ( .A(n408), .B(n454), .ZN(n611) );
  INV_X1 U412 ( .A(G902), .ZN(n454) );
  XNOR2_X1 U413 ( .A(G119), .B(G116), .ZN(n431) );
  XNOR2_X1 U414 ( .A(KEYINPUT77), .B(G110), .ZN(n447) );
  XNOR2_X1 U415 ( .A(n399), .B(KEYINPUT70), .ZN(n442) );
  INV_X1 U416 ( .A(G137), .ZN(n399) );
  XNOR2_X1 U417 ( .A(G128), .B(G110), .ZN(n400) );
  XNOR2_X1 U418 ( .A(G134), .B(G116), .ZN(n387) );
  NOR2_X1 U419 ( .A1(n518), .A2(n666), .ZN(n519) );
  XNOR2_X1 U420 ( .A(n594), .B(KEYINPUT78), .ZN(n518) );
  OR2_X1 U421 ( .A1(n496), .A2(n534), .ZN(n497) );
  OR2_X1 U422 ( .A1(n670), .A2(n673), .ZN(n495) );
  BUF_X1 U423 ( .A(n533), .Z(n546) );
  NAND2_X1 U424 ( .A1(n366), .A2(n357), .ZN(n367) );
  AND2_X1 U425 ( .A1(n370), .A2(n369), .ZN(n368) );
  INV_X1 U426 ( .A(n480), .ZN(n371) );
  INV_X1 U427 ( .A(n671), .ZN(n510) );
  NAND2_X1 U428 ( .A1(G953), .A2(G224), .ZN(n722) );
  XNOR2_X1 U429 ( .A(n615), .B(n614), .ZN(n616) );
  INV_X1 U430 ( .A(KEYINPUT105), .ZN(n525) );
  AND2_X1 U431 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U432 ( .A1(n733), .A2(G953), .ZN(n734) );
  XNOR2_X1 U433 ( .A(n628), .B(n627), .ZN(n629) );
  AND2_X1 U434 ( .A1(n551), .A2(n550), .ZN(n352) );
  XOR2_X1 U435 ( .A(n514), .B(n513), .Z(n353) );
  OR2_X1 U436 ( .A1(n485), .A2(n484), .ZN(n354) );
  XOR2_X1 U437 ( .A(n595), .B(n539), .Z(n355) );
  OR2_X1 U438 ( .A1(n478), .A2(n660), .ZN(n356) );
  AND2_X1 U439 ( .A1(n663), .A2(n480), .ZN(n357) );
  AND2_X1 U440 ( .A1(n368), .A2(n367), .ZN(n358) );
  XNOR2_X1 U441 ( .A(KEYINPUT62), .B(n621), .ZN(n359) );
  NAND2_X1 U442 ( .A1(n550), .A2(n361), .ZN(n537) );
  AND2_X1 U443 ( .A1(n691), .A2(n361), .ZN(n692) );
  NAND2_X1 U444 ( .A1(n669), .A2(n361), .ZN(n686) );
  INV_X1 U445 ( .A(n478), .ZN(n366) );
  XNOR2_X2 U446 ( .A(n476), .B(n475), .ZN(n478) );
  NAND2_X1 U447 ( .A1(n371), .A2(n660), .ZN(n369) );
  NAND2_X1 U448 ( .A1(n478), .A2(n371), .ZN(n370) );
  INV_X1 U449 ( .A(n508), .ZN(n509) );
  INV_X1 U450 ( .A(n511), .ZN(n512) );
  INV_X1 U451 ( .A(n611), .ZN(n612) );
  INV_X1 U452 ( .A(n649), .ZN(n623) );
  XOR2_X1 U453 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n373) );
  NAND2_X1 U454 ( .A1(G214), .A2(n426), .ZN(n372) );
  XNOR2_X1 U455 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U456 ( .A(n374), .B(KEYINPUT12), .Z(n378) );
  XNOR2_X1 U457 ( .A(G146), .B(G125), .ZN(n463) );
  INV_X1 U458 ( .A(KEYINPUT10), .ZN(n375) );
  XNOR2_X1 U459 ( .A(n375), .B(G140), .ZN(n376) );
  XNOR2_X1 U460 ( .A(n463), .B(n376), .ZN(n729) );
  INV_X1 U461 ( .A(n729), .ZN(n377) );
  XNOR2_X1 U462 ( .A(n378), .B(n377), .ZN(n384) );
  XOR2_X1 U463 ( .A(KEYINPUT99), .B(G122), .Z(n380) );
  XNOR2_X1 U464 ( .A(n380), .B(n379), .ZN(n382) );
  XNOR2_X1 U465 ( .A(G143), .B(G131), .ZN(n381) );
  XNOR2_X1 U466 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U467 ( .A(n384), .B(n383), .ZN(n615) );
  NAND2_X1 U468 ( .A1(n615), .A2(n454), .ZN(n386) );
  XNOR2_X1 U469 ( .A(KEYINPUT13), .B(G475), .ZN(n385) );
  XNOR2_X1 U470 ( .A(n386), .B(n385), .ZN(n553) );
  XOR2_X1 U471 ( .A(G122), .B(G107), .Z(n388) );
  XNOR2_X1 U472 ( .A(n388), .B(n387), .ZN(n390) );
  XNOR2_X2 U473 ( .A(G143), .B(G128), .ZN(n429) );
  XNOR2_X1 U474 ( .A(n429), .B(KEYINPUT101), .ZN(n389) );
  XNOR2_X1 U475 ( .A(n390), .B(n389), .ZN(n395) );
  NAND2_X1 U476 ( .A1(G217), .A2(n397), .ZN(n393) );
  XOR2_X1 U477 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n392) );
  XNOR2_X1 U478 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U479 ( .A(n395), .B(n394), .ZN(n646) );
  NAND2_X1 U480 ( .A1(n646), .A2(n454), .ZN(n396) );
  XNOR2_X1 U481 ( .A(n396), .B(G478), .ZN(n552) );
  OR2_X1 U482 ( .A1(n553), .A2(n552), .ZN(n699) );
  NAND2_X1 U483 ( .A1(G221), .A2(n397), .ZN(n398) );
  XNOR2_X1 U484 ( .A(n398), .B(n729), .ZN(n406) );
  XNOR2_X1 U485 ( .A(n400), .B(n442), .ZN(n404) );
  XOR2_X1 U486 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n402) );
  XNOR2_X1 U487 ( .A(G119), .B(KEYINPUT94), .ZN(n401) );
  XNOR2_X1 U488 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U489 ( .A(n404), .B(n403), .Z(n405) );
  XNOR2_X1 U490 ( .A(n406), .B(n405), .ZN(n643) );
  NOR2_X1 U491 ( .A1(n643), .A2(G902), .ZN(n407) );
  XNOR2_X1 U492 ( .A(n407), .B(KEYINPUT96), .ZN(n413) );
  XOR2_X1 U493 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n410) );
  XNOR2_X1 U494 ( .A(KEYINPUT89), .B(KEYINPUT15), .ZN(n408) );
  NAND2_X1 U495 ( .A1(G234), .A2(n611), .ZN(n409) );
  XNOR2_X1 U496 ( .A(n410), .B(n409), .ZN(n422) );
  NAND2_X1 U497 ( .A1(n422), .A2(G217), .ZN(n411) );
  XNOR2_X1 U498 ( .A(KEYINPUT25), .B(n411), .ZN(n412) );
  XNOR2_X1 U499 ( .A(n413), .B(n412), .ZN(n506) );
  INV_X1 U500 ( .A(n506), .ZN(n414) );
  INV_X1 U501 ( .A(n414), .ZN(n673) );
  XOR2_X1 U502 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n416) );
  NAND2_X1 U503 ( .A1(G234), .A2(G237), .ZN(n415) );
  XNOR2_X1 U504 ( .A(n416), .B(n415), .ZN(n418) );
  NAND2_X1 U505 ( .A1(G952), .A2(n418), .ZN(n689) );
  XNOR2_X1 U506 ( .A(n417), .B(KEYINPUT92), .ZN(n485) );
  INV_X1 U507 ( .A(n485), .ZN(n421) );
  NAND2_X1 U508 ( .A1(G902), .A2(n418), .ZN(n481) );
  NOR2_X1 U509 ( .A1(G900), .A2(n481), .ZN(n419) );
  NAND2_X1 U510 ( .A1(n421), .A2(n420), .ZN(n511) );
  AND2_X1 U511 ( .A1(n422), .A2(G221), .ZN(n424) );
  INV_X1 U512 ( .A(KEYINPUT21), .ZN(n423) );
  XNOR2_X1 U513 ( .A(n424), .B(n423), .ZN(n489) );
  INV_X1 U514 ( .A(n489), .ZN(n674) );
  NAND2_X1 U515 ( .A1(n511), .A2(n674), .ZN(n425) );
  NOR2_X1 U516 ( .A1(n673), .A2(n425), .ZN(n569) );
  NAND2_X1 U517 ( .A1(n426), .A2(G210), .ZN(n428) );
  XOR2_X1 U518 ( .A(G137), .B(G146), .Z(n427) );
  XNOR2_X1 U519 ( .A(n429), .B(KEYINPUT4), .ZN(n465) );
  XNOR2_X1 U520 ( .A(G134), .B(G131), .ZN(n430) );
  XNOR2_X1 U521 ( .A(n465), .B(n430), .ZN(n444) );
  XNOR2_X1 U522 ( .A(n431), .B(KEYINPUT3), .ZN(n433) );
  XNOR2_X1 U523 ( .A(G113), .B(KEYINPUT71), .ZN(n432) );
  XNOR2_X1 U524 ( .A(n433), .B(n432), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n444), .B(n470), .ZN(n434) );
  NAND2_X1 U526 ( .A1(n621), .A2(n454), .ZN(n437) );
  INV_X1 U527 ( .A(KEYINPUT97), .ZN(n435) );
  XNOR2_X1 U528 ( .A(n435), .B(G472), .ZN(n436) );
  XNOR2_X1 U529 ( .A(n437), .B(n436), .ZN(n438) );
  BUF_X2 U530 ( .A(n438), .Z(n527) );
  INV_X1 U531 ( .A(KEYINPUT6), .ZN(n439) );
  NAND2_X1 U532 ( .A1(n569), .A2(n534), .ZN(n440) );
  NOR2_X1 U533 ( .A1(n699), .A2(n440), .ZN(n580) );
  INV_X1 U534 ( .A(G237), .ZN(n441) );
  NAND2_X1 U535 ( .A1(n454), .A2(n441), .ZN(n472) );
  NAND2_X1 U536 ( .A1(n472), .A2(G214), .ZN(n663) );
  NAND2_X1 U537 ( .A1(n580), .A2(n663), .ZN(n457) );
  INV_X1 U538 ( .A(n442), .ZN(n443) );
  XNOR2_X1 U539 ( .A(n444), .B(n443), .ZN(n730) );
  INV_X1 U540 ( .A(KEYINPUT72), .ZN(n445) );
  XNOR2_X1 U541 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U542 ( .A(n351), .B(n447), .ZN(n717) );
  XNOR2_X1 U543 ( .A(n448), .B(n717), .ZN(n459) );
  BUF_X1 U544 ( .A(n460), .Z(n449) );
  NAND2_X1 U545 ( .A1(G227), .A2(n449), .ZN(n451) );
  XOR2_X1 U546 ( .A(G146), .B(G140), .Z(n450) );
  XNOR2_X1 U547 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U548 ( .A(n459), .B(n452), .ZN(n453) );
  XNOR2_X1 U549 ( .A(n730), .B(n453), .ZN(n628) );
  NAND2_X1 U550 ( .A1(n628), .A2(n454), .ZN(n456) );
  INV_X1 U551 ( .A(G469), .ZN(n455) );
  INV_X1 U552 ( .A(n670), .ZN(n523) );
  NOR2_X1 U553 ( .A1(n457), .A2(n523), .ZN(n458) );
  XOR2_X1 U554 ( .A(KEYINPUT43), .B(n458), .Z(n477) );
  INV_X1 U555 ( .A(n459), .ZN(n468) );
  NAND2_X1 U556 ( .A1(n460), .A2(G224), .ZN(n461) );
  XNOR2_X1 U557 ( .A(n462), .B(n461), .ZN(n464) );
  XNOR2_X1 U558 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U559 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U560 ( .A(n468), .B(n467), .ZN(n471) );
  XNOR2_X1 U561 ( .A(KEYINPUT16), .B(G122), .ZN(n469) );
  XNOR2_X1 U562 ( .A(n470), .B(n469), .ZN(n719) );
  XNOR2_X1 U563 ( .A(n471), .B(n719), .ZN(n633) );
  NAND2_X1 U564 ( .A1(n633), .A2(n611), .ZN(n476) );
  NAND2_X1 U565 ( .A1(n472), .A2(G210), .ZN(n474) );
  XNOR2_X1 U566 ( .A(KEYINPUT82), .B(KEYINPUT90), .ZN(n473) );
  XNOR2_X1 U567 ( .A(n474), .B(n473), .ZN(n475) );
  BUF_X1 U568 ( .A(n478), .Z(n596) );
  NAND2_X1 U569 ( .A1(n477), .A2(n596), .ZN(n608) );
  XNOR2_X1 U570 ( .A(n608), .B(G140), .ZN(G42) );
  INV_X1 U571 ( .A(n663), .ZN(n660) );
  INV_X1 U572 ( .A(KEYINPUT66), .ZN(n479) );
  XOR2_X1 U573 ( .A(n479), .B(KEYINPUT19), .Z(n480) );
  INV_X1 U574 ( .A(n481), .ZN(n482) );
  NOR2_X1 U575 ( .A1(G898), .A2(n449), .ZN(n720) );
  NAND2_X1 U576 ( .A1(n482), .A2(n720), .ZN(n483) );
  XNOR2_X1 U577 ( .A(n483), .B(KEYINPUT93), .ZN(n484) );
  XNOR2_X1 U578 ( .A(KEYINPUT88), .B(KEYINPUT0), .ZN(n486) );
  INV_X1 U579 ( .A(n533), .ZN(n492) );
  INV_X1 U580 ( .A(n552), .ZN(n488) );
  AND2_X1 U581 ( .A1(n553), .A2(n488), .ZN(n661) );
  INV_X1 U582 ( .A(n661), .ZN(n490) );
  NOR2_X1 U583 ( .A1(n490), .A2(n489), .ZN(n491) );
  NAND2_X1 U584 ( .A1(n492), .A2(n491), .ZN(n494) );
  XNOR2_X1 U585 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n493) );
  XNOR2_X1 U586 ( .A(n495), .B(KEYINPUT104), .ZN(n496) );
  OR2_X2 U587 ( .A1(n524), .A2(n497), .ZN(n500) );
  INV_X1 U588 ( .A(KEYINPUT81), .ZN(n498) );
  XNOR2_X1 U589 ( .A(n498), .B(KEYINPUT32), .ZN(n499) );
  XNOR2_X2 U590 ( .A(n500), .B(n499), .ZN(n530) );
  XOR2_X1 U591 ( .A(G119), .B(KEYINPUT127), .Z(n501) );
  XNOR2_X1 U592 ( .A(n530), .B(n501), .ZN(G21) );
  OR2_X1 U593 ( .A1(n524), .A2(n523), .ZN(n504) );
  INV_X1 U594 ( .A(n534), .ZN(n502) );
  NAND2_X1 U595 ( .A1(n502), .A2(n673), .ZN(n503) );
  NOR2_X1 U596 ( .A1(n504), .A2(n503), .ZN(n505) );
  XOR2_X1 U597 ( .A(KEYINPUT103), .B(n505), .Z(n557) );
  XOR2_X1 U598 ( .A(G101), .B(n557), .Z(G3) );
  NAND2_X1 U599 ( .A1(n506), .A2(n674), .ZN(n507) );
  NAND2_X1 U600 ( .A1(n510), .A2(n509), .ZN(n549) );
  XNOR2_X1 U601 ( .A(KEYINPUT30), .B(KEYINPUT106), .ZN(n514) );
  NAND2_X1 U602 ( .A1(n527), .A2(n663), .ZN(n513) );
  INV_X1 U603 ( .A(KEYINPUT76), .ZN(n516) );
  XNOR2_X1 U604 ( .A(n516), .B(KEYINPUT38), .ZN(n517) );
  XNOR2_X1 U605 ( .A(n596), .B(n517), .ZN(n666) );
  XNOR2_X1 U606 ( .A(n519), .B(KEYINPUT39), .ZN(n605) );
  NOR2_X1 U607 ( .A1(n605), .A2(n699), .ZN(n522) );
  XNOR2_X1 U608 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n520) );
  XOR2_X1 U609 ( .A(n520), .B(KEYINPUT110), .Z(n521) );
  XNOR2_X1 U610 ( .A(n522), .B(n521), .ZN(n577) );
  XOR2_X1 U611 ( .A(G131), .B(n577), .Z(G33) );
  XNOR2_X1 U612 ( .A(n526), .B(n525), .ZN(n529) );
  NOR2_X1 U613 ( .A1(n673), .A2(n527), .ZN(n528) );
  NAND2_X1 U614 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U615 ( .A(n531), .B(G110), .ZN(G12) );
  INV_X1 U616 ( .A(KEYINPUT73), .ZN(n544) );
  NAND2_X1 U617 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U618 ( .A(n532), .B(KEYINPUT86), .ZN(n563) );
  INV_X1 U619 ( .A(n546), .ZN(n550) );
  NOR2_X1 U620 ( .A1(n671), .A2(n670), .ZN(n545) );
  NAND2_X1 U621 ( .A1(n545), .A2(n534), .ZN(n535) );
  XOR2_X1 U622 ( .A(KEYINPUT80), .B(KEYINPUT34), .Z(n536) );
  XNOR2_X1 U623 ( .A(n537), .B(n536), .ZN(n540) );
  INV_X1 U624 ( .A(n553), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n538), .A2(n552), .ZN(n595) );
  INV_X1 U626 ( .A(KEYINPUT79), .ZN(n539) );
  NAND2_X1 U627 ( .A1(n540), .A2(n355), .ZN(n541) );
  OR2_X2 U628 ( .A1(n640), .A2(KEYINPUT44), .ZN(n542) );
  NOR2_X1 U629 ( .A1(n563), .A2(n542), .ZN(n543) );
  XNOR2_X1 U630 ( .A(n544), .B(n543), .ZN(n562) );
  NAND2_X1 U631 ( .A1(n545), .A2(n527), .ZN(n680) );
  NOR2_X1 U632 ( .A1(n680), .A2(n546), .ZN(n548) );
  XOR2_X1 U633 ( .A(KEYINPUT31), .B(KEYINPUT98), .Z(n547) );
  XNOR2_X1 U634 ( .A(n548), .B(n547), .ZN(n712) );
  NOR2_X1 U635 ( .A1(n549), .A2(n527), .ZN(n551) );
  NOR2_X1 U636 ( .A1(n712), .A2(n352), .ZN(n555) );
  AND2_X1 U637 ( .A1(n553), .A2(n552), .ZN(n711) );
  INV_X1 U638 ( .A(n711), .ZN(n606) );
  NAND2_X1 U639 ( .A1(n606), .A2(n699), .ZN(n664) );
  INV_X1 U640 ( .A(n664), .ZN(n554) );
  NOR2_X1 U641 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U642 ( .A(n556), .B(KEYINPUT102), .ZN(n558) );
  NOR2_X1 U643 ( .A1(n558), .A2(n557), .ZN(n560) );
  NAND2_X1 U644 ( .A1(n640), .A2(KEYINPUT44), .ZN(n559) );
  NAND2_X1 U645 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U646 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U647 ( .A1(n563), .A2(KEYINPUT44), .ZN(n564) );
  XOR2_X1 U648 ( .A(n564), .B(KEYINPUT65), .Z(n565) );
  NAND2_X1 U649 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U650 ( .A(n509), .B(KEYINPUT108), .ZN(n572) );
  NAND2_X1 U651 ( .A1(n527), .A2(n569), .ZN(n570) );
  XOR2_X1 U652 ( .A(KEYINPUT28), .B(n570), .Z(n571) );
  NAND2_X1 U653 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U654 ( .A(n573), .B(KEYINPUT109), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n661), .A2(n663), .ZN(n574) );
  OR2_X1 U656 ( .A1(n666), .A2(n574), .ZN(n575) );
  XNOR2_X1 U657 ( .A(n575), .B(KEYINPUT41), .ZN(n691) );
  NAND2_X1 U658 ( .A1(n585), .A2(n691), .ZN(n576) );
  XOR2_X1 U659 ( .A(n576), .B(KEYINPUT42), .Z(n742) );
  XOR2_X1 U660 ( .A(KEYINPUT85), .B(KEYINPUT46), .Z(n578) );
  XNOR2_X1 U661 ( .A(n579), .B(n578), .ZN(n602) );
  XOR2_X1 U662 ( .A(KEYINPUT112), .B(n580), .Z(n581) );
  NOR2_X1 U663 ( .A1(n581), .A2(n356), .ZN(n582) );
  XOR2_X1 U664 ( .A(KEYINPUT36), .B(n582), .Z(n583) );
  NOR2_X1 U665 ( .A1(n583), .A2(n670), .ZN(n714) );
  XOR2_X1 U666 ( .A(KEYINPUT47), .B(KEYINPUT69), .Z(n586) );
  AND2_X1 U667 ( .A1(n586), .A2(KEYINPUT75), .ZN(n584) );
  NOR2_X1 U668 ( .A1(n714), .A2(n584), .ZN(n593) );
  AND2_X1 U669 ( .A1(n585), .A2(n358), .ZN(n706) );
  NAND2_X1 U670 ( .A1(n706), .A2(n664), .ZN(n589) );
  NOR2_X1 U671 ( .A1(n586), .A2(KEYINPUT75), .ZN(n587) );
  OR2_X1 U672 ( .A1(n589), .A2(n587), .ZN(n591) );
  NOR2_X1 U673 ( .A1(KEYINPUT75), .A2(KEYINPUT47), .ZN(n588) );
  NAND2_X1 U674 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U675 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U676 ( .A1(n593), .A2(n592), .ZN(n600) );
  XOR2_X1 U677 ( .A(KEYINPUT78), .B(n594), .Z(n598) );
  NOR2_X1 U678 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U680 ( .A(n599), .B(KEYINPUT107), .ZN(n741) );
  NOR2_X1 U681 ( .A1(n600), .A2(n741), .ZN(n601) );
  NAND2_X1 U682 ( .A1(n602), .A2(n601), .ZN(n604) );
  XNOR2_X1 U683 ( .A(KEYINPUT84), .B(KEYINPUT48), .ZN(n603) );
  NOR2_X1 U684 ( .A1(n605), .A2(n606), .ZN(n607) );
  XNOR2_X1 U685 ( .A(n607), .B(KEYINPUT113), .ZN(n740) );
  NAND2_X1 U686 ( .A1(n740), .A2(n608), .ZN(n609) );
  INV_X1 U687 ( .A(KEYINPUT2), .ZN(n655) );
  NAND2_X1 U688 ( .A1(n641), .A2(G475), .ZN(n617) );
  XOR2_X1 U689 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n614) );
  XNOR2_X1 U690 ( .A(n617), .B(n616), .ZN(n618) );
  NOR2_X2 U691 ( .A1(n618), .A2(n649), .ZN(n620) );
  XNOR2_X1 U692 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n620), .B(n619), .ZN(G60) );
  NAND2_X1 U694 ( .A1(n641), .A2(G472), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(n359), .ZN(n624) );
  XNOR2_X1 U696 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n626), .B(n625), .ZN(G57) );
  NAND2_X1 U698 ( .A1(n641), .A2(G469), .ZN(n630) );
  XNOR2_X1 U699 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X2 U701 ( .A1(n631), .A2(n649), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n632), .B(KEYINPUT120), .ZN(G54) );
  NAND2_X1 U703 ( .A1(n641), .A2(G210), .ZN(n637) );
  BUF_X1 U704 ( .A(n633), .Z(n634) );
  XNOR2_X1 U705 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n634), .B(n635), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X2 U708 ( .A1(n638), .A2(n649), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U710 ( .A(G122), .B(n640), .Z(G24) );
  BUF_X1 U711 ( .A(n641), .Z(n642) );
  NAND2_X1 U712 ( .A1(n642), .A2(G217), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X1 U714 ( .A1(n645), .A2(n649), .ZN(G66) );
  NAND2_X1 U715 ( .A1(n642), .A2(G478), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n646), .B(KEYINPUT123), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n650), .A2(n649), .ZN(G63) );
  BUF_X1 U719 ( .A(n651), .Z(n652) );
  NOR2_X1 U720 ( .A1(n652), .A2(KEYINPUT2), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n653), .B(KEYINPUT83), .ZN(n659) );
  NAND2_X1 U722 ( .A1(n654), .A2(KEYINPUT2), .ZN(n657) );
  NAND2_X1 U723 ( .A1(n736), .A2(n655), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  AND2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n697) );
  NAND2_X1 U726 ( .A1(n666), .A2(n660), .ZN(n662) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n668) );
  NAND2_X1 U728 ( .A1(n664), .A2(n663), .ZN(n665) );
  OR2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U730 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U731 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U732 ( .A(KEYINPUT50), .B(n672), .ZN(n678) );
  NOR2_X1 U733 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U734 ( .A(KEYINPUT49), .B(n675), .Z(n676) );
  NOR2_X1 U735 ( .A1(n438), .A2(n676), .ZN(n677) );
  NAND2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U737 ( .A(n679), .B(KEYINPUT116), .ZN(n681) );
  NAND2_X1 U738 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U739 ( .A(n682), .B(KEYINPUT51), .ZN(n683) );
  XNOR2_X1 U740 ( .A(n683), .B(KEYINPUT117), .ZN(n684) );
  NAND2_X1 U741 ( .A1(n684), .A2(n691), .ZN(n685) );
  NAND2_X1 U742 ( .A1(n686), .A2(n685), .ZN(n688) );
  XOR2_X1 U743 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n687) );
  XNOR2_X1 U744 ( .A(n688), .B(n687), .ZN(n690) );
  NOR2_X1 U745 ( .A1(n690), .A2(n689), .ZN(n693) );
  OR2_X1 U746 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U747 ( .A(n694), .B(KEYINPUT119), .ZN(n695) );
  NAND2_X1 U748 ( .A1(n695), .A2(n449), .ZN(n696) );
  NOR2_X1 U749 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U750 ( .A(n698), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U751 ( .A(n699), .ZN(n708) );
  NAND2_X1 U752 ( .A1(n352), .A2(n708), .ZN(n700) );
  XNOR2_X1 U753 ( .A(n700), .B(G104), .ZN(G6) );
  XOR2_X1 U754 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n702) );
  NAND2_X1 U755 ( .A1(n352), .A2(n711), .ZN(n701) );
  XNOR2_X1 U756 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U757 ( .A(G107), .B(n703), .ZN(G9) );
  XOR2_X1 U758 ( .A(G128), .B(KEYINPUT29), .Z(n705) );
  NAND2_X1 U759 ( .A1(n706), .A2(n711), .ZN(n704) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(G30) );
  NAND2_X1 U761 ( .A1(n706), .A2(n708), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n707), .B(G146), .ZN(G48) );
  NAND2_X1 U763 ( .A1(n712), .A2(n708), .ZN(n709) );
  XNOR2_X1 U764 ( .A(n709), .B(KEYINPUT114), .ZN(n710) );
  XNOR2_X1 U765 ( .A(G113), .B(n710), .ZN(G15) );
  NAND2_X1 U766 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U767 ( .A(n713), .B(G116), .ZN(G18) );
  XOR2_X1 U768 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n716) );
  XNOR2_X1 U769 ( .A(G125), .B(n714), .ZN(n715) );
  XNOR2_X1 U770 ( .A(n716), .B(n715), .ZN(G27) );
  XOR2_X1 U771 ( .A(G101), .B(n717), .Z(n718) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n721) );
  NOR2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n728) );
  NAND2_X1 U774 ( .A1(n652), .A2(n449), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n722), .B(KEYINPUT124), .ZN(n723) );
  XNOR2_X1 U776 ( .A(KEYINPUT61), .B(n723), .ZN(n724) );
  NAND2_X1 U777 ( .A1(G898), .A2(n724), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(G69) );
  XOR2_X1 U780 ( .A(n730), .B(n729), .Z(n731) );
  XOR2_X1 U781 ( .A(KEYINPUT125), .B(n731), .Z(n735) );
  XOR2_X1 U782 ( .A(G227), .B(n735), .Z(n732) );
  NAND2_X1 U783 ( .A1(n732), .A2(G900), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n734), .B(KEYINPUT126), .ZN(n739) );
  XNOR2_X1 U785 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n737), .A2(n449), .ZN(n738) );
  NAND2_X1 U787 ( .A1(n739), .A2(n738), .ZN(G72) );
  XNOR2_X1 U788 ( .A(G134), .B(n740), .ZN(G36) );
  XOR2_X1 U789 ( .A(G143), .B(n741), .Z(G45) );
  XOR2_X1 U790 ( .A(G137), .B(n742), .Z(G39) );
endmodule

