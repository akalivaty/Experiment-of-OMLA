//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n573, new_n574,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n467), .A2(KEYINPUT71), .A3(G137), .A4(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(KEYINPUT3), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n462), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n472), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n466), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G101), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n462), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n486), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n487), .A2(new_n470), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G160));
  INV_X1    g065(.A(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n467), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G136), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n478), .A2(new_n470), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G124), .ZN(new_n496));
  OAI221_X1 g071(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n468), .A2(new_n469), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n501), .A2(new_n486), .A3(KEYINPUT74), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n504));
  INV_X1    g079(.A(new_n469), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(G138), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n462), .A2(new_n485), .A3(new_n502), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n501), .A2(new_n511), .A3(new_n477), .A4(new_n462), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT4), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n467), .B2(new_n501), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(G126), .A2(G2105), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n477), .A2(new_n462), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  OR2_X1    g093(.A1(G102), .A2(G2105), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n519), .B(G2104), .C1(G114), .C2(new_n491), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n518), .B1(new_n517), .B2(new_n520), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G164));
  AND2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G50), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT75), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT5), .B(G543), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n526), .A2(new_n527), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n534), .ZN(new_n537));
  INV_X1    g112(.A(G88), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n533), .A2(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n532), .A2(new_n539), .ZN(G303));
  INV_X1    g115(.A(G303), .ZN(G166));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT77), .Z(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT76), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT7), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g122(.A1(G63), .A2(G651), .ZN(new_n548));
  INV_X1    g123(.A(G89), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n528), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(new_n534), .B1(new_n530), .B2(G51), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  NAND2_X1  g128(.A1(new_n534), .A2(G64), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n533), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(KEYINPUT78), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(KEYINPUT78), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT5), .B(G543), .Z(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n528), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G90), .B1(new_n530), .B2(G52), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(G301));
  INV_X1    g137(.A(G301), .ZN(G171));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n536), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G81), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n564), .A2(new_n565), .B1(new_n537), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n533), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(new_n530), .A2(G53), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT9), .Z(new_n577));
  NAND2_X1  g152(.A1(new_n560), .A2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  XOR2_X1   g154(.A(new_n579), .B(KEYINPUT79), .Z(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(G65), .B2(new_n534), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n578), .B1(new_n581), .B2(new_n533), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n577), .A2(new_n582), .ZN(G299));
  OAI21_X1  g158(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT80), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n560), .A2(G87), .B1(new_n530), .B2(G49), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G288));
  INV_X1    g163(.A(G48), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n589), .A2(new_n565), .B1(new_n537), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n534), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n533), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n559), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n533), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n599), .B2(new_n598), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n560), .A2(G85), .B1(new_n530), .B2(G47), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n560), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT10), .Z(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n559), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(new_n530), .B2(G54), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G868), .ZN(G284));
  XNOR2_X1  g187(.A(G284), .B(KEYINPUT82), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n577), .A2(new_n582), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n570), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n482), .A2(new_n486), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT83), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n493), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n495), .A2(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n626), .A2(new_n627), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n629), .B(new_n636), .C1(new_n630), .C2(new_n635), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(G14), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n648), .ZN(G401));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(new_n627), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n630), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT85), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n668), .A2(new_n670), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n673), .A3(new_n671), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n678), .C1(new_n673), .C2(new_n677), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  NAND2_X1  g261(.A1(new_n482), .A2(G105), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT98), .ZN(new_n688));
  INV_X1    g263(.A(G141), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n492), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n495), .A2(G129), .ZN(new_n691));
  NAND3_X1  g266(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT26), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n696), .B2(G32), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT27), .B(G1996), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(G33), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT25), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(KEYINPUT97), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(new_n470), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(KEYINPUT97), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI211_X1 g283(.A(new_n703), .B(new_n708), .C1(G139), .C2(new_n493), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n701), .B1(new_n709), .B2(new_n696), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n700), .B1(G2072), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G20), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT23), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n615), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1956), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n698), .B2(new_n699), .ZN(new_n717));
  INV_X1    g292(.A(G2078), .ZN(new_n718));
  NOR2_X1   g293(.A1(G164), .A2(new_n696), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G27), .B2(new_n696), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n711), .B(new_n717), .C1(new_n718), .C2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n718), .B2(new_n720), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT96), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n696), .A2(G26), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n493), .A2(G140), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n495), .A2(G128), .ZN(new_n728));
  OAI221_X1 g303(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n726), .B1(new_n731), .B2(new_n696), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n634), .A2(new_n696), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT31), .B(G11), .Z(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT99), .B(G28), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n736), .B2(KEYINPUT30), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT100), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(KEYINPUT30), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n737), .B2(new_n738), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n735), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n570), .A2(G16), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G16), .B2(G19), .ZN(new_n744));
  INV_X1    g319(.A(G1341), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n734), .B(new_n746), .C1(new_n745), .C2(new_n744), .ZN(new_n747));
  AND2_X1   g322(.A1(KEYINPUT24), .A2(G34), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n696), .B1(KEYINPUT24), .B2(G34), .ZN(new_n749));
  OAI22_X1  g324(.A1(G160), .A2(new_n696), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n747), .B1(G2084), .B2(new_n750), .C1(G2072), .C2(new_n710), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n733), .B(new_n751), .C1(G2084), .C2(new_n750), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n712), .A2(G4), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n611), .B2(new_n712), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT94), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT93), .B(G1348), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n712), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n712), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1966), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G35), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G162), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT29), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2090), .ZN(new_n765));
  NOR2_X1   g340(.A1(G5), .A2(G16), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT101), .Z(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G301), .B2(new_n712), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT102), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n722), .A2(new_n752), .A3(new_n761), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G6), .A2(G16), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n594), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n775), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(G166), .A2(G16), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G16), .B2(G22), .ZN(new_n781));
  INV_X1    g356(.A(G1971), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n782), .B2(new_n781), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n712), .A2(G23), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n587), .B2(new_n712), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT91), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT33), .B(G1976), .Z(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n787), .A2(new_n789), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n784), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT92), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n495), .A2(G119), .ZN(new_n796));
  NOR2_X1   g371(.A1(G95), .A2(G2105), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT86), .Z(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n799));
  INV_X1    g374(.A(G131), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n796), .B(new_n799), .C1(new_n800), .C2(new_n492), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT87), .Z(new_n802));
  MUX2_X1   g377(.A(G25), .B(new_n802), .S(G29), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT88), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G24), .B(G290), .S(G16), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1986), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n795), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n794), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT36), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n794), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n773), .B1(new_n811), .B2(new_n813), .ZN(G311));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n813), .ZN(new_n815));
  INV_X1    g390(.A(new_n773), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(G150));
  INV_X1    g392(.A(G55), .ZN(new_n818));
  INV_X1    g393(.A(G93), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n818), .A2(new_n565), .B1(new_n537), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n533), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT104), .B(G860), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT37), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n606), .A2(new_n610), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n618), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  OR3_X1    g404(.A1(new_n820), .A2(KEYINPUT103), .A3(new_n822), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT103), .B1(new_n820), .B2(new_n822), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n570), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n830), .A2(new_n570), .A3(new_n831), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n829), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n824), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n826), .B1(new_n839), .B2(new_n841), .ZN(G145));
  NAND2_X1  g417(.A1(new_n493), .A2(G142), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT107), .Z(new_n844));
  OAI221_X1 g419(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n470), .C2(G118), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n495), .A2(G130), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n801), .B(new_n625), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n847), .B(new_n848), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT106), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n515), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n517), .A2(new_n520), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OAI211_X1 g429(.A(KEYINPUT106), .B(new_n510), .C1(new_n513), .C2(new_n514), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n730), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n695), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n859), .A2(new_n709), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n709), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n850), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n858), .B(new_n709), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n849), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n489), .B(KEYINPUT105), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n634), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT108), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n863), .A2(KEYINPUT108), .A3(new_n849), .ZN(new_n872));
  INV_X1    g447(.A(new_n868), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n862), .A4(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n869), .A2(new_n874), .A3(KEYINPUT40), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT40), .B1(new_n869), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(G395));
  OAI21_X1  g452(.A(KEYINPUT109), .B1(new_n611), .B2(G299), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n611), .A2(G299), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT109), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n827), .A2(new_n615), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT110), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT110), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n878), .A2(new_n884), .A3(new_n879), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n878), .A2(new_n888), .A3(new_n879), .A4(new_n881), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n836), .B(new_n620), .ZN(new_n891));
  MUX2_X1   g466(.A(new_n886), .B(new_n890), .S(new_n891), .Z(new_n892));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G303), .B(G288), .ZN(new_n895));
  XNOR2_X1  g470(.A(G290), .B(G305), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n895), .B(new_n896), .Z(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(new_n893), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n894), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(G868), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(G868), .B2(new_n823), .ZN(G295));
  OAI21_X1  g477(.A(new_n901), .B1(G868), .B2(new_n823), .ZN(G331));
  NAND2_X1  g478(.A1(new_n836), .A2(G168), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n834), .A2(G286), .A3(new_n835), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n904), .A2(G171), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G171), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n887), .B(new_n889), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(G301), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n904), .A2(G171), .A3(new_n905), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n882), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(KEYINPUT111), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n890), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n897), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n897), .B1(new_n913), .B2(new_n916), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n913), .A2(new_n916), .ZN(new_n923));
  INV_X1    g498(.A(new_n897), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n886), .A2(new_n911), .A3(new_n910), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n908), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n897), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n925), .A2(new_n926), .A3(new_n918), .A4(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n921), .A2(new_n922), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n918), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n932), .B2(new_n920), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g510(.A(KEYINPUT112), .B(KEYINPUT43), .C1(new_n932), .C2(new_n920), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n925), .A2(new_n926), .A3(new_n918), .A4(new_n917), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n931), .B1(new_n938), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g514(.A(G1384), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n856), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n481), .A2(new_n488), .A3(G40), .A4(new_n483), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n695), .B(G1996), .ZN(new_n946));
  INV_X1    g521(.A(G2067), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n730), .B(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n801), .B(new_n804), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(G290), .B(G1986), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1956), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n856), .B2(new_n940), .ZN(new_n955));
  INV_X1    g530(.A(new_n944), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n524), .A2(new_n940), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(KEYINPUT50), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n856), .A2(KEYINPUT45), .A3(new_n940), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n944), .B1(new_n957), .B2(new_n942), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT56), .B(G2072), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n615), .B(KEYINPUT57), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AND4_X1   g542(.A1(new_n940), .A2(new_n856), .A3(new_n947), .A4(new_n956), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n856), .A2(new_n954), .A3(new_n940), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n944), .B1(new_n957), .B2(KEYINPUT50), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1348), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n827), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n959), .A2(new_n963), .A3(new_n965), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT117), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n959), .A2(new_n963), .A3(KEYINPUT117), .A4(new_n965), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n973), .A2(KEYINPUT60), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n853), .B1(new_n515), .B2(new_n851), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n982), .B2(new_n855), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n947), .A3(new_n956), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n515), .B2(new_n523), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n956), .B1(new_n985), .B2(new_n954), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n954), .B2(new_n983), .ZN(new_n987));
  OAI211_X1 g562(.A(KEYINPUT60), .B(new_n984), .C1(new_n987), .C2(G1348), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT119), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n988), .A2(new_n989), .A3(new_n611), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n988), .B2(new_n611), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI211_X1 g567(.A(KEYINPUT50), .B(G1384), .C1(new_n982), .C2(new_n855), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n972), .B1(new_n993), .B2(new_n986), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n994), .A2(KEYINPUT60), .A3(new_n827), .A4(new_n984), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n973), .A2(KEYINPUT118), .A3(KEYINPUT60), .A4(new_n827), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n981), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n983), .A2(new_n956), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT58), .B(G1341), .Z(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n960), .A2(new_n961), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(new_n1004), .B2(G1996), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n570), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT59), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(KEYINPUT59), .A3(new_n570), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT61), .B1(new_n977), .B2(new_n978), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT61), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n967), .B2(new_n975), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1008), .B(new_n1009), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n980), .B1(new_n1000), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT122), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n1004), .B2(G2078), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(G2078), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n944), .B1(new_n985), .B2(KEYINPUT45), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1019), .B(new_n1020), .C1(new_n983), .C2(KEYINPUT45), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1961), .B1(new_n969), .B2(new_n970), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT121), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n770), .B1(new_n993), .B2(new_n986), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT121), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n1021), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1018), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1015), .B1(new_n1028), .B2(G301), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1022), .A2(new_n1023), .A3(KEYINPUT121), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1026), .B1(new_n1025), .B2(new_n1021), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1017), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n960), .A2(new_n1019), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n484), .A2(KEYINPUT123), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n481), .A2(new_n483), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n488), .A2(G40), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(KEYINPUT45), .B2(new_n983), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT124), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1035), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n943), .A2(KEYINPUT124), .A3(new_n1041), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT125), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT45), .B1(new_n856), .B2(new_n940), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1043), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1035), .ZN(new_n1050));
  AND4_X1   g625(.A1(KEYINPUT125), .A2(new_n1045), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1034), .B(G301), .C1(new_n1046), .C2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1029), .A2(new_n1033), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1034), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1054), .B1(new_n1056), .B2(G171), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT126), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1032), .B2(G171), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1028), .A2(KEYINPUT126), .A3(G301), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  INV_X1    g638(.A(G1966), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n956), .B1(new_n957), .B2(new_n942), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1047), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G2084), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n969), .A2(new_n970), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1063), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G286), .A2(G8), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1062), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(new_n1071), .ZN(new_n1075));
  AOI211_X1 g650(.A(KEYINPUT120), .B(new_n1070), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1069), .A2(new_n1062), .A3(new_n1071), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1063), .B1(new_n983), .B2(new_n956), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n587), .A2(G1976), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(KEYINPUT114), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1001), .A2(G8), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1001), .A2(G8), .A3(new_n1081), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1089));
  OR2_X1    g664(.A1(G305), .A2(G1981), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G305), .A2(G1981), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT49), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(KEYINPUT49), .A3(new_n1091), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1080), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AND4_X1   g671(.A1(new_n1084), .A2(new_n1087), .A3(new_n1089), .A4(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G303), .A2(G8), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT55), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT113), .B(G2090), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n993), .A2(new_n986), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1971), .B1(new_n960), .B2(new_n961), .ZN(new_n1104));
  OAI211_X1 g679(.A(G8), .B(new_n1100), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n944), .B1(new_n985), .B2(new_n954), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(new_n1101), .C1(new_n983), .C2(new_n954), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(G8), .B1(new_n1108), .B2(new_n1104), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1100), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1097), .A2(new_n1105), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1079), .A2(new_n1112), .ZN(new_n1113));
  AND4_X1   g688(.A1(new_n1014), .A2(new_n1055), .A3(new_n1061), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1004), .A2(new_n782), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1063), .B1(new_n1116), .B2(new_n1107), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1105), .B1(new_n1117), .B2(new_n1100), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1087), .A2(new_n1089), .A3(new_n1084), .A4(new_n1096), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1069), .A2(G168), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1115), .B1(new_n1121), .B2(KEYINPUT63), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT115), .B(new_n1123), .C1(new_n1112), .C2(new_n1120), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1116), .B1(new_n971), .B2(new_n1102), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(G8), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1097), .B(KEYINPUT116), .C1(new_n1126), .C2(new_n1100), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1100), .B1(new_n1125), .B2(G8), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n1119), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1105), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1131), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1122), .A2(new_n1124), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT62), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1078), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n1072), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1112), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1135), .A2(new_n1136), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1096), .A2(new_n1082), .A3(new_n587), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1090), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1097), .A2(new_n1131), .B1(new_n1144), .B2(new_n1080), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1134), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n952), .B1(new_n1114), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n948), .A2(new_n695), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n945), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT46), .ZN(new_n1150));
  INV_X1    g725(.A(G1996), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1150), .B1(new_n945), .B2(new_n1151), .ZN(new_n1152));
  NOR4_X1   g727(.A1(new_n943), .A2(KEYINPUT46), .A3(G1996), .A4(new_n944), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT47), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n950), .A2(new_n945), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1156), .B(KEYINPUT127), .Z(new_n1157));
  NOR2_X1   g732(.A1(G290), .A2(G1986), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n945), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT48), .Z(new_n1160));
  NOR2_X1   g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n804), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n802), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n946), .A2(new_n948), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(G2067), .B2(new_n730), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n1155), .B(new_n1161), .C1(new_n945), .C2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1147), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g742(.A1(new_n869), .A2(new_n874), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n921), .A2(new_n930), .ZN(new_n1170));
  INV_X1    g744(.A(G319), .ZN(new_n1171));
  NOR3_X1   g745(.A1(G401), .A2(new_n1171), .A3(G227), .ZN(new_n1172));
  NAND4_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n685), .A4(new_n1172), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


