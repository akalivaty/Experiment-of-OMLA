//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G8gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n208), .C1(G1gat), .C2(new_n202), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(G57gat), .A2(G64gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G57gat), .A2(G64gat), .ZN(new_n212));
  AND2_X1   g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(KEYINPUT9), .ZN(new_n214));
  NOR2_X1   g013(.A1(G71gat), .A2(G78gat), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n215), .A2(KEYINPUT91), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n213), .A2(new_n215), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n214), .B(new_n216), .C1(new_n215), .C2(new_n213), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n210), .B1(KEYINPUT21), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G127gat), .B(G155gat), .Z(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT20), .ZN(new_n226));
  NAND2_X1  g025(.A1(G231gat), .A2(G233gat), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n227), .B(KEYINPUT92), .Z(new_n228));
  XNOR2_X1  g027(.A(new_n226), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n224), .B(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n221), .A2(KEYINPUT21), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G211gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n230), .B(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G43gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G50gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(G50gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(KEYINPUT15), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G50gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT83), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT83), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G50gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n239), .B1(new_n248), .B2(new_n238), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT84), .B1(new_n249), .B2(KEYINPUT15), .ZN(new_n250));
  INV_X1    g049(.A(G29gat), .ZN(new_n251));
  INV_X1    g050(.A(G36gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT14), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT14), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(G29gat), .B2(G36gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(G29gat), .A2(G36gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n243), .B1(new_n250), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT84), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT15), .ZN(new_n261));
  AOI21_X1  g060(.A(G43gat), .B1(new_n245), .B2(new_n247), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n239), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n257), .B1(new_n263), .B2(new_n242), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT17), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT83), .B(G50gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n240), .B1(new_n266), .B2(G43gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n260), .B1(new_n267), .B2(new_n261), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n242), .B1(new_n268), .B2(new_n257), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n242), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n258), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT17), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G99gat), .B(G106gat), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G85gat), .A2(G92gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT7), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT7), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(G85gat), .A3(G92gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G99gat), .A2(G106gat), .ZN(new_n281));
  INV_X1    g080(.A(G85gat), .ZN(new_n282));
  INV_X1    g081(.A(G92gat), .ZN(new_n283));
  AOI22_X1  g082(.A1(KEYINPUT8), .A2(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT95), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n280), .B2(new_n284), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n275), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n280), .A2(new_n284), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT95), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n274), .A3(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n265), .A2(new_n273), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n246), .A2(G50gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n244), .A2(KEYINPUT83), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n238), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT15), .B1(new_n297), .B2(new_n240), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n258), .B1(new_n298), .B2(new_n260), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n264), .B1(new_n242), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(new_n292), .A3(new_n289), .ZN(new_n301));
  AND2_X1   g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT41), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n294), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(G190gat), .B(G218gat), .Z(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT96), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n304), .B(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n302), .A2(KEYINPUT41), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT94), .ZN(new_n309));
  INV_X1    g108(.A(G134gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(G162gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n307), .B(new_n312), .Z(new_n313));
  NAND2_X1  g112(.A1(G230gat), .A2(G233gat), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n219), .A2(new_n220), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n287), .A2(new_n275), .A3(new_n288), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n274), .B1(new_n291), .B2(new_n286), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT10), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n289), .A2(new_n221), .A3(new_n292), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n289), .A2(new_n221), .A3(KEYINPUT10), .A4(new_n292), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n321), .A2(KEYINPUT97), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT97), .B1(new_n321), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n314), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n314), .ZN(new_n326));
  INV_X1    g125(.A(new_n320), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n221), .B1(new_n289), .B2(new_n292), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT98), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G120gat), .B(G148gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(G176gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n333), .B(G204gat), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n329), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(KEYINPUT98), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n325), .A2(new_n331), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT99), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n322), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(new_n314), .ZN(new_n341));
  AOI211_X1 g140(.A(KEYINPUT99), .B(new_n326), .C1(new_n321), .C2(new_n322), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n341), .A2(new_n342), .A3(new_n336), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n338), .B1(new_n343), .B2(new_n334), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n237), .A2(new_n313), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n347));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348));
  INV_X1    g147(.A(G218gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n234), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(KEYINPUT22), .B2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G211gat), .B(G218gat), .Z(new_n352));
  AND2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n351), .A2(new_n352), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n347), .B1(new_n355), .B2(KEYINPUT29), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  OR2_X1    g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(G141gat), .A2(G148gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT2), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(G155gat), .B2(G162gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n357), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G155gat), .B(G162gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G155gat), .ZN(new_n367));
  INV_X1    g166(.A(G162gat), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT2), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n358), .A3(new_n359), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n364), .B1(new_n370), .B2(new_n357), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(new_n365), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n357), .A3(new_n364), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n347), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n355), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G228gat), .ZN(new_n382));
  INV_X1    g181(.A(G233gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n351), .B(new_n352), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n377), .B2(new_n378), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n381), .B(new_n385), .C1(KEYINPUT77), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G22gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n373), .B(new_n380), .C1(new_n390), .C2(new_n384), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT78), .ZN(new_n393));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT31), .B(G50gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n387), .B1(new_n372), .B2(new_n356), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n385), .B1(new_n387), .B2(KEYINPUT77), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  OAI21_X1  g199(.A(G22gat), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n393), .A2(new_n396), .B1(new_n392), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT78), .ZN(new_n403));
  AND4_X1   g202(.A1(new_n403), .A2(new_n401), .A3(new_n392), .A4(new_n396), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT76), .B(KEYINPUT0), .Z(new_n407));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G57gat), .B(G85gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT67), .B1(new_n310), .B2(G127gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G127gat), .B(G134gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(KEYINPUT67), .ZN(new_n416));
  INV_X1    g215(.A(G113gat), .ZN(new_n417));
  INV_X1    g216(.A(G120gat), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT1), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G113gat), .A2(G120gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n420), .A3(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n372), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n423), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n421), .B2(new_n416), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n376), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n413), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n374), .A2(KEYINPUT3), .A3(new_n375), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n377), .A2(new_n424), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n431), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n372), .A2(new_n424), .A3(KEYINPUT4), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n427), .B2(new_n376), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n434), .B(new_n435), .C1(new_n436), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(new_n439), .A3(KEYINPUT75), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n434), .B1(new_n436), .B2(new_n438), .ZN(new_n445));
  OR3_X1    g244(.A1(new_n445), .A2(KEYINPUT5), .A3(new_n431), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT80), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n432), .A2(new_n439), .A3(KEYINPUT75), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT75), .B1(new_n432), .B2(new_n439), .ZN(new_n449));
  OAI211_X1 g248(.A(KEYINPUT80), .B(new_n446), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n412), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G226gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(new_n383), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT27), .B(G183gat), .ZN(new_n455));
  INV_X1    g254(.A(G190gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(KEYINPUT28), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT66), .B(G183gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT27), .ZN(new_n459));
  OR2_X1    g258(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n460));
  AOI21_X1  g259(.A(G190gat), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n457), .B1(new_n461), .B2(KEYINPUT28), .ZN(new_n462));
  INV_X1    g261(.A(G169gat), .ZN(new_n463));
  INV_X1    g262(.A(G176gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT26), .ZN(new_n466));
  NOR2_X1   g265(.A1(G169gat), .A2(G176gat), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n468), .A2(new_n469), .B1(G183gat), .B2(G190gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n467), .A2(KEYINPUT23), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n467), .A2(KEYINPUT23), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n472), .A2(new_n473), .A3(new_n465), .ZN(new_n474));
  NAND3_X1  g273(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  OR2_X1    g275(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n456), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n479), .B2(KEYINPUT65), .ZN(new_n480));
  OAI22_X1  g279(.A1(new_n223), .A2(new_n456), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n481));
  AND2_X1   g280(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483));
  OAI22_X1  g282(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n475), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n474), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT25), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT25), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n223), .B2(new_n456), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(new_n475), .C1(G183gat), .C2(G190gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n471), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n454), .B1(new_n492), .B2(new_n378), .ZN(new_n493));
  INV_X1    g292(.A(new_n454), .ZN(new_n494));
  INV_X1    g293(.A(new_n491), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n462), .B2(new_n470), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n496), .B2(new_n486), .ZN(new_n497));
  OR3_X1    g296(.A1(new_n493), .A2(new_n355), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n355), .B1(new_n493), .B2(new_n497), .ZN(new_n499));
  XNOR2_X1  g298(.A(G8gat), .B(G36gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(G64gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(new_n283), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n502), .ZN(new_n506));
  INV_X1    g305(.A(new_n499), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n493), .A2(new_n355), .A3(new_n497), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT30), .A4(new_n502), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n505), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT79), .B1(new_n445), .B2(new_n431), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n445), .A2(KEYINPUT79), .A3(new_n431), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n425), .A2(new_n430), .A3(new_n428), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n513), .A2(KEYINPUT39), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT39), .ZN(new_n517));
  INV_X1    g316(.A(new_n514), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n512), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n519), .A3(new_n411), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT40), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n516), .A2(new_n519), .A3(KEYINPUT40), .A4(new_n411), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n452), .A2(new_n511), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT37), .B1(new_n507), .B2(new_n508), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT37), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n498), .A2(new_n499), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n506), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT38), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT38), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n525), .A2(new_n530), .A3(new_n527), .A4(new_n506), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n503), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(KEYINPUT6), .A3(new_n412), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT80), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n411), .B1(new_n536), .B2(new_n450), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n411), .B(new_n446), .C1(new_n448), .C2(new_n449), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n534), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n406), .B(new_n524), .C1(new_n532), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n492), .A2(new_n424), .ZN(new_n543));
  INV_X1    g342(.A(G227gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(new_n383), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n496), .A2(new_n427), .A3(new_n486), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT34), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n543), .A2(KEYINPUT34), .A3(new_n547), .A4(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT72), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n492), .A2(new_n424), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n427), .B1(new_n496), .B2(new_n486), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n545), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT70), .ZN(new_n559));
  XNOR2_X1  g358(.A(G71gat), .B(G99gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT68), .ZN(new_n561));
  INV_X1    g360(.A(G15gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n561), .A2(new_n562), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n564), .A2(new_n238), .A3(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n560), .B(KEYINPUT68), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(G15gat), .ZN(new_n568));
  AOI21_X1  g367(.A(G43gat), .B1(new_n568), .B2(new_n563), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n559), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n238), .B1(new_n564), .B2(new_n565), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n563), .A3(G43gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT70), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n573), .A3(KEYINPUT33), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n574), .A3(KEYINPUT32), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT71), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n558), .A2(new_n574), .A3(new_n577), .A4(KEYINPUT32), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n558), .A2(new_n580), .B1(new_n572), .B2(new_n571), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n558), .A2(KEYINPUT32), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT69), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT69), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n558), .A2(KEYINPUT32), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n546), .B1(new_n543), .B2(new_n547), .ZN(new_n587));
  OAI22_X1  g386(.A1(new_n587), .A2(KEYINPUT33), .B1(new_n566), .B2(new_n569), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n585), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n550), .A2(KEYINPUT72), .A3(new_n551), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n555), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n581), .A2(new_n582), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n593), .B1(new_n585), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n595), .A2(new_n554), .A3(new_n583), .A4(new_n579), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n592), .A2(new_n596), .A3(KEYINPUT36), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n542), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n411), .B1(new_n444), .B2(new_n446), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n534), .B1(new_n540), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n509), .A2(new_n510), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT73), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT73), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n509), .A2(new_n510), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n603), .A2(new_n505), .A3(new_n605), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n405), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n601), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT81), .ZN(new_n612));
  INV_X1    g411(.A(new_n540), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n452), .A2(new_n613), .B1(KEYINPUT6), .B2(new_n602), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n612), .B1(new_n614), .B2(new_n511), .ZN(new_n615));
  INV_X1    g414(.A(new_n511), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n541), .A2(KEYINPUT81), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g417(.A(KEYINPUT35), .B(new_n405), .C1(new_n592), .C2(new_n596), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n405), .B1(new_n592), .B2(new_n596), .ZN(new_n620));
  INV_X1    g419(.A(new_n608), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n618), .A2(new_n619), .B1(new_n622), .B2(KEYINPUT35), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n611), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT88), .ZN(new_n625));
  INV_X1    g424(.A(new_n210), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n265), .A2(new_n273), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n300), .B2(new_n210), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(KEYINPUT18), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT86), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT86), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n627), .A2(new_n630), .A3(new_n633), .A4(KEYINPUT18), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n627), .A2(new_n630), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n628), .B(KEYINPUT13), .Z(new_n639));
  NAND3_X1  g438(.A1(new_n269), .A2(new_n271), .A3(new_n210), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n210), .B1(new_n269), .B2(new_n271), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT87), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n300), .A2(KEYINPUT87), .A3(new_n210), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G169gat), .B(G197gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT12), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n638), .A2(new_n645), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n625), .B1(new_n635), .B2(new_n652), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n638), .A2(new_n645), .A3(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n632), .A2(new_n634), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(KEYINPUT88), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT87), .B1(new_n300), .B2(new_n210), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n642), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n640), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n639), .A2(new_n660), .B1(new_n636), .B2(new_n637), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n651), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT89), .B1(new_n657), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT89), .ZN(new_n665));
  AOI211_X1 g464(.A(new_n665), .B(new_n662), .C1(new_n653), .C2(new_n656), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT90), .B1(new_n624), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT35), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n597), .A2(new_n669), .A3(new_n406), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n617), .B2(new_n615), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n620), .B2(new_n621), .ZN(new_n672));
  OAI22_X1  g471(.A1(new_n671), .A2(new_n672), .B1(new_n610), .B2(new_n601), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT90), .ZN(new_n674));
  INV_X1    g473(.A(new_n667), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n346), .B1(new_n668), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n603), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT100), .B(G1gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1324gat));
  NAND2_X1  g480(.A1(new_n668), .A2(new_n676), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n511), .A3(new_n345), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT16), .B(G8gat), .Z(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT42), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n677), .A2(new_n687), .A3(new_n511), .A4(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n690));
  INV_X1    g489(.A(new_n683), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(new_n208), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n683), .A2(KEYINPUT101), .A3(G8gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n689), .A2(new_n692), .A3(new_n696), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1325gat));
  INV_X1    g497(.A(new_n600), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT36), .B1(new_n592), .B2(new_n596), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT103), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n562), .B1(new_n677), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n597), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(G15gat), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(new_n677), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT104), .ZN(G1326gat));
  NAND2_X1  g506(.A1(new_n677), .A2(new_n405), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(new_n344), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n237), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n313), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n682), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n251), .A3(new_n678), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n673), .B2(new_n313), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n609), .A2(KEYINPUT105), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n608), .A2(new_n722), .A3(new_n405), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n601), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n719), .B(new_n313), .C1(new_n725), .C2(new_n623), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT106), .ZN(new_n727));
  OAI22_X1  g526(.A1(new_n671), .A2(new_n672), .B1(new_n724), .B2(new_n601), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n728), .A2(new_n729), .A3(new_n719), .A4(new_n313), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n720), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n662), .B1(new_n653), .B2(new_n656), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n712), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G29gat), .B1(new_n736), .B2(new_n603), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n716), .A2(new_n717), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n718), .A2(new_n737), .A3(new_n738), .ZN(G1328gat));
  NAND3_X1  g538(.A1(new_n715), .A2(new_n252), .A3(new_n511), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n736), .A2(new_n616), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(KEYINPUT107), .ZN(new_n744));
  OAI21_X1  g543(.A(G36gat), .B1(new_n743), .B2(KEYINPUT107), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(G1329gat));
  OAI21_X1  g545(.A(G43gat), .B1(new_n736), .B2(new_n701), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n704), .A2(G43gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n715), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(KEYINPUT47), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n238), .B1(new_n735), .B2(new_n702), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n715), .B2(new_n748), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n752), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n682), .A2(new_n266), .A3(new_n405), .A4(new_n714), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(KEYINPUT109), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n731), .A2(new_n406), .A3(new_n734), .ZN(new_n757));
  OAI221_X1 g556(.A(new_n756), .B1(KEYINPUT109), .B2(new_n755), .C1(new_n266), .C2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n757), .B2(new_n266), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n727), .A2(new_n730), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n405), .B(new_n733), .C1(new_n761), .C2(new_n720), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(KEYINPUT108), .A3(new_n248), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n760), .A2(new_n763), .A3(new_n755), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n758), .B1(new_n764), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g564(.A1(new_n635), .A2(new_n625), .A3(new_n652), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT88), .B1(new_n654), .B2(new_n655), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n663), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n768), .A2(new_n237), .A3(new_n313), .A4(new_n711), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n728), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n678), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g572(.A1(new_n770), .A2(new_n616), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  AND2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(G1333gat));
  INV_X1    g577(.A(new_n702), .ZN(new_n779));
  OAI21_X1  g578(.A(G71gat), .B1(new_n770), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n704), .A2(G71gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g582(.A1(new_n771), .A2(new_n405), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g584(.A1(new_n768), .A2(new_n236), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n344), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n731), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n603), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n728), .A2(new_n313), .A3(new_n786), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT110), .Z(new_n794));
  NAND3_X1  g593(.A1(new_n678), .A2(new_n282), .A3(new_n344), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n790), .B1(new_n794), .B2(new_n795), .ZN(G1336gat));
  NOR2_X1   g595(.A1(new_n616), .A2(G92gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n344), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT111), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n793), .A2(new_n800), .A3(new_n344), .A4(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n283), .B1(new_n788), .B2(new_n511), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT52), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n798), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n803), .B2(new_n806), .ZN(G1337gat));
  OAI21_X1  g606(.A(G99gat), .B1(new_n789), .B2(new_n779), .ZN(new_n808));
  OR3_X1    g607(.A1(new_n704), .A2(G99gat), .A3(new_n711), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n794), .B2(new_n809), .ZN(G1338gat));
  INV_X1    g609(.A(G106gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n788), .B2(new_n405), .ZN(new_n812));
  AND4_X1   g611(.A1(new_n811), .A2(new_n793), .A3(new_n405), .A4(new_n344), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n812), .A2(new_n813), .A3(KEYINPUT53), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT53), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1339gat));
  NAND3_X1  g615(.A1(new_n321), .A2(new_n326), .A3(new_n322), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(KEYINPUT54), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n325), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n341), .B2(new_n342), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n819), .A2(new_n821), .A3(KEYINPUT55), .A4(new_n335), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n335), .A3(new_n821), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n768), .A2(new_n338), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n650), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n660), .A2(new_n639), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n628), .B1(new_n627), .B2(new_n640), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n344), .B(new_n830), .C1(new_n766), .C2(new_n767), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n657), .A2(KEYINPUT113), .A3(new_n344), .A4(new_n830), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n826), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n713), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n825), .A2(new_n338), .A3(new_n822), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n837), .A2(new_n657), .A3(new_n313), .A4(new_n830), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n237), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n346), .A2(new_n768), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n603), .A2(new_n511), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n620), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n768), .ZN(new_n848));
  INV_X1    g647(.A(new_n844), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n840), .B2(new_n842), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n620), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(new_n417), .A3(new_n667), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n848), .A2(new_n852), .ZN(G1340gat));
  AOI21_X1  g652(.A(G120gat), .B1(new_n847), .B2(new_n344), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n851), .A2(new_n418), .A3(new_n711), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(G1341gat));
  NAND4_X1  g655(.A1(new_n850), .A2(G127gat), .A3(new_n620), .A4(new_n236), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(KEYINPUT114), .ZN(new_n858));
  AOI21_X1  g657(.A(G127gat), .B1(new_n847), .B2(new_n236), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n857), .A2(KEYINPUT114), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G1342gat));
  NOR3_X1   g660(.A1(new_n846), .A2(G134gat), .A3(new_n713), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT56), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n851), .B2(new_n713), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1343gat));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n702), .A2(new_n406), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n850), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(G141gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n870), .A3(new_n675), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n236), .B1(new_n836), .B2(new_n838), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n873), .B(new_n405), .C1(new_n874), .C2(new_n841), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n699), .A2(new_n700), .A3(new_n849), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n825), .A2(new_n338), .A3(new_n822), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n768), .A2(new_n665), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n732), .A2(KEYINPUT89), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n831), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n657), .A2(KEYINPUT115), .A3(new_n344), .A4(new_n830), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n878), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n837), .B1(new_n664), .B2(new_n666), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(KEYINPUT116), .A3(new_n884), .A4(new_n885), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n889), .A3(new_n713), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n236), .B1(new_n890), .B2(new_n838), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n405), .B1(new_n891), .B2(new_n841), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n877), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n870), .B1(new_n893), .B2(new_n768), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT58), .B1(new_n872), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n877), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n890), .A2(new_n838), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n237), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n406), .B1(new_n898), .B2(new_n842), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n675), .B(new_n896), .C1(new_n899), .C2(new_n873), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT117), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n893), .A2(new_n902), .A3(new_n675), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n901), .A2(G141gat), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n871), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n866), .B(new_n895), .C1(new_n904), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n870), .B1(new_n900), .B2(KEYINPUT117), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n908), .B2(new_n903), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n896), .B1(new_n899), .B2(new_n873), .ZN(new_n910));
  OAI21_X1  g709(.A(G141gat), .B1(new_n910), .B2(new_n732), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n905), .B1(new_n911), .B2(new_n871), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT118), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n907), .A2(new_n913), .ZN(G1344gat));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  AOI211_X1 g714(.A(new_n915), .B(G148gat), .C1(new_n869), .C2(new_n344), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n873), .B1(new_n843), .B2(new_n405), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n667), .A2(new_n345), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT119), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n891), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n406), .A2(KEYINPUT57), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(new_n344), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(KEYINPUT59), .A3(new_n876), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n915), .B1(new_n910), .B2(new_n711), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n916), .B1(new_n926), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g726(.A(G155gat), .B1(new_n910), .B2(new_n237), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n869), .A2(new_n367), .A3(new_n236), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1346gat));
  OAI21_X1  g729(.A(G162gat), .B1(new_n910), .B2(new_n713), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n869), .A2(new_n368), .A3(new_n313), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT120), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n678), .A2(new_n616), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n843), .A2(new_n620), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G169gat), .B1(new_n936), .B2(new_n768), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n667), .A2(new_n463), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n936), .B2(new_n938), .ZN(G1348gat));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n344), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g740(.A1(new_n936), .A2(new_n236), .ZN(new_n942));
  MUX2_X1   g741(.A(new_n455), .B(new_n458), .S(new_n942), .Z(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g743(.A1(new_n936), .A2(new_n313), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G190gat), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(KEYINPUT121), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(G190gat), .A3(new_n949), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n948), .B(new_n950), .C1(G190gat), .C2(new_n945), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT122), .ZN(G1351gat));
  INV_X1    g751(.A(new_n935), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n702), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n405), .A3(new_n843), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n955), .A2(G197gat), .A3(new_n732), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT123), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n954), .B(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n922), .A3(new_n675), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G197gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n957), .A2(new_n961), .ZN(G1352gat));
  NAND2_X1  g761(.A1(new_n923), .A2(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G204gat), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n955), .A2(G204gat), .A3(new_n711), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1353gat));
  NAND2_X1  g766(.A1(new_n236), .A2(new_n234), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n955), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n959), .A2(new_n922), .A3(new_n236), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n234), .B1(KEYINPUT125), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n971), .A2(KEYINPUT125), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n975), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  NAND2_X1  g775(.A1(new_n313), .A2(G218gat), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n959), .A2(new_n922), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n349), .B1(new_n955), .B2(new_n713), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


