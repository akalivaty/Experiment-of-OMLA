//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  INV_X1    g0003(.A(G244), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G107), .A2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  AOI211_X1 g0010(.A(new_n205), .B(new_n210), .C1(G116), .C2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G1), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n220), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  OR2_X1    g0025(.A1(KEYINPUT64), .A2(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(KEYINPUT64), .A2(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AND2_X1   g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n214), .A2(new_n208), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n222), .B(new_n225), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT67), .B(G264), .ZN(new_n241));
  INV_X1    g0041(.A(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  AND2_X1   g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT69), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT69), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n230), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G222), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n265), .B(new_n267), .C1(new_n268), .C2(new_n266), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n260), .B(new_n269), .C1(G77), .C2(new_n265), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n217), .B(G274), .C1(G41), .C2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(new_n217), .A4(G274), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n217), .A2(new_n275), .B1(new_n230), .B2(new_n258), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G226), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n270), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G200), .ZN(new_n282));
  INV_X1    g0082(.A(G190), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n284), .A2(new_n255), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n228), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(G20), .B1(new_n232), .B2(G50), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(KEYINPUT71), .A2(G20), .A3(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G150), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n286), .B1(new_n291), .B2(new_n298), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n217), .A2(G13), .A3(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G50), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n285), .B1(G1), .B2(new_n218), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(G50), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT73), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n300), .A2(new_n301), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n282), .B1(new_n283), .B2(new_n281), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n310), .A2(KEYINPUT10), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT10), .B1(new_n310), .B2(new_n311), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n281), .A2(G179), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n281), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT74), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n285), .B2(new_n302), .ZN(new_n321));
  AND4_X1   g0121(.A1(new_n320), .A2(new_n302), .A3(new_n255), .A4(new_n284), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n217), .B2(G20), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n229), .A2(G77), .ZN(new_n325));
  XOR2_X1   g0125(.A(KEYINPUT15), .B(G87), .Z(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n325), .B1(new_n296), .B2(new_n287), .C1(new_n327), .C2(new_n290), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n324), .A2(G77), .B1(new_n286), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n303), .A2(new_n203), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n266), .A2(G232), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n265), .B(new_n332), .C1(new_n209), .C2(new_n266), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n260), .B(new_n333), .C1(G107), .C2(new_n265), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n279), .A2(G244), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n278), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n316), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n336), .A2(G179), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n331), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n319), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT7), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n265), .B2(G20), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n228), .A2(new_n347), .A3(KEYINPUT7), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n208), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(G58), .B(G68), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G20), .ZN(new_n351));
  INV_X1    g0151(.A(G159), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n296), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n342), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT7), .B1(new_n265), .B2(G20), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n228), .A2(new_n347), .A3(new_n343), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n356), .A3(G68), .ZN(new_n357));
  INV_X1    g0157(.A(new_n295), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n293), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G159), .B1(new_n350), .B2(G20), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n360), .A3(KEYINPUT16), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n354), .A2(new_n286), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n289), .A2(new_n302), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n287), .B(KEYINPUT70), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n305), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n256), .A2(new_n259), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G87), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n268), .A2(new_n266), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n213), .A2(G1698), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n369), .B(new_n370), .C1(new_n345), .C2(new_n346), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n367), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n275), .A2(new_n217), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n230), .A2(new_n258), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(G232), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n278), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(G200), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n371), .A2(new_n368), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n260), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(G232), .A2(new_n279), .B1(new_n272), .B2(new_n277), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(G190), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n362), .A2(new_n366), .A3(new_n377), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n362), .A2(new_n366), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n316), .B1(new_n372), .B2(new_n376), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT75), .ZN(new_n387));
  INV_X1    g0187(.A(G179), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n379), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n386), .B2(new_n389), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT76), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT76), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n372), .A2(new_n376), .A3(G179), .ZN(new_n394));
  AOI21_X1  g0194(.A(G169), .B1(new_n379), .B2(new_n380), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT75), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n385), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT76), .B1(new_n390), .B2(new_n391), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(new_n393), .A3(new_n397), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT18), .A3(new_n385), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n384), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n215), .A2(G1698), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n407), .B1(G226), .B2(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n260), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  AOI22_X1  g0212(.A1(G238), .A2(new_n279), .B1(new_n272), .B2(new_n277), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT14), .B1(new_n417), .B2(new_n316), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(G179), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT14), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n420), .B(G169), .C1(new_n415), .C2(new_n416), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n290), .A2(new_n203), .B1(new_n218), .B2(G68), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n296), .A2(new_n212), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n286), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT11), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n217), .A2(new_n208), .A3(G13), .A4(G20), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT12), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n426), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n321), .A2(new_n322), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(G68), .C1(G1), .C2(new_n218), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n427), .A2(new_n429), .A3(new_n430), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n422), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n417), .B2(G190), .ZN(new_n435));
  INV_X1    g0235(.A(G200), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(new_n417), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n406), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n336), .A2(new_n283), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n331), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n336), .A2(G200), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n341), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OR3_X1    g0245(.A1(new_n228), .A2(KEYINPUT23), .A3(G107), .ZN(new_n446));
  INV_X1    g0246(.A(G116), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n262), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G20), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n448), .A2(new_n218), .B1(new_n450), .B2(KEYINPUT23), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT22), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n226), .A2(new_n227), .B1(new_n263), .B2(new_n264), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(new_n453), .B2(G87), .ZN(new_n454));
  AND4_X1   g0254(.A1(new_n452), .A2(new_n228), .A3(new_n265), .A4(G87), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n446), .B(new_n451), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT24), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n228), .A2(new_n265), .ZN(new_n459));
  INV_X1    g0259(.A(G87), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT22), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n453), .A2(new_n452), .A3(G87), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(KEYINPUT24), .A3(new_n446), .A4(new_n451), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n458), .A2(new_n464), .A3(new_n286), .ZN(new_n465));
  INV_X1    g0265(.A(G13), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n450), .A2(G1), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n217), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n302), .A2(new_n471), .A3(new_n255), .A4(new_n284), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n469), .A2(new_n470), .B1(G107), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n274), .A2(G1), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G274), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(G264), .A3(new_n374), .ZN(new_n482));
  INV_X1    g0282(.A(G250), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n266), .ZN(new_n484));
  INV_X1    g0284(.A(G257), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G1698), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n484), .B(new_n486), .C1(new_n345), .C2(new_n346), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G294), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n481), .B(new_n482), .C1(new_n489), .C2(new_n367), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G169), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT80), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(new_n488), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n260), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(G179), .A3(new_n481), .A4(new_n482), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n491), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n492), .B1(new_n491), .B2(new_n495), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT81), .B1(new_n475), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n497), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n491), .A2(new_n492), .A3(new_n495), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n465), .A2(new_n474), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n494), .A2(new_n482), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(new_n283), .A4(new_n481), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT82), .B1(new_n490), .B2(G190), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n490), .A2(new_n436), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n474), .A3(new_n465), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(G97), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n472), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n449), .B1(new_n344), .B2(new_n348), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n296), .A2(new_n203), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n515), .A2(new_n449), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n449), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n228), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n517), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n516), .B1(new_n526), .B2(new_n286), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n303), .A2(new_n515), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n483), .B1(new_n263), .B2(new_n264), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT4), .ZN(new_n530));
  OAI21_X1  g0330(.A(G1698), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  OAI21_X1  g0332(.A(G244), .B1(new_n345), .B2(new_n346), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n530), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n260), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n479), .A2(new_n374), .ZN(new_n538));
  INV_X1    g0338(.A(G274), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n538), .A2(new_n485), .B1(new_n539), .B2(new_n479), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n540), .B1(new_n536), .B2(new_n260), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n527), .A2(new_n528), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n326), .A2(new_n302), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n472), .A2(new_n460), .ZN(new_n548));
  AND2_X1   g0348(.A1(KEYINPUT64), .A2(G20), .ZN(new_n549));
  NOR2_X1   g0349(.A1(KEYINPUT64), .A2(G20), .ZN(new_n550));
  OAI211_X1 g0350(.A(G33), .B(G97), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n228), .A2(new_n265), .A3(G68), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n549), .A2(new_n550), .B1(new_n552), .B2(new_n409), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n521), .A2(new_n460), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n547), .B(new_n548), .C1(new_n558), .C2(new_n286), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n483), .B1(new_n274), .B2(G1), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n217), .A2(new_n539), .A3(G45), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n374), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n209), .A2(new_n266), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n204), .A2(G1698), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n345), .C2(new_n346), .ZN(new_n566));
  INV_X1    g0366(.A(new_n448), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n563), .B1(new_n260), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G190), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n569), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G200), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n316), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n547), .B1(new_n558), .B2(new_n286), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n473), .A2(new_n326), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n575), .A2(new_n576), .B1(new_n388), .B2(new_n569), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n571), .A2(new_n573), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n516), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n528), .B(new_n579), .C1(new_n525), .C2(new_n285), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n542), .A2(new_n316), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n544), .A2(new_n388), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n546), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n266), .A2(G257), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G264), .A2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n586), .B(new_n587), .C1(new_n345), .C2(new_n346), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT77), .ZN(new_n589));
  INV_X1    g0389(.A(G303), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n263), .A2(new_n590), .A3(new_n264), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n588), .B2(new_n591), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n592), .A2(new_n593), .A3(new_n367), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n481), .B1(new_n538), .B2(new_n242), .ZN(new_n595));
  OAI21_X1  g0395(.A(G169), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n262), .A2(G97), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(new_n532), .C1(new_n549), .C2(new_n550), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n284), .A2(new_n255), .B1(G20), .B2(new_n447), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT20), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(KEYINPUT20), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(G116), .B(new_n471), .C1(new_n321), .C2(new_n322), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n303), .A2(new_n447), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n585), .B1(new_n596), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT78), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n588), .A2(new_n591), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT77), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n260), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n479), .A2(new_n374), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n616), .A2(G270), .B1(G274), .B2(new_n480), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n585), .B(new_n316), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n617), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n388), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n611), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n316), .B1(new_n615), .B2(new_n617), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n611), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(KEYINPUT78), .A3(new_n585), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(G200), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n625), .B(new_n607), .C1(new_n283), .C2(new_n619), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n610), .A2(new_n621), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n584), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n445), .A2(new_n514), .A3(new_n628), .ZN(G372));
  NAND3_X1  g0429(.A1(new_n610), .A2(new_n621), .A3(new_n624), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n465), .A2(new_n474), .B1(new_n491), .B2(new_n495), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT84), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n260), .A2(new_n568), .A3(KEYINPUT83), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT83), .B1(new_n260), .B2(new_n568), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n633), .A2(new_n634), .A3(new_n563), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n570), .B(new_n559), .C1(new_n635), .C2(new_n436), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n513), .A2(new_n546), .A3(new_n583), .A4(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT78), .B1(new_n623), .B2(new_n585), .ZN(new_n638));
  AOI211_X1 g0438(.A(new_n609), .B(KEYINPUT21), .C1(new_n622), .C2(new_n611), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT84), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n491), .A2(new_n495), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n504), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n640), .A2(new_n641), .A3(new_n621), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n632), .A2(new_n637), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT83), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n263), .A2(new_n264), .B1(new_n204), .B2(G1698), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n448), .B1(new_n647), .B2(new_n564), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n646), .B1(new_n648), .B2(new_n367), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n260), .A2(new_n568), .A3(KEYINPUT83), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n562), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n316), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n577), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n636), .A2(new_n653), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(new_n583), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT85), .ZN(new_n657));
  INV_X1    g0457(.A(new_n583), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n578), .A3(KEYINPUT26), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT85), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n660), .B(new_n654), .C1(new_n655), .C2(new_n583), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n657), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n645), .A2(new_n653), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n445), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT86), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT87), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n437), .A2(new_n340), .B1(new_n433), .B2(new_n422), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(new_n384), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n396), .A2(new_n397), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n385), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n400), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(KEYINPUT18), .A3(new_n385), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n666), .B1(new_n668), .B2(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n666), .B(new_n673), .C1(new_n667), .C2(new_n384), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n314), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n318), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n665), .A2(new_n678), .ZN(G369));
  INV_X1    g0479(.A(new_n630), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n228), .A2(G13), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT27), .B1(new_n681), .B2(G1), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT27), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n228), .A2(new_n683), .A3(new_n217), .A4(G13), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n687), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n514), .A2(new_n688), .B1(new_n631), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n514), .B1(new_n475), .B2(new_n689), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n502), .A2(new_n504), .A3(new_n687), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n689), .A2(new_n607), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n630), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n627), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n690), .B1(new_n694), .B2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n223), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n556), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n233), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n663), .A2(new_n689), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT88), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n663), .A2(KEYINPUT88), .A3(new_n689), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n546), .A2(new_n513), .A3(new_n583), .A4(new_n636), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n506), .B2(new_n680), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n658), .A2(new_n578), .A3(new_n654), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT26), .B1(new_n655), .B2(new_n583), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(new_n653), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT29), .B1(new_n719), .B2(new_n687), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n628), .A2(new_n506), .A3(new_n513), .A4(new_n689), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n635), .A2(G179), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n490), .A3(new_n542), .A4(new_n619), .ZN(new_n725));
  INV_X1    g0525(.A(new_n619), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n569), .A2(new_n494), .A3(new_n482), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(G179), .A4(new_n544), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n620), .A2(KEYINPUT30), .A3(new_n544), .A4(new_n727), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n687), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT31), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(new_n735), .A3(new_n687), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n722), .B1(new_n723), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n721), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n706), .B1(new_n739), .B2(G1), .ZN(G364));
  XOR2_X1   g0540(.A(new_n681), .B(KEYINPUT89), .Z(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G45), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G1), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n701), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n698), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n697), .A2(G330), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n255), .B1(G20), .B2(new_n316), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT93), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n228), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G179), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n750), .B1(new_n752), .B2(new_n436), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n751), .A2(KEYINPUT93), .A3(G179), .A4(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G179), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n229), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n756), .A2(new_n208), .B1(new_n515), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n436), .A2(G179), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n751), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n761), .B1(G107), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n229), .A2(G179), .A3(G190), .ZN(new_n766));
  OR3_X1    g0566(.A1(new_n766), .A2(KEYINPUT91), .A3(G200), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT91), .B1(new_n766), .B2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n766), .A2(new_n436), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n770), .A2(new_n214), .B1(new_n212), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n752), .A2(G200), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n773), .B1(G77), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(KEYINPUT92), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n762), .A2(G20), .A3(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n776), .B1(G87), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n347), .B1(new_n775), .B2(KEYINPUT92), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n751), .A2(new_n757), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n352), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  AND4_X1   g0583(.A1(new_n765), .A2(new_n779), .A3(new_n780), .A4(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G322), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT33), .B(G317), .Z(new_n786));
  OAI22_X1  g0586(.A1(new_n770), .A2(new_n785), .B1(new_n756), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G326), .B2(new_n771), .ZN(new_n788));
  INV_X1    g0588(.A(G329), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n347), .B1(new_n590), .B2(new_n777), .C1(new_n781), .C2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G283), .B2(new_n764), .ZN(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n788), .B(new_n791), .C1(new_n792), .C2(new_n760), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G311), .B2(new_n774), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n749), .B1(new_n784), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n795), .B1(new_n697), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n798), .A2(new_n749), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n223), .A2(new_n265), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT90), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G355), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n249), .A2(new_n274), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n700), .A2(new_n265), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G45), .B2(new_n233), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n804), .B1(G116), .B2(new_n223), .C1(new_n805), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n800), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n748), .B1(new_n809), .B2(new_n745), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT94), .Z(G396));
  AOI21_X1  g0611(.A(new_n689), .B1(new_n329), .B2(new_n330), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n339), .B1(new_n442), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n340), .A2(new_n689), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n663), .A2(new_n689), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n711), .B2(new_n815), .ZN(new_n817));
  INV_X1    g0617(.A(new_n738), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n744), .B1(new_n817), .B2(new_n818), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n813), .A2(new_n814), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n745), .B1(new_n823), .B2(new_n796), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n749), .A2(new_n796), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n769), .A2(G294), .B1(G97), .B2(new_n759), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT95), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n772), .A2(new_n590), .B1(new_n460), .B2(new_n763), .ZN(new_n829));
  INV_X1    g0629(.A(new_n781), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n265), .B(new_n829), .C1(G311), .C2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G283), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n832), .B1(new_n449), .B2(new_n777), .C1(new_n833), .C2(new_n756), .ZN(new_n834));
  INV_X1    g0634(.A(new_n774), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n447), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n755), .A2(G150), .B1(G159), .B2(new_n774), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n769), .A2(G143), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n772), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n830), .A2(G132), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n764), .A2(G68), .B1(G58), .B2(new_n759), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n347), .B1(new_n778), .B2(G50), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n834), .A2(new_n836), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT96), .ZN(new_n849));
  INV_X1    g0649(.A(new_n749), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n824), .B1(G77), .B2(new_n826), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n822), .A2(new_n851), .ZN(G384));
  NAND2_X1  g0652(.A1(new_n433), .A2(new_n687), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT99), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n422), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n854), .B2(new_n422), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n437), .A2(new_n434), .A3(new_n853), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n823), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n723), .A2(new_n737), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n685), .B(KEYINPUT100), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n385), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n865), .A2(new_n382), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n399), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n361), .A2(new_n286), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT16), .B1(new_n357), .B2(new_n360), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n366), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n685), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n669), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n873), .A2(new_n382), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n868), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n872), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n406), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n875), .B(KEYINPUT38), .C1(new_n406), .C2(new_n876), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n863), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT37), .B1(new_n404), .B2(new_n385), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n670), .A2(new_n382), .A3(new_n865), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n884), .A2(new_n866), .B1(KEYINPUT37), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n382), .B(KEYINPUT17), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n865), .B1(new_n673), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n878), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n883), .B1(new_n880), .B2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n882), .A2(new_n883), .B1(new_n863), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(G330), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n341), .A2(G330), .A3(new_n443), .A4(new_n862), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT102), .Z(new_n895));
  NAND3_X1  g0695(.A1(new_n891), .A2(new_n445), .A3(new_n862), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n434), .A2(new_n687), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n880), .A2(new_n899), .A3(new_n889), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n880), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT18), .B1(new_n404), .B2(new_n385), .ZN(new_n903));
  INV_X1    g0703(.A(new_n366), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n361), .A2(new_n286), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n905), .B2(new_n354), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n400), .B(new_n906), .C1(new_n402), .C2(new_n403), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n887), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n876), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n910), .B2(new_n875), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT39), .B1(new_n902), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n901), .B1(new_n912), .B2(KEYINPUT101), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT101), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n900), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n898), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n673), .A2(new_n864), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n816), .A2(new_n814), .ZN(new_n918));
  INV_X1    g0718(.A(new_n858), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n860), .A2(new_n919), .A3(new_n856), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n917), .B1(new_n921), .B2(new_n881), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n897), .B(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n677), .B1(new_n721), .B2(new_n445), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n217), .B2(new_n741), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n522), .A2(new_n523), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT35), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n231), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(G116), .C1(new_n929), .C2(new_n928), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  OAI21_X1  g0732(.A(G77), .B1(new_n214), .B2(new_n208), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n233), .A2(new_n933), .B1(G50), .B2(new_n208), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(G1), .A3(new_n466), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT98), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n927), .A2(new_n932), .A3(new_n936), .ZN(G367));
  XNOR2_X1  g0737(.A(new_n701), .B(KEYINPUT41), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n694), .A2(new_n698), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(KEYINPUT104), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n514), .A2(new_n688), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n693), .B2(new_n688), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(new_n746), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n739), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n580), .A2(new_n687), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n546), .A2(new_n583), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n583), .B2(new_n689), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n690), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT103), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT44), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n690), .A2(KEYINPUT103), .A3(new_n947), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n690), .A2(new_n947), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT45), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n951), .B1(new_n950), .B2(new_n952), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n939), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n940), .B(new_n944), .C1(new_n958), .C2(KEYINPUT104), .ZN(new_n959));
  INV_X1    g0759(.A(new_n739), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n938), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n743), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n514), .A2(new_n583), .A3(new_n546), .A4(new_n688), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT42), .Z(new_n965));
  OAI21_X1  g0765(.A(new_n583), .B1(new_n506), .B2(new_n946), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n689), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n689), .A2(new_n559), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n577), .A3(new_n652), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n655), .B2(new_n968), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n965), .A2(new_n967), .B1(KEYINPUT43), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n939), .A2(new_n947), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n971), .B(new_n972), .Z(new_n973));
  NOR2_X1   g0773(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n973), .B(new_n974), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n963), .A2(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n781), .A2(new_n839), .B1(new_n214), .B2(new_n777), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT105), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n347), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n212), .B2(new_n835), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n771), .A2(G143), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n203), .B2(new_n763), .C1(new_n977), .C2(new_n978), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(G68), .C2(new_n759), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n297), .B2(new_n770), .C1(new_n352), .C2(new_n756), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n347), .B1(new_n760), .B2(new_n449), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n764), .A2(G97), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n777), .A2(new_n447), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(KEYINPUT46), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n985), .B(new_n988), .C1(G317), .C2(new_n830), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n774), .A2(G283), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n755), .A2(G294), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n769), .A2(G303), .B1(G311), .B2(new_n771), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n987), .A2(KEYINPUT46), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n984), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n749), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n970), .A2(new_n799), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n245), .A2(new_n806), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n999), .B(new_n801), .C1(new_n223), .C2(new_n327), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n997), .A2(new_n744), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n976), .A2(new_n1001), .ZN(G387));
  OR3_X1    g0802(.A1(new_n287), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1003));
  AOI21_X1  g0803(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT50), .B1(new_n287), .B2(G50), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1003), .A2(new_n703), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n806), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n240), .B2(G45), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n803), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n703), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1006), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n700), .A2(new_n449), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n798), .B(new_n749), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n777), .A2(new_n203), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n830), .B2(G150), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT106), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n759), .A2(new_n326), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n755), .A2(new_n364), .B1(G68), .B2(new_n774), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT107), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(G159), .C2(new_n771), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n769), .A2(G50), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1021), .A2(new_n265), .A3(new_n986), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n755), .A2(G311), .B1(G322), .B2(new_n771), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n590), .B2(new_n835), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G317), .B2(new_n769), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT48), .Z(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n833), .B2(new_n760), .C1(new_n792), .C2(new_n777), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n764), .A2(G116), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n830), .A2(G326), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1030), .A2(new_n347), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n745), .B(new_n1013), .C1(new_n1035), .C2(new_n749), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n694), .A2(new_n798), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1036), .A2(new_n1037), .B1(new_n743), .B2(new_n943), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n739), .A2(new_n943), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1039), .A2(new_n701), .A3(new_n944), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(G393));
  AOI21_X1  g0841(.A(new_n944), .B1(new_n958), .B2(KEYINPUT104), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT104), .B2(new_n939), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n958), .A2(new_n944), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n701), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n958), .A2(new_n962), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n781), .A2(new_n785), .B1(new_n833), .B2(new_n777), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT111), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n347), .B1(new_n763), .B2(new_n449), .C1(new_n447), .C2(new_n760), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n769), .A2(G311), .B1(G317), .B2(new_n771), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1048), .B(new_n1049), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n792), .B2(new_n835), .C1(new_n590), .C2(new_n756), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT112), .Z(new_n1056));
  AOI22_X1  g0856(.A1(new_n769), .A2(G159), .B1(G150), .B2(new_n771), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT51), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G87), .B2(new_n764), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n287), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n755), .A2(G50), .B1(new_n1060), .B2(new_n774), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT109), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n830), .A2(G143), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n760), .A2(new_n203), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n265), .B1(new_n777), .B2(new_n208), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n1061), .C2(KEYINPUT109), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1059), .A2(new_n1062), .A3(new_n1063), .A4(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT110), .Z(new_n1068));
  OAI21_X1  g0868(.A(new_n749), .B1(new_n1056), .B2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n801), .B1(new_n515), .B2(new_n223), .C1(new_n1007), .C2(new_n252), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1069), .A2(new_n744), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n947), .A2(new_n799), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT108), .Z(new_n1073));
  AOI21_X1  g0873(.A(new_n1046), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1045), .A2(new_n1074), .ZN(G390));
  INV_X1    g0875(.A(new_n720), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n711), .B2(new_n712), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n678), .B(new_n893), .C1(new_n1077), .C2(new_n444), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT115), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n812), .B1(new_n440), .B2(new_n441), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n814), .B(new_n1079), .C1(new_n1080), .C2(new_n340), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n859), .A2(new_n860), .A3(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n738), .A2(new_n815), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1082), .B1(new_n738), .B2(new_n815), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n813), .B(new_n689), .C1(new_n715), .C2(new_n718), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n814), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n862), .A2(G330), .A3(new_n815), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1088), .A2(new_n920), .B1(new_n861), .B2(new_n738), .ZN(new_n1089));
  OAI21_X1  g0889(.A(KEYINPUT114), .B1(new_n1089), .B2(new_n918), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT114), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n816), .A2(new_n814), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n861), .A2(new_n738), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n859), .A2(new_n860), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n738), .B2(new_n815), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1091), .B(new_n1092), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1087), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1078), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n899), .B1(new_n879), .B2(new_n880), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n900), .B1(new_n1100), .B2(new_n914), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n915), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n921), .C2(new_n898), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT113), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n898), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n880), .A2(new_n889), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1106), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n920), .B1(new_n1085), .B2(new_n814), .ZN(new_n1110));
  OAI21_X1  g0910(.A(KEYINPUT113), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1103), .A2(new_n1112), .A3(new_n1093), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1093), .B1(new_n1103), .B2(new_n1112), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1099), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1078), .A2(new_n1098), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n898), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n913), .A2(new_n915), .A3(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1094), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1121), .A3(new_n1113), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1116), .A2(new_n701), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n743), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n913), .A2(new_n797), .A3(new_n915), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n830), .A2(G294), .B1(G87), .B2(new_n778), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n208), .B2(new_n763), .C1(new_n515), .C2(new_n835), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n265), .B(new_n1129), .C1(G107), .C2(new_n755), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1064), .B1(new_n769), .B2(G116), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT116), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(new_n833), .C2(new_n772), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n777), .A2(new_n297), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1135), .B1(new_n835), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n756), .A2(new_n839), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(G132), .C2(new_n769), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n764), .A2(G50), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n830), .A2(G125), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n265), .B1(new_n760), .B2(new_n352), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n771), .B2(G128), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1133), .A2(new_n1145), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n744), .B1(new_n364), .B2(new_n826), .C1(new_n1146), .C2(new_n850), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1126), .B1(new_n1127), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n1127), .B2(new_n1147), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1123), .A2(new_n1125), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(G378));
  INV_X1    g0951(.A(new_n1078), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1122), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n308), .A2(new_n872), .ZN(new_n1154));
  XOR2_X1   g0954(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n314), .B2(new_n318), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n318), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1158), .B(new_n1155), .C1(new_n312), .C2(new_n313), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1154), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1157), .A2(new_n1159), .A3(new_n1154), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT120), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n916), .B2(new_n922), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT120), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1168), .A2(new_n892), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n916), .A2(new_n1163), .A3(new_n922), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1165), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n892), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1170), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n1164), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1153), .A2(KEYINPUT57), .A3(new_n1171), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n701), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT121), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1153), .A2(new_n1171), .A3(new_n1174), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(new_n1181), .A3(new_n701), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1177), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1171), .A2(new_n1174), .A3(new_n743), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n212), .B1(new_n345), .B2(G41), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n774), .A2(new_n326), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n771), .A2(G116), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n830), .A2(G283), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n273), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n764), .A2(G58), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n208), .B2(new_n760), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1189), .A2(new_n1191), .A3(new_n265), .A4(new_n1014), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n515), .B2(new_n756), .C1(new_n449), .C2(new_n770), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT58), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1137), .A2(new_n777), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n771), .A2(G125), .B1(G150), .B2(new_n759), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT118), .Z(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(G132), .C2(new_n755), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n769), .A2(G128), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n839), .C2(new_n835), .ZN(new_n1200));
  XOR2_X1   g1000(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1201));
  OR2_X1    g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n764), .A2(G159), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G41), .B1(new_n830), .B2(G124), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n262), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1185), .B(new_n1194), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n745), .B1(new_n1207), .B2(new_n749), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(G50), .B2(new_n826), .C1(new_n1166), .C2(new_n797), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1184), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1183), .A2(new_n1210), .ZN(G375));
  OR3_X1    g1011(.A1(new_n1098), .A2(KEYINPUT122), .A3(new_n962), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n265), .B1(new_n771), .B2(G294), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(new_n1017), .C1(new_n449), .C2(new_n835), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n756), .A2(new_n447), .B1(new_n203), .B2(new_n763), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(G97), .C2(new_n778), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n833), .B2(new_n770), .C1(new_n590), .C2(new_n781), .ZN(new_n1217));
  INV_X1    g1017(.A(G128), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1190), .B1(new_n1218), .B2(new_n781), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n347), .B(new_n1219), .C1(G159), .C2(new_n778), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n212), .B2(new_n760), .C1(new_n297), .C2(new_n835), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT123), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n769), .A2(G137), .B1(G132), .B2(new_n771), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n756), .B2(new_n1137), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n749), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n825), .A2(new_n208), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n920), .A2(new_n796), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1226), .A2(new_n744), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT122), .B1(new_n1098), .B2(new_n962), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1212), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1078), .A2(new_n1098), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1099), .A2(new_n938), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(G381));
  INV_X1    g1034(.A(G390), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n976), .A2(new_n1235), .A3(new_n1001), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1236), .A2(G396), .A3(G393), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1183), .A2(new_n1150), .A3(new_n1210), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1238), .A2(G384), .A3(G381), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1237), .A2(KEYINPUT124), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT124), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1240), .A2(new_n1241), .ZN(G407));
  OAI221_X1 g1042(.A(G213), .B1(new_n1238), .B2(G343), .C1(new_n1240), .C2(new_n1241), .ZN(G409));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  INV_X1    g1044(.A(G213), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(G343), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1183), .A2(G378), .A3(new_n1210), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1153), .A2(new_n938), .A3(new_n1171), .A4(new_n1174), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1184), .A3(new_n1209), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT125), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1249), .A2(new_n1150), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1249), .B2(new_n1150), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1246), .B1(new_n1247), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1232), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1078), .A2(new_n1098), .A3(KEYINPUT60), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(new_n1099), .A3(new_n701), .A4(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G384), .A2(new_n1231), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1231), .B2(new_n1258), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(G2897), .A3(new_n1246), .ZN(new_n1264));
  INV_X1    g1064(.A(G2897), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1246), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1262), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1244), .B1(new_n1254), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT127), .B(new_n1244), .C1(new_n1254), .C2(new_n1268), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n975), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n961), .B2(new_n962), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1001), .ZN(new_n1276));
  OAI21_X1  g1076(.A(G390), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1236), .A2(new_n1277), .ZN(new_n1278));
  XOR2_X1   g1078(.A(G393), .B(G396), .Z(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1236), .A2(new_n1279), .A3(new_n1277), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1254), .A2(new_n1262), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT62), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1254), .A2(KEYINPUT62), .A3(new_n1262), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1283), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1247), .A2(new_n1253), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1266), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1268), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1284), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1254), .A2(KEYINPUT63), .A3(new_n1262), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1292), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1273), .A2(new_n1288), .B1(new_n1283), .B2(new_n1296), .ZN(G405));
  NAND2_X1  g1097(.A1(G375), .A2(new_n1150), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1247), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1262), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1247), .A3(new_n1263), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  XOR2_X1   g1102(.A(new_n1302), .B(new_n1283), .Z(G402));
endmodule


