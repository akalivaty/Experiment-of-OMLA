

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589;

  NOR2_X1 U319 ( .A1(n516), .A2(n472), .ZN(n575) );
  XOR2_X1 U320 ( .A(G1GAT), .B(G127GAT), .Z(n399) );
  INV_X1 U321 ( .A(KEYINPUT91), .ZN(n323) );
  XNOR2_X1 U322 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U323 ( .A(n326), .B(n325), .ZN(n329) );
  XNOR2_X1 U324 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n468) );
  XNOR2_X1 U325 ( .A(KEYINPUT102), .B(KEYINPUT36), .ZN(n313) );
  XNOR2_X1 U326 ( .A(n469), .B(n468), .ZN(n548) );
  XNOR2_X1 U327 ( .A(n569), .B(n313), .ZN(n587) );
  XNOR2_X1 U328 ( .A(n476), .B(KEYINPUT123), .ZN(n567) );
  XNOR2_X1 U329 ( .A(KEYINPUT93), .B(n392), .ZN(n516) );
  XNOR2_X1 U330 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U331 ( .A(n453), .B(G50GAT), .ZN(n454) );
  XNOR2_X1 U332 ( .A(n480), .B(n479), .ZN(G1349GAT) );
  XNOR2_X1 U333 ( .A(n455), .B(n454), .ZN(G1331GAT) );
  INV_X1 U334 ( .A(KEYINPUT103), .ZN(n448) );
  INV_X1 U335 ( .A(KEYINPUT79), .ZN(n312) );
  XOR2_X1 U336 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n289) );
  XNOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .ZN(n287) );
  XNOR2_X1 U338 ( .A(n287), .B(G218GAT), .ZN(n334) );
  XOR2_X1 U339 ( .A(G134GAT), .B(G162GAT), .Z(n318) );
  XNOR2_X1 U340 ( .A(n334), .B(n318), .ZN(n288) );
  XNOR2_X1 U341 ( .A(n289), .B(n288), .ZN(n293) );
  XOR2_X1 U342 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n291) );
  NAND2_X1 U343 ( .A1(G232GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U344 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n302) );
  INV_X1 U346 ( .A(G92GAT), .ZN(n294) );
  NAND2_X1 U347 ( .A1(KEYINPUT76), .A2(n294), .ZN(n297) );
  INV_X1 U348 ( .A(KEYINPUT76), .ZN(n295) );
  NAND2_X1 U349 ( .A1(n295), .A2(G92GAT), .ZN(n296) );
  NAND2_X1 U350 ( .A1(n297), .A2(n296), .ZN(n299) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(G85GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U353 ( .A(G106GAT), .B(n300), .Z(n419) );
  INV_X1 U354 ( .A(KEYINPUT10), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n419), .B(n301), .ZN(n303) );
  NAND2_X1 U356 ( .A1(n302), .A2(n303), .ZN(n307) );
  INV_X1 U357 ( .A(n302), .ZN(n305) );
  INV_X1 U358 ( .A(n303), .ZN(n304) );
  NAND2_X1 U359 ( .A1(n305), .A2(n304), .ZN(n306) );
  NAND2_X1 U360 ( .A1(n307), .A2(n306), .ZN(n311) );
  XOR2_X1 U361 ( .A(KEYINPUT8), .B(G50GAT), .Z(n309) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(G29GAT), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U364 ( .A(KEYINPUT7), .B(n310), .Z(n434) );
  XOR2_X1 U365 ( .A(n311), .B(n434), .Z(n561) );
  XNOR2_X1 U366 ( .A(n312), .B(n561), .ZN(n569) );
  XOR2_X1 U367 ( .A(G155GAT), .B(KEYINPUT2), .Z(n315) );
  XNOR2_X1 U368 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n357) );
  XOR2_X1 U370 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n317) );
  XNOR2_X1 U371 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n322) );
  XOR2_X1 U373 ( .A(G85GAT), .B(n399), .Z(n320) );
  XNOR2_X1 U374 ( .A(G29GAT), .B(n318), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U376 ( .A(n322), .B(n321), .Z(n326) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n327), .B(KEYINPUT0), .ZN(n373) );
  XNOR2_X1 U380 ( .A(n373), .B(KEYINPUT92), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U382 ( .A(n357), .B(n330), .Z(n332) );
  XOR2_X1 U383 ( .A(G120GAT), .B(G148GAT), .Z(n331) );
  XOR2_X1 U384 ( .A(G57GAT), .B(n331), .Z(n426) );
  XNOR2_X1 U385 ( .A(n332), .B(n426), .ZN(n392) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(G204GAT), .ZN(n333) );
  XOR2_X1 U387 ( .A(n333), .B(G64GAT), .Z(n425) );
  XOR2_X1 U388 ( .A(n334), .B(G92GAT), .Z(n336) );
  NAND2_X1 U389 ( .A1(G226GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n338) );
  XNOR2_X1 U391 ( .A(G8GAT), .B(G183GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n337), .B(G211GAT), .ZN(n400) );
  XOR2_X1 U393 ( .A(n338), .B(n400), .Z(n344) );
  XOR2_X1 U394 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n340) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n375) );
  XOR2_X1 U397 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n342) );
  XNOR2_X1 U398 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n360) );
  XNOR2_X1 U400 ( .A(n375), .B(n360), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n425), .B(n345), .ZN(n518) );
  XNOR2_X1 U403 ( .A(n518), .B(KEYINPUT27), .ZN(n388) );
  NAND2_X1 U404 ( .A1(n516), .A2(n388), .ZN(n547) );
  XOR2_X1 U405 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n347) );
  XNOR2_X1 U406 ( .A(KEYINPUT85), .B(KEYINPUT90), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U408 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n349) );
  XNOR2_X1 U409 ( .A(G148GAT), .B(KEYINPUT23), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U412 ( .A(G211GAT), .B(G162GAT), .Z(n353) );
  XNOR2_X1 U413 ( .A(G50GAT), .B(G22GAT), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U416 ( .A(n356), .B(G78GAT), .Z(n359) );
  XNOR2_X1 U417 ( .A(n357), .B(G204GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n365) );
  XOR2_X1 U419 ( .A(n360), .B(G106GAT), .Z(n362) );
  NAND2_X1 U420 ( .A1(G228GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U422 ( .A(G218GAT), .B(n363), .Z(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n473) );
  XOR2_X1 U424 ( .A(KEYINPUT28), .B(n473), .Z(n524) );
  NOR2_X1 U425 ( .A1(n547), .A2(n524), .ZN(n531) );
  XOR2_X1 U426 ( .A(G176GAT), .B(KEYINPUT67), .Z(n367) );
  XNOR2_X1 U427 ( .A(G120GAT), .B(KEYINPUT20), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n383) );
  XOR2_X1 U429 ( .A(G127GAT), .B(G71GAT), .Z(n369) );
  XNOR2_X1 U430 ( .A(G43GAT), .B(G134GAT), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n371) );
  XOR2_X1 U432 ( .A(G99GAT), .B(G190GAT), .Z(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n379) );
  XNOR2_X1 U434 ( .A(G183GAT), .B(KEYINPUT84), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n372), .B(KEYINPUT83), .ZN(n374) );
  XOR2_X1 U436 ( .A(n374), .B(n373), .Z(n377) );
  XNOR2_X1 U437 ( .A(G15GAT), .B(n375), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n381) );
  NAND2_X1 U440 ( .A1(G227GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n520) );
  INV_X1 U443 ( .A(n520), .ZN(n529) );
  NAND2_X1 U444 ( .A1(n531), .A2(n529), .ZN(n395) );
  NAND2_X1 U445 ( .A1(n520), .A2(n518), .ZN(n384) );
  NAND2_X1 U446 ( .A1(n384), .A2(n473), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n385), .B(KEYINPUT25), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n386), .B(KEYINPUT94), .ZN(n390) );
  NOR2_X1 U449 ( .A1(n520), .A2(n473), .ZN(n387) );
  XNOR2_X1 U450 ( .A(KEYINPUT26), .B(n387), .ZN(n574) );
  AND2_X1 U451 ( .A1(n388), .A2(n574), .ZN(n389) );
  NOR2_X1 U452 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n391), .B(KEYINPUT95), .ZN(n393) );
  NAND2_X1 U454 ( .A1(n393), .A2(n392), .ZN(n394) );
  NAND2_X1 U455 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n396), .B(KEYINPUT96), .ZN(n483) );
  XOR2_X1 U457 ( .A(KEYINPUT81), .B(G64GAT), .Z(n398) );
  XNOR2_X1 U458 ( .A(G155GAT), .B(G57GAT), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n413) );
  XOR2_X1 U460 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U461 ( .A1(G231GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U463 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n404) );
  XNOR2_X1 U464 ( .A(KEYINPUT80), .B(KEYINPUT15), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U466 ( .A(n406), .B(n405), .Z(n411) );
  XNOR2_X1 U467 ( .A(G15GAT), .B(G22GAT), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n407), .B(KEYINPUT70), .ZN(n433) );
  XOR2_X1 U469 ( .A(KEYINPUT13), .B(KEYINPUT73), .Z(n409) );
  XNOR2_X1 U470 ( .A(G71GAT), .B(G78GAT), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n420) );
  XNOR2_X1 U472 ( .A(n433), .B(n420), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U474 ( .A(n413), .B(n412), .Z(n481) );
  INV_X1 U475 ( .A(n481), .ZN(n583) );
  NAND2_X1 U476 ( .A1(n483), .A2(n583), .ZN(n414) );
  NOR2_X1 U477 ( .A1(n587), .A2(n414), .ZN(n415) );
  XNOR2_X1 U478 ( .A(KEYINPUT37), .B(n415), .ZN(n515) );
  XOR2_X1 U479 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n417) );
  XNOR2_X1 U480 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n419), .B(n418), .ZN(n430) );
  XOR2_X1 U483 ( .A(KEYINPUT75), .B(n420), .Z(n422) );
  NAND2_X1 U484 ( .A1(G230GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n424) );
  INV_X1 U486 ( .A(KEYINPUT77), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U488 ( .A(n426), .B(n425), .Z(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n580) );
  XOR2_X1 U491 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n432) );
  XNOR2_X1 U492 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n438) );
  XOR2_X1 U494 ( .A(G8GAT), .B(KEYINPUT69), .Z(n436) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n446) );
  NAND2_X1 U498 ( .A1(G229GAT), .A2(G233GAT), .ZN(n444) );
  XOR2_X1 U499 ( .A(G1GAT), .B(G197GAT), .Z(n440) );
  XNOR2_X1 U500 ( .A(G113GAT), .B(G141GAT), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U502 ( .A(G169GAT), .B(G36GAT), .Z(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n576) );
  XOR2_X1 U506 ( .A(n576), .B(KEYINPUT72), .Z(n563) );
  NAND2_X1 U507 ( .A1(n580), .A2(n563), .ZN(n486) );
  NOR2_X1 U508 ( .A1(n515), .A2(n486), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n447), .B(KEYINPUT38), .ZN(n449) );
  NAND2_X1 U510 ( .A1(n448), .A2(n449), .ZN(n452) );
  INV_X1 U511 ( .A(n449), .ZN(n450) );
  NAND2_X1 U512 ( .A1(KEYINPUT103), .A2(n450), .ZN(n451) );
  NAND2_X1 U513 ( .A1(n452), .A2(n451), .ZN(n501) );
  NAND2_X1 U514 ( .A1(n501), .A2(n524), .ZN(n455) );
  XOR2_X1 U515 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n453) );
  XNOR2_X1 U516 ( .A(KEYINPUT65), .B(KEYINPUT41), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n580), .B(n456), .ZN(n555) );
  XOR2_X1 U518 ( .A(n555), .B(KEYINPUT106), .Z(n535) );
  NOR2_X1 U519 ( .A1(n587), .A2(n583), .ZN(n458) );
  INV_X1 U520 ( .A(KEYINPUT45), .ZN(n457) );
  XNOR2_X1 U521 ( .A(n458), .B(n457), .ZN(n461) );
  INV_X1 U522 ( .A(n563), .ZN(n459) );
  NAND2_X1 U523 ( .A1(n580), .A2(n459), .ZN(n460) );
  NOR2_X1 U524 ( .A1(n461), .A2(n460), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n481), .B(KEYINPUT112), .ZN(n565) );
  NOR2_X1 U526 ( .A1(n555), .A2(n576), .ZN(n462) );
  XNOR2_X1 U527 ( .A(n462), .B(KEYINPUT46), .ZN(n463) );
  NOR2_X1 U528 ( .A1(n565), .A2(n463), .ZN(n464) );
  NAND2_X1 U529 ( .A1(n561), .A2(n464), .ZN(n465) );
  XNOR2_X1 U530 ( .A(n465), .B(KEYINPUT47), .ZN(n466) );
  NOR2_X1 U531 ( .A1(n467), .A2(n466), .ZN(n469) );
  XOR2_X1 U532 ( .A(KEYINPUT122), .B(n518), .Z(n470) );
  NOR2_X1 U533 ( .A1(n548), .A2(n470), .ZN(n471) );
  XOR2_X1 U534 ( .A(KEYINPUT54), .B(n471), .Z(n472) );
  NAND2_X1 U535 ( .A1(n575), .A2(n473), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n474), .B(KEYINPUT55), .ZN(n475) );
  NAND2_X1 U537 ( .A1(n475), .A2(n520), .ZN(n476) );
  NAND2_X1 U538 ( .A1(n535), .A2(n567), .ZN(n480) );
  XOR2_X1 U539 ( .A(G176GAT), .B(KEYINPUT56), .Z(n478) );
  XNOR2_X1 U540 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n477) );
  XOR2_X1 U541 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n488) );
  NAND2_X1 U542 ( .A1(n569), .A2(n481), .ZN(n482) );
  XOR2_X1 U543 ( .A(KEYINPUT16), .B(n482), .Z(n484) );
  NAND2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n485) );
  XOR2_X1 U545 ( .A(KEYINPUT97), .B(n485), .Z(n504) );
  NOR2_X1 U546 ( .A1(n486), .A2(n504), .ZN(n495) );
  NAND2_X1 U547 ( .A1(n495), .A2(n516), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U549 ( .A(G1GAT), .B(n489), .Z(G1324GAT) );
  NAND2_X1 U550 ( .A1(n495), .A2(n518), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n492) );
  NAND2_X1 U553 ( .A1(n495), .A2(n520), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n494) );
  XOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT99), .Z(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  XOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT101), .Z(n497) );
  NAND2_X1 U558 ( .A1(n495), .A2(n524), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(G1327GAT) );
  NAND2_X1 U560 ( .A1(n516), .A2(n501), .ZN(n499) );
  XOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U563 ( .A1(n501), .A2(n518), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U565 ( .A1(n501), .A2(n520), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n535), .A2(n576), .ZN(n514) );
  NOR2_X1 U569 ( .A1(n514), .A2(n504), .ZN(n505) );
  XOR2_X1 U570 ( .A(KEYINPUT107), .B(n505), .Z(n511) );
  NAND2_X1 U571 ( .A1(n511), .A2(n516), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(KEYINPUT42), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n518), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n520), .A2(n511), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n509), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U580 ( .A1(n511), .A2(n524), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n515), .A2(n514), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n516), .A2(n525), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n525), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n522) );
  NAND2_X1 U588 ( .A1(n525), .A2(n520), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n527) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n548), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(KEYINPUT113), .B(n532), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n563), .A2(n541), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT114), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U602 ( .A1(n541), .A2(n535), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n539) );
  NAND2_X1 U605 ( .A1(n541), .A2(n565), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  INV_X1 U608 ( .A(n541), .ZN(n542) );
  NOR2_X1 U609 ( .A1(n542), .A2(n569), .ZN(n546) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n544) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n549), .A2(n574), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n576), .A2(n560), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n555), .A2(n560), .ZN(n556) );
  XOR2_X1 U624 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U625 ( .A1(n583), .A2(n560), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NAND2_X1 U630 ( .A1(n567), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n567), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U634 ( .A(n567), .ZN(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n573) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT125), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT126), .B(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1351GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n586) );
  NOR2_X1 U641 ( .A1(n576), .A2(n586), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n586), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n586), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

