//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT11), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n193), .B2(G134), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n190), .A2(KEYINPUT64), .A3(G137), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n190), .A2(KEYINPUT64), .A3(G137), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT64), .B1(new_n190), .B2(G137), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n196), .B1(new_n204), .B2(new_n195), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT0), .A4(G128), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT0), .B(G128), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT82), .B1(new_n217), .B2(G104), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G107), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n217), .A2(KEYINPUT3), .A3(G104), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT3), .B1(new_n217), .B2(G104), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n218), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G101), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n216), .B1(new_n225), .B2(KEYINPUT4), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n220), .B2(G107), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n217), .A2(KEYINPUT3), .A3(G104), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G101), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n230), .A2(new_n231), .A3(new_n218), .A4(new_n221), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n225), .A2(KEYINPUT4), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT83), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n224), .B2(G101), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT83), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(new_n232), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n226), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT10), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT1), .B1(new_n210), .B2(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT85), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(KEYINPUT1), .C1(new_n210), .C2(G146), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(G128), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n209), .A2(new_n211), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n209), .A3(new_n211), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT65), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n213), .A2(new_n251), .A3(new_n248), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n245), .A2(new_n246), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT84), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n220), .B2(G107), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n220), .A2(G107), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n217), .A2(KEYINPUT84), .A3(G104), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G101), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n232), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n240), .B1(new_n253), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n250), .A2(new_n252), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT66), .A2(G128), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT66), .A2(G128), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n241), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n246), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n240), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n232), .A2(new_n259), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n207), .B1(new_n239), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n226), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n236), .A2(new_n237), .A3(new_n232), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n237), .B1(new_n236), .B2(new_n232), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n244), .A2(G128), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n243), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n246), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n262), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n268), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n280), .A2(new_n240), .B1(new_n268), .B2(new_n267), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n275), .A2(new_n281), .A3(new_n206), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n271), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G110), .B(G140), .ZN(new_n284));
  INV_X1    g098(.A(G953), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(G227), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n284), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n253), .A2(new_n260), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n250), .A2(new_n252), .B1(new_n246), .B2(new_n265), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n290), .A2(new_n260), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n207), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT12), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n260), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n260), .B2(new_n253), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT12), .A3(new_n207), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n287), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n282), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n288), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n189), .B1(new_n301), .B2(new_n187), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n299), .B1(new_n298), .B2(new_n282), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n271), .A2(new_n282), .A3(new_n299), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n293), .B(new_n206), .C1(new_n280), .C2(new_n295), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT12), .B1(new_n296), .B2(new_n207), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n239), .A2(new_n270), .A3(new_n207), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n287), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n271), .A2(new_n282), .A3(new_n299), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(KEYINPUT86), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n306), .A2(G469), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n302), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G221), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT9), .B(G234), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT81), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n316), .B1(new_n319), .B2(new_n188), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G475), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n324));
  AND2_X1   g138(.A1(KEYINPUT76), .A2(G140), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT76), .A2(G140), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n324), .B(G125), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  OR2_X1    g142(.A1(KEYINPUT76), .A2(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT76), .A2(G140), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n327), .B(KEYINPUT16), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n328), .A2(G140), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G146), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n208), .A3(new_n337), .ZN(new_n340));
  NOR2_X1   g154(.A1(G237), .A2(G953), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G214), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n210), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(G143), .A3(G214), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT17), .A3(G131), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(G131), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT17), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(new_n196), .A3(new_n344), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n339), .A2(new_n340), .A3(new_n346), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT18), .A2(G131), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n345), .B(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n335), .A2(new_n332), .A3(new_n208), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n327), .B(G146), .C1(new_n331), .C2(new_n333), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n353), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G113), .B(G122), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(new_n220), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n359), .B1(new_n351), .B2(new_n357), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n188), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n323), .B1(new_n363), .B2(KEYINPUT94), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(new_n188), .C1(new_n361), .C2(new_n362), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n327), .B(KEYINPUT19), .C1(new_n331), .C2(new_n333), .ZN(new_n367));
  OR2_X1    g181(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n335), .A2(new_n332), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n208), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n347), .A2(new_n349), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n339), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n357), .ZN(new_n375));
  INV_X1    g189(.A(new_n359), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n360), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n379));
  NOR2_X1   g193(.A1(G475), .A2(G902), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n359), .B1(new_n374), .B2(new_n357), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(new_n361), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT20), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n364), .A2(new_n366), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G116), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n217), .B1(new_n387), .B2(KEYINPUT14), .ZN(new_n388));
  INV_X1    g202(.A(G116), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G122), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n391), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n264), .A2(new_n263), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G143), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n210), .A2(G128), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n395), .A2(new_n190), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n190), .B1(new_n395), .B2(new_n396), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n392), .B(new_n393), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT13), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n396), .B(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n264), .A2(new_n263), .A3(new_n210), .ZN(new_n402));
  OAI21_X1  g216(.A(G134), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n391), .B(G107), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n395), .A2(new_n190), .A3(new_n396), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G217), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n318), .A2(new_n407), .A3(G953), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n399), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n399), .B2(new_n406), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n188), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT95), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  OAI211_X1 g229(.A(KEYINPUT95), .B(new_n188), .C1(new_n409), .C2(new_n410), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n411), .A2(new_n415), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n285), .A2(G952), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(G234), .B2(G237), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n188), .B(new_n285), .C1(G234), .C2(G237), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(G898), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n417), .A2(new_n418), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT96), .B1(new_n385), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n385), .A2(KEYINPUT96), .A3(new_n425), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n322), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G214), .B1(G237), .B2(G902), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G210), .B1(G237), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n290), .A2(new_n328), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT90), .B(G224), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n285), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n215), .A2(G125), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n435), .B2(new_n438), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n224), .A2(G101), .ZN(new_n442));
  INV_X1    g256(.A(G119), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G116), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n389), .A2(G119), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT67), .ZN(new_n447));
  XNOR2_X1  g261(.A(G116), .B(G119), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT67), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT2), .B(G113), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n446), .A2(new_n451), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n442), .A2(new_n235), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n273), .B2(new_n274), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n453), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n446), .A2(KEYINPUT67), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n448), .A2(new_n449), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT5), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G113), .ZN(new_n462));
  INV_X1    g276(.A(new_n444), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT5), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n458), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n268), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT87), .B(new_n454), .C1(new_n273), .C2(new_n274), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n457), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G122), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT89), .B(KEYINPUT6), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n467), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n234), .A2(new_n238), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT87), .B1(new_n476), .B2(new_n454), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n471), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n457), .A2(new_n470), .A3(new_n467), .A4(new_n468), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(KEYINPUT6), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT88), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n478), .A2(new_n479), .A3(new_n482), .A4(KEYINPUT6), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n441), .B(new_n474), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n470), .B(KEYINPUT8), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n448), .A2(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n465), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n487), .A2(new_n232), .A3(new_n453), .A4(new_n259), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n466), .A2(new_n268), .B1(KEYINPUT91), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n488), .A2(KEYINPUT91), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n437), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n439), .B2(new_n440), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n435), .A2(new_n438), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n492), .A3(new_n437), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n491), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n497), .B2(new_n479), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT92), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n434), .B1(new_n484), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n441), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n469), .B2(new_n471), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n482), .B1(new_n503), .B2(new_n479), .ZN(new_n504));
  INV_X1    g318(.A(new_n483), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n501), .B(new_n473), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n494), .A2(new_n496), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n507), .A2(new_n479), .A3(new_n491), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT92), .B1(new_n508), .B2(G902), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n498), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(new_n512), .A3(new_n433), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n432), .B1(new_n500), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n430), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(G472), .A2(G902), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n452), .A2(new_n453), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n193), .A2(G134), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n190), .A2(G137), .ZN(new_n520));
  OAI21_X1  g334(.A(G131), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n200), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n290), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n191), .A2(new_n194), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n198), .A2(new_n199), .ZN(new_n525));
  OAI21_X1  g339(.A(G131), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n215), .B1(new_n526), .B2(new_n200), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n523), .A2(new_n527), .A3(KEYINPUT30), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n251), .B1(new_n213), .B2(new_n248), .ZN(new_n530));
  AND4_X1   g344(.A1(new_n251), .A2(new_n248), .A3(new_n209), .A4(new_n211), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n266), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n521), .A3(new_n200), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n216), .B1(new_n201), .B2(new_n205), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n518), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n341), .A2(G210), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT27), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT26), .B(G101), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n518), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n533), .A2(new_n534), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n536), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n523), .A2(new_n527), .A3(new_n518), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT30), .B1(new_n523), .B2(new_n527), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n533), .A2(new_n534), .A3(new_n529), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n546), .B1(new_n549), .B2(new_n518), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT31), .A3(new_n540), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n540), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT28), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n542), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n518), .B1(new_n523), .B2(new_n527), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n554), .B1(new_n556), .B2(new_n542), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT68), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI211_X1 g373(.A(KEYINPUT68), .B(new_n554), .C1(new_n556), .C2(new_n542), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n553), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT32), .B(new_n517), .C1(new_n552), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT31), .B1(new_n550), .B2(new_n540), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n541), .B1(new_n547), .B2(new_n548), .ZN(new_n565));
  NOR4_X1   g379(.A1(new_n565), .A2(new_n544), .A3(new_n553), .A4(new_n546), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n561), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n563), .B1(new_n567), .B2(new_n516), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G472), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n536), .A2(new_n542), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT70), .B1(new_n571), .B2(new_n553), .ZN(new_n572));
  OAI211_X1 g386(.A(KEYINPUT70), .B(new_n553), .C1(new_n565), .C2(new_n546), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n541), .B1(new_n533), .B2(new_n534), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT28), .B1(new_n546), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT68), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n558), .B(KEYINPUT28), .C1(new_n546), .C2(new_n576), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n578), .A2(new_n540), .A3(new_n579), .A4(new_n555), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT69), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n582));
  INV_X1    g396(.A(new_n555), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n577), .B2(KEYINPUT68), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT69), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n540), .A4(new_n579), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n575), .A2(new_n581), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n583), .A2(KEYINPUT71), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT71), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n555), .A2(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n588), .A2(new_n557), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n553), .A2(new_n582), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n570), .B1(new_n587), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT72), .B1(new_n569), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT79), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT22), .B(G137), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n285), .A2(G221), .A3(G234), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n264), .A2(new_n263), .A3(new_n443), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n247), .A2(G119), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT73), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g417(.A1(KEYINPUT66), .A2(G128), .ZN(new_n604));
  NAND2_X1  g418(.A1(KEYINPUT66), .A2(G128), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(G119), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT73), .ZN(new_n607));
  INV_X1    g421(.A(new_n602), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G110), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT24), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT24), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G110), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n612), .A2(new_n614), .A3(KEYINPUT74), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT74), .B1(new_n612), .B2(new_n614), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n394), .A2(KEYINPUT23), .A3(G119), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT23), .B1(new_n247), .B2(G119), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n602), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n610), .A2(new_n617), .B1(G110), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n354), .B1(new_n338), .B2(G146), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n618), .A2(new_n620), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n611), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n339), .B2(new_n340), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n607), .B1(new_n606), .B2(new_n608), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n617), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT75), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g445(.A(KEYINPUT75), .B(new_n617), .C1(new_n627), .C2(new_n628), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI221_X4 g447(.A(new_n600), .B1(new_n622), .B2(new_n623), .C1(new_n626), .C2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n600), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n626), .A2(new_n633), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n623), .A2(new_n622), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n634), .A2(new_n638), .A3(G902), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT78), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n596), .B(new_n597), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n407), .B1(G234), .B2(new_n188), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT25), .B1(new_n639), .B2(new_n596), .ZN(new_n643));
  INV_X1    g457(.A(new_n632), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT75), .B1(new_n610), .B2(new_n617), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n334), .A2(new_n208), .A3(new_n337), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n208), .B1(new_n334), .B2(new_n337), .ZN(new_n648));
  OAI22_X1  g462(.A1(new_n647), .A2(new_n648), .B1(new_n611), .B2(new_n624), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n637), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n600), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n636), .A2(new_n637), .A3(new_n635), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n188), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT79), .B1(new_n653), .B2(KEYINPUT78), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n634), .A2(new_n638), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT80), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n642), .A2(G902), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT70), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n550), .B2(new_n540), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n586), .A2(new_n582), .A3(new_n663), .A4(new_n573), .ZN(new_n664));
  INV_X1    g478(.A(new_n581), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n593), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G472), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n584), .A2(new_n579), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n668), .A2(new_n553), .B1(new_n545), .B2(new_n551), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT32), .B1(new_n669), .B2(new_n517), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n517), .B1(new_n552), .B2(new_n561), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n563), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT72), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n667), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n595), .A2(new_n661), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n515), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n231), .ZN(G3));
  AND2_X1   g492(.A1(new_n413), .A2(new_n416), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT97), .B(G478), .Z(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR3_X1    g495(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT33), .ZN(new_n682));
  OAI21_X1  g496(.A(KEYINPUT33), .B1(new_n409), .B2(new_n410), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n188), .A2(G478), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n385), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n514), .A2(new_n424), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n552), .B2(new_n561), .ZN(new_n690));
  OAI22_X1  g504(.A1(new_n690), .A2(new_n570), .B1(new_n669), .B2(new_n517), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n660), .A2(new_n322), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n220), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G6));
  AOI21_X1  g510(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n364), .A2(new_n366), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n381), .A2(new_n384), .A3(KEYINPUT99), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n417), .A2(new_n418), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n514), .A2(new_n424), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n692), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT35), .B(G107), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G9));
  NOR2_X1   g522(.A1(new_n600), .A2(KEYINPUT36), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n650), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n658), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n655), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n567), .A2(new_n188), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n671), .B1(new_n713), .B2(G472), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT100), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n711), .ZN(new_n716));
  INV_X1    g530(.A(new_n642), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n654), .B2(new_n597), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n597), .B1(new_n653), .B2(KEYINPUT79), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n640), .B1(new_n656), .B2(new_n188), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n719), .B1(new_n720), .B2(KEYINPUT79), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n716), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n691), .A3(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n715), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n515), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT37), .B(G110), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT101), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n726), .B(new_n728), .ZN(G12));
  INV_X1    g543(.A(G900), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n421), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n420), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n699), .A2(new_n702), .A3(new_n700), .A4(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n322), .A2(new_n722), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n514), .A2(new_n735), .A3(new_n595), .A4(new_n675), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G128), .ZN(G30));
  AND3_X1   g551(.A1(new_n506), .A2(new_n512), .A3(new_n433), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n433), .B1(new_n506), .B2(new_n512), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT38), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT38), .B1(new_n500), .B2(new_n513), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n571), .A2(new_n540), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n556), .A2(new_n553), .A3(new_n542), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n188), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n570), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n670), .B2(new_n672), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n385), .A2(new_n703), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n431), .A2(new_n750), .A3(new_n722), .A4(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n320), .B1(new_n302), .B2(new_n314), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n733), .B(KEYINPUT39), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT40), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n743), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G143), .ZN(G45));
  NAND2_X1  g573(.A1(new_n364), .A2(new_n366), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n381), .A2(new_n384), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n686), .A2(new_n762), .A3(new_n733), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n322), .A2(new_n722), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n514), .A2(new_n764), .A3(new_n595), .A4(new_n675), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G146), .ZN(G48));
  NAND3_X1  g580(.A1(new_n514), .A2(new_n424), .A3(new_n688), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n288), .A2(new_n300), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n188), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(G469), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n301), .A2(new_n187), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n320), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n595), .A2(new_n675), .A3(new_n661), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT41), .B(G113), .Z(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G15));
  NAND3_X1  g591(.A1(new_n514), .A2(new_n424), .A3(new_n704), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n774), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n389), .ZN(G18));
  AOI21_X1  g594(.A(new_n722), .B1(new_n429), .B2(new_n427), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n595), .A3(new_n675), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n514), .A2(new_n773), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n443), .ZN(G21));
  OAI22_X1  g599(.A1(new_n591), .A2(new_n540), .B1(new_n564), .B2(new_n566), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n516), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(new_n570), .B2(new_n690), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n660), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n772), .A2(new_n320), .A3(new_n423), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n514), .A2(new_n751), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G122), .ZN(G24));
  NOR3_X1   g606(.A1(new_n722), .A2(new_n788), .A3(new_n763), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n514), .A2(new_n773), .A3(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(KEYINPUT102), .B(G125), .Z(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(G27));
  NOR3_X1   g610(.A1(new_n569), .A2(new_n594), .A3(KEYINPUT72), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n674), .B1(new_n667), .B2(new_n673), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n189), .B(KEYINPUT103), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n311), .A2(new_n312), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n801), .B2(new_n187), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n320), .B1(new_n803), .B2(new_n771), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n500), .A2(new_n431), .A3(new_n513), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n763), .A2(KEYINPUT42), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n799), .A2(new_n806), .A3(new_n661), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n667), .A2(new_n673), .ZN(new_n809));
  INV_X1    g623(.A(new_n763), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n661), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT42), .B1(new_n811), .B2(new_n805), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n196), .ZN(G33));
  NOR3_X1   g628(.A1(new_n676), .A2(new_n734), .A3(new_n805), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(new_n190), .ZN(G36));
  NAND3_X1  g630(.A1(new_n500), .A2(new_n431), .A3(new_n513), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n686), .A2(new_n385), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT43), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT43), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n686), .A2(new_n385), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT105), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n712), .A2(new_n823), .A3(new_n691), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT105), .B1(new_n722), .B2(new_n714), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n817), .B1(new_n826), .B2(KEYINPUT44), .ZN(new_n827));
  INV_X1    g641(.A(new_n822), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n823), .B1(new_n712), .B2(new_n691), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n722), .A2(new_n714), .A3(KEYINPUT105), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT44), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT104), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT45), .B1(new_n306), .B2(new_n313), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT45), .ZN(new_n836));
  OAI21_X1  g650(.A(G469), .B1(new_n801), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(KEYINPUT46), .B(new_n800), .C1(new_n835), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n834), .B1(new_n838), .B2(new_n771), .ZN(new_n839));
  INV_X1    g653(.A(new_n837), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n306), .A2(new_n313), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n840), .B1(new_n841), .B2(KEYINPUT45), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT46), .B1(new_n842), .B2(new_n800), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n838), .A2(new_n834), .A3(new_n771), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n320), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n827), .A2(new_n833), .A3(new_n846), .A4(new_n754), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G137), .ZN(G39));
  XNOR2_X1  g662(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n838), .A2(new_n834), .A3(new_n771), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n839), .A3(new_n843), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n852), .B2(new_n320), .ZN(new_n853));
  INV_X1    g667(.A(new_n839), .ZN(new_n854));
  INV_X1    g668(.A(new_n843), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n855), .A3(new_n845), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n321), .A3(new_n849), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n810), .A2(new_n660), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n799), .A2(new_n817), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n853), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(G140), .ZN(G42));
  INV_X1    g675(.A(KEYINPUT108), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n733), .B(KEYINPUT107), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n301), .A2(new_n187), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n321), .B(new_n863), .C1(new_n864), .C2(new_n802), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n749), .A2(new_n712), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n514), .A3(new_n751), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n736), .A2(new_n765), .A3(new_n867), .A4(new_n794), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n862), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n722), .A2(new_n788), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n810), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n805), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n703), .A2(new_n699), .A3(new_n700), .A4(new_n733), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n878), .A2(new_n712), .A3(new_n753), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n879), .A2(new_n595), .A3(new_n675), .ZN(new_n880));
  INV_X1    g694(.A(new_n817), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n676), .ZN(new_n883));
  INV_X1    g697(.A(new_n734), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n806), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n882), .A2(new_n812), .A3(new_n808), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n715), .A2(new_n724), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n514), .B(new_n430), .C1(new_n883), .C2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n774), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n689), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n705), .A2(new_n889), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n688), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n762), .B2(new_n703), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(new_n692), .A3(new_n514), .A4(new_n424), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n791), .C1(new_n783), .C2(new_n782), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n886), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT53), .B1(new_n874), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n892), .A2(new_n896), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n799), .A2(new_n881), .A3(new_n879), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n806), .A2(new_n793), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n813), .A2(new_n902), .A3(new_n815), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n799), .B(new_n514), .C1(new_n735), .C2(new_n764), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n904), .A2(KEYINPUT52), .A3(new_n794), .A4(new_n867), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n871), .A2(new_n905), .ZN(new_n906));
  AND4_X1   g720(.A1(KEYINPUT53), .A2(new_n899), .A3(new_n903), .A4(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT54), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n772), .A2(new_n320), .A3(new_n732), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n500), .A3(new_n431), .A4(new_n513), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n822), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n661), .A3(new_n809), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT48), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n828), .A2(new_n420), .A3(new_n789), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n783), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n419), .ZN(new_n916));
  INV_X1    g730(.A(new_n909), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n817), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n750), .A2(new_n660), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n913), .B(new_n916), .C1(new_n893), .C2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n301), .B(G469), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT109), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n432), .A4(new_n321), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n770), .A2(new_n432), .A3(new_n321), .A4(new_n771), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT109), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n741), .B2(new_n742), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT110), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(KEYINPUT110), .B(new_n927), .C1(new_n741), .C2(new_n742), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n914), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT50), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT50), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n935), .B(new_n914), .C1(new_n930), .C2(new_n931), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n686), .A2(new_n762), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n920), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n918), .A2(new_n828), .ZN(new_n941));
  INV_X1    g755(.A(new_n875), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT111), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR4_X1   g757(.A1(new_n910), .A2(new_n942), .A3(new_n822), .A4(KEYINPUT111), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n940), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n772), .A2(new_n321), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n853), .B2(new_n857), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n914), .A2(new_n817), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n946), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT51), .B1(new_n937), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n500), .A2(new_n513), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n740), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n500), .A2(KEYINPUT38), .A3(new_n513), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT110), .B1(new_n956), .B2(new_n927), .ZN(new_n957));
  INV_X1    g771(.A(new_n931), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n933), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n935), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n932), .A2(KEYINPUT50), .A3(new_n933), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT111), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n911), .B2(new_n875), .ZN(new_n964));
  OAI22_X1  g778(.A1(new_n964), .A2(new_n944), .B1(new_n920), .B2(new_n939), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n853), .A2(new_n857), .ZN(new_n966));
  INV_X1    g780(.A(new_n947), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n965), .B1(new_n968), .B2(new_n949), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT51), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n962), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n921), .B1(new_n952), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n874), .A2(new_n897), .A3(KEYINPUT53), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT53), .ZN(new_n974));
  INV_X1    g788(.A(new_n896), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n515), .B1(new_n725), .B2(new_n676), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n976), .A2(new_n775), .A3(new_n779), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n903), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n906), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT54), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n973), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n908), .A2(new_n972), .A3(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(G952), .A2(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n818), .A2(new_n432), .A3(new_n320), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n922), .B(KEYINPUT49), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n956), .A2(new_n919), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT112), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n985), .A2(KEYINPUT112), .A3(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(G75));
  NOR2_X1   g807(.A1(new_n285), .A2(G952), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n973), .A2(new_n980), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n996), .A2(G210), .A3(G902), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT56), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n473), .B1(new_n504), .B2(new_n505), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(new_n501), .ZN(new_n1001));
  XNOR2_X1  g815(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1001), .B(new_n1002), .Z(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT115), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n995), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1003), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(KEYINPUT114), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT114), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n999), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1005), .B1(new_n1008), .B2(new_n1010), .ZN(G51));
  INV_X1    g825(.A(new_n982), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n981), .B1(new_n973), .B2(new_n980), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n800), .B(KEYINPUT57), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n768), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n842), .B(KEYINPUT116), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n996), .A2(G902), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n994), .B1(new_n1016), .B2(new_n1018), .ZN(G54));
  AND4_X1   g833(.A1(KEYINPUT58), .A2(new_n996), .A3(G475), .A4(G902), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n995), .B1(new_n1020), .B2(new_n378), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n378), .B2(new_n1020), .ZN(G60));
  XNOR2_X1  g836(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n414), .A2(new_n188), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(new_n908), .B2(new_n982), .ZN(new_n1026));
  INV_X1    g840(.A(new_n684), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n995), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n684), .A2(new_n1025), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1029), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT118), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g846(.A(KEYINPUT118), .B(new_n1029), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1028), .B1(new_n1032), .B2(new_n1033), .ZN(G63));
  NAND2_X1  g848(.A1(G217), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT60), .Z(new_n1036));
  NAND2_X1  g850(.A1(new_n996), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(new_n657), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n996), .A2(new_n710), .A3(new_n1036), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1039), .A2(new_n995), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(KEYINPUT61), .B1(new_n1040), .B2(KEYINPUT119), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1041), .B(new_n1042), .ZN(G66));
  OAI21_X1  g857(.A(KEYINPUT120), .B1(new_n892), .B2(new_n896), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT120), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n977), .A2(new_n1045), .A3(new_n975), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1044), .A2(new_n1046), .A3(new_n285), .ZN(new_n1047));
  INV_X1    g861(.A(new_n436), .ZN(new_n1048));
  OAI21_X1  g862(.A(G953), .B1(new_n1048), .B2(new_n422), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n1050), .B(KEYINPUT121), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1000), .B1(G898), .B2(new_n285), .ZN(new_n1052));
  XOR2_X1   g866(.A(new_n1051), .B(new_n1052), .Z(G69));
  XNOR2_X1  g867(.A(new_n549), .B(new_n371), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1054), .B1(new_n730), .B2(new_n285), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n765), .A2(new_n736), .A3(new_n794), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1056), .A2(KEYINPUT123), .ZN(new_n1057));
  INV_X1    g871(.A(KEYINPUT123), .ZN(new_n1058));
  NAND4_X1  g872(.A1(new_n765), .A2(new_n736), .A3(new_n1058), .A4(new_n794), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  AND4_X1   g874(.A1(new_n661), .A2(new_n514), .A3(new_n809), .A4(new_n751), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1061), .A2(new_n846), .A3(new_n754), .ZN(new_n1062));
  NOR2_X1   g876(.A1(new_n813), .A2(new_n815), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n860), .A2(new_n847), .ZN(new_n1065));
  NOR2_X1   g879(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1055), .B1(new_n1066), .B2(new_n285), .ZN(new_n1067));
  AND2_X1   g881(.A1(new_n753), .A2(new_n754), .ZN(new_n1068));
  NAND4_X1  g882(.A1(new_n883), .A2(new_n1068), .A3(new_n881), .A4(new_n894), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n860), .A2(new_n847), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1058), .B1(new_n904), .B2(new_n794), .ZN(new_n1071));
  AND4_X1   g885(.A1(new_n1058), .A2(new_n765), .A3(new_n736), .A4(new_n794), .ZN(new_n1072));
  OAI21_X1  g886(.A(new_n758), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g887(.A(new_n1070), .B1(KEYINPUT62), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g888(.A(KEYINPUT62), .ZN(new_n1075));
  AND4_X1   g889(.A1(KEYINPUT124), .A2(new_n1060), .A3(new_n1075), .A4(new_n758), .ZN(new_n1076));
  INV_X1    g890(.A(new_n758), .ZN(new_n1077));
  AOI21_X1  g891(.A(new_n1077), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1078));
  AOI21_X1  g892(.A(KEYINPUT124), .B1(new_n1078), .B2(new_n1075), .ZN(new_n1079));
  OAI21_X1  g893(.A(new_n1074), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g894(.A1(new_n1080), .A2(new_n285), .ZN(new_n1081));
  XOR2_X1   g895(.A(new_n1054), .B(KEYINPUT122), .Z(new_n1082));
  AOI21_X1  g896(.A(new_n1067), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g897(.A(new_n285), .B1(G227), .B2(G900), .ZN(new_n1084));
  XOR2_X1   g898(.A(new_n1083), .B(new_n1084), .Z(G72));
  NAND2_X1  g899(.A1(G472), .A2(G902), .ZN(new_n1086));
  XOR2_X1   g900(.A(new_n1086), .B(KEYINPUT63), .Z(new_n1087));
  INV_X1    g901(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g902(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1089));
  AOI21_X1  g903(.A(new_n1088), .B1(new_n1066), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g904(.A1(new_n550), .A2(new_n553), .ZN(new_n1091));
  OAI21_X1  g905(.A(new_n995), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g906(.A1(new_n575), .A2(new_n543), .ZN(new_n1093));
  NAND2_X1  g907(.A1(new_n1093), .A2(new_n1087), .ZN(new_n1094));
  NAND2_X1  g908(.A1(new_n874), .A2(new_n897), .ZN(new_n1095));
  NAND2_X1  g909(.A1(new_n1095), .A2(new_n974), .ZN(new_n1096));
  NAND3_X1  g910(.A1(new_n897), .A2(KEYINPUT53), .A3(new_n906), .ZN(new_n1097));
  AOI21_X1  g911(.A(new_n1094), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g912(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g913(.A(KEYINPUT125), .ZN(new_n1100));
  OAI211_X1 g914(.A(new_n1074), .B(new_n1089), .C1(new_n1076), .C2(new_n1079), .ZN(new_n1101));
  NAND2_X1  g915(.A1(new_n1101), .A2(new_n1087), .ZN(new_n1102));
  INV_X1    g916(.A(new_n744), .ZN(new_n1103));
  AOI21_X1  g917(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g918(.A(KEYINPUT125), .B(new_n744), .C1(new_n1101), .C2(new_n1087), .ZN(new_n1105));
  OAI21_X1  g919(.A(new_n1099), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g920(.A(KEYINPUT126), .ZN(new_n1107));
  NAND2_X1  g921(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g922(.A(new_n1099), .B(KEYINPUT126), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1109));
  NAND2_X1  g923(.A1(new_n1108), .A2(new_n1109), .ZN(G57));
endmodule


