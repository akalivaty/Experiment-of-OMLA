//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(new_n465), .B2(G125), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT67), .A4(G125), .ZN(new_n467));
  INV_X1    g042(.A(G113), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(new_n461), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT68), .B1(new_n463), .B2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n473), .A3(new_n464), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n461), .A2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n477), .A2(KEYINPUT69), .B1(G101), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n480), .B1(new_n474), .B2(new_n476), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n470), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT70), .Z(G160));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n474), .B(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n485), .A2(new_n475), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  MUX2_X1   g064(.A(G100), .B(G112), .S(G2105), .Z(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2104), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n487), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NOR2_X1   g069(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(KEYINPUT68), .B2(new_n462), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(KEYINPUT73), .A3(new_n473), .A4(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n471), .A2(new_n473), .A3(new_n464), .A4(new_n497), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n475), .A2(G138), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT4), .B1(new_n474), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n465), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n475), .A2(G102), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT74), .B(G114), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(new_n475), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G2104), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n502), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OR3_X1    g091(.A1(new_n515), .A2(KEYINPUT75), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT75), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(new_n514), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n524), .A2(G88), .B1(new_n525), .B2(G50), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n521), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n523), .B2(new_n531), .ZN(new_n532));
  XOR2_X1   g107(.A(new_n532), .B(KEYINPUT76), .Z(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n525), .A2(G51), .B1(new_n514), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G168));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n522), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n523), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n515), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n542), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n549), .B1(new_n548), .B2(new_n547), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n524), .A2(G81), .B1(new_n525), .B2(G43), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT78), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  XOR2_X1   g131(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n557));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n525), .A2(G53), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n524), .A2(G91), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n542), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(G299));
  XNOR2_X1  g141(.A(G171), .B(KEYINPUT80), .ZN(G301));
  NAND2_X1  g142(.A1(new_n533), .A2(new_n535), .ZN(G286));
  NAND2_X1  g143(.A1(new_n524), .A2(G87), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n525), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT81), .ZN(G288));
  AOI22_X1  g148(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n542), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT82), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n575), .B(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n524), .A2(G86), .B1(new_n525), .B2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G305));
  INV_X1    g154(.A(G85), .ZN(new_n580));
  INV_X1    g155(.A(G47), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n523), .A2(new_n580), .B1(new_n538), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n542), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n514), .A2(new_n522), .A3(G92), .ZN(new_n588));
  XOR2_X1   g163(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n589));
  XOR2_X1   g164(.A(new_n588), .B(new_n589), .Z(new_n590));
  XNOR2_X1  g165(.A(KEYINPUT84), .B(G66), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n514), .A2(new_n591), .B1(G79), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n592), .A2(new_n542), .B1(new_n593), .B2(new_n538), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n587), .B1(G868), .B2(new_n595), .ZN(G284));
  OAI21_X1  g171(.A(new_n587), .B1(G868), .B2(new_n595), .ZN(G321));
  MUX2_X1   g172(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g173(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n595), .B1(new_n600), .B2(G860), .ZN(G148));
  INV_X1    g176(.A(new_n595), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G559), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n552), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(G282));
  INV_X1    g184(.A(new_n607), .ZN(G323));
  NAND2_X1  g185(.A1(new_n465), .A2(new_n478), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT12), .Z(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT13), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n488), .A2(G135), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n486), .A2(G123), .ZN(new_n616));
  AND2_X1   g191(.A1(G111), .A2(G2105), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(G99), .B2(new_n475), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(new_n461), .C2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2096), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2096), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n614), .A2(new_n620), .A3(new_n621), .ZN(G156));
  XOR2_X1   g197(.A(KEYINPUT15), .B(G2435), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2427), .ZN(new_n625));
  INV_X1    g200(.A(G2430), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XOR2_X1   g207(.A(new_n631), .B(new_n632), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n629), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT86), .ZN(new_n637));
  OAI21_X1  g212(.A(G14), .B1(new_n634), .B2(new_n635), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  INV_X1    g221(.A(new_n642), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n643), .B1(new_n649), .B2(new_n640), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n641), .B2(new_n648), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n641), .A2(new_n644), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n647), .B1(new_n652), .B2(KEYINPUT17), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n646), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT20), .Z(new_n665));
  AOI211_X1 g240(.A(new_n663), .B(new_n665), .C1(new_n658), .C2(new_n662), .ZN(new_n666));
  XOR2_X1   g241(.A(G1981), .B(G1986), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n668), .B(new_n672), .ZN(G229));
  MUX2_X1   g248(.A(G6), .B(G305), .S(G16), .Z(new_n674));
  XOR2_X1   g249(.A(KEYINPUT32), .B(G1981), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(G166), .A2(G16), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G16), .B2(G22), .ZN(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G23), .ZN(new_n683));
  INV_X1    g258(.A(new_n572), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT33), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n676), .A2(new_n680), .A3(new_n681), .A4(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n690));
  NOR2_X1   g265(.A1(G25), .A2(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n488), .A2(G131), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n486), .A2(G119), .ZN(new_n693));
  MUX2_X1   g268(.A(G95), .B(G107), .S(G2105), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G2104), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n691), .B1(new_n697), .B2(G29), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G16), .A2(G24), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n585), .B2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n689), .A2(new_n690), .A3(new_n700), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT36), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n488), .A2(G139), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n708));
  AOI21_X1  g283(.A(KEYINPUT25), .B1(new_n478), .B2(G103), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n478), .A2(KEYINPUT25), .A3(G103), .ZN(new_n710));
  OAI221_X1 g285(.A(new_n707), .B1(new_n475), .B2(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G33), .B(new_n711), .S(G29), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G2072), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G32), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n488), .A2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n486), .A2(G129), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT26), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n720), .A2(new_n721), .B1(G105), .B2(new_n478), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n716), .A2(new_n717), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n715), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n713), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(G168), .A2(G16), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G21), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(KEYINPUT92), .B2(new_n727), .ZN(new_n731));
  INV_X1    g306(.A(G1966), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n724), .A2(new_n725), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT31), .B(G11), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT30), .B(G28), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n714), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n619), .B2(new_n714), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT93), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n682), .A2(G20), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT23), .Z(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G299), .B2(G16), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(G1956), .Z(new_n744));
  NAND2_X1  g319(.A1(G164), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G27), .B2(G29), .ZN(new_n746));
  INV_X1    g321(.A(G2078), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n682), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n682), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1961), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n744), .A2(new_n748), .A3(new_n749), .A4(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n726), .A2(new_n735), .A3(new_n740), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G29), .A2(G35), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G162), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2090), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(KEYINPUT24), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(KEYINPUT24), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n714), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n714), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT91), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2084), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n754), .A2(new_n758), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n714), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n488), .A2(G140), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT88), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(new_n475), .B2(G116), .ZN(new_n771));
  OR3_X1    g346(.A1(KEYINPUT89), .A2(G104), .A3(G2105), .ZN(new_n772));
  OAI21_X1  g347(.A(KEYINPUT89), .B1(G104), .B2(G2105), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n486), .B2(G128), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G16), .A2(G19), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n552), .B2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n595), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G4), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1348), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n779), .A2(new_n782), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT90), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n706), .A2(new_n766), .A3(new_n789), .ZN(G150));
  INV_X1    g365(.A(G150), .ZN(G311));
  INV_X1    g366(.A(G93), .ZN(new_n792));
  INV_X1    g367(.A(G55), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n523), .A2(new_n792), .B1(new_n538), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(new_n542), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n552), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n595), .A2(G559), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT39), .ZN(new_n804));
  INV_X1    g379(.A(G860), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(KEYINPUT39), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n797), .A2(new_n805), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT37), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT95), .ZN(G145));
  XNOR2_X1  g386(.A(new_n776), .B(new_n512), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n711), .B(new_n723), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n812), .B(new_n813), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n696), .B(new_n612), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n486), .A2(G130), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n475), .A2(KEYINPUT96), .A3(G118), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT96), .B1(new_n475), .B2(G118), .ZN(new_n818));
  OR2_X1    g393(.A1(G106), .A2(G2105), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n818), .A2(G2104), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n816), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G142), .B2(new_n488), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n815), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n814), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n825), .A2(new_n826), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n814), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n828), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(G160), .B(new_n619), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G162), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n812), .B(new_n813), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n835), .B1(new_n837), .B2(new_n823), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n827), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n836), .A2(new_n841), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n839), .A2(new_n840), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT99), .B1(new_n827), .B2(new_n838), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n835), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n831), .B1(KEYINPUT98), .B2(new_n827), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(new_n828), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n843), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n845), .A2(new_n852), .ZN(G395));
  NOR2_X1   g428(.A1(new_n798), .A2(G868), .ZN(new_n854));
  XNOR2_X1  g429(.A(G305), .B(G303), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n585), .B(new_n572), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT103), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT42), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(KEYINPUT42), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(KEYINPUT104), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(KEYINPUT104), .B2(new_n859), .ZN(new_n862));
  INV_X1    g437(.A(G299), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n602), .ZN(new_n864));
  NAND2_X1  g439(.A1(G299), .A2(new_n595), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n865), .B(KEYINPUT101), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n864), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n871), .A2(KEYINPUT102), .A3(KEYINPUT41), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT102), .B1(new_n871), .B2(KEYINPUT41), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n799), .B(new_n603), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n871), .B2(new_n875), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n862), .B(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n854), .B1(new_n878), .B2(G868), .ZN(G295));
  AOI21_X1  g454(.A(new_n854), .B1(new_n878), .B2(G868), .ZN(G331));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n881));
  NAND3_X1  g456(.A1(G286), .A2(KEYINPUT105), .A3(G171), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(G168), .B2(G301), .ZN(new_n884));
  INV_X1    g459(.A(G171), .ZN(new_n885));
  NOR2_X1   g460(.A1(G168), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n882), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n887), .A2(new_n799), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n799), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n888), .A2(new_n892), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n874), .A2(new_n893), .B1(new_n870), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n895), .B2(new_n858), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n870), .A2(new_n897), .A3(new_n867), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT107), .B1(new_n864), .B2(new_n865), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n867), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n870), .A2(new_n897), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n893), .A2(new_n871), .B1(new_n902), .B2(new_n894), .ZN(new_n903));
  INV_X1    g478(.A(new_n858), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n895), .A2(new_n858), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n909), .A3(new_n896), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n881), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n909), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(KEYINPUT43), .A3(new_n896), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n911), .A2(new_n914), .ZN(G397));
  INV_X1    g490(.A(G1384), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n499), .A2(new_n500), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n499), .A2(new_n500), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n511), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n504), .A2(new_n506), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n470), .A2(new_n479), .A3(G40), .A4(new_n481), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n776), .A2(G2067), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n770), .A2(new_n778), .A3(new_n775), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT108), .ZN(new_n930));
  INV_X1    g505(.A(G1996), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n723), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n929), .A2(KEYINPUT108), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n697), .A2(new_n699), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n926), .B1(new_n937), .B2(new_n928), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n927), .A2(new_n928), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n925), .B1(new_n939), .B2(new_n723), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n925), .B(new_n931), .C1(KEYINPUT127), .C2(KEYINPUT46), .ZN(new_n941));
  NAND2_X1  g516(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n941), .B(new_n942), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT47), .Z(new_n945));
  NOR2_X1   g520(.A1(new_n697), .A2(new_n699), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n925), .B1(new_n936), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(G290), .A2(G1986), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n925), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT48), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n935), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n938), .A2(new_n945), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n585), .A2(new_n703), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n925), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n935), .A2(new_n954), .A3(new_n947), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT109), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n935), .A2(new_n957), .A3(new_n954), .A4(new_n947), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n924), .B1(new_n921), .B2(new_n922), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n916), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT56), .B(G2072), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n921), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n512), .A2(KEYINPUT110), .A3(new_n916), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(KEYINPUT50), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n921), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n924), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n963), .B1(new_n970), .B2(G1956), .ZN(new_n971));
  XNOR2_X1  g546(.A(G299), .B(KEYINPUT57), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n924), .B1(new_n921), .B2(KEYINPUT50), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n498), .A2(new_n501), .B1(G2104), .B2(new_n510), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n964), .B(G1384), .C1(new_n977), .C2(new_n507), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT110), .B1(new_n512), .B2(new_n916), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n980), .B2(new_n968), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n965), .A2(new_n976), .A3(new_n968), .A4(new_n966), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n975), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT120), .ZN(new_n985));
  INV_X1    g560(.A(new_n975), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n965), .A2(new_n968), .A3(new_n966), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n988), .B2(new_n982), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT120), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n785), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT119), .ZN(new_n993));
  INV_X1    g568(.A(new_n924), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n965), .A2(new_n966), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n965), .A2(new_n994), .A3(KEYINPUT118), .A4(new_n966), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n999), .B2(new_n778), .ZN(new_n1000));
  AOI211_X1 g575(.A(KEYINPUT119), .B(G2067), .C1(new_n997), .C2(new_n998), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n602), .B1(new_n992), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n972), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n963), .C1(new_n970), .C2(G1956), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n974), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n973), .A2(KEYINPUT61), .A3(new_n1005), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT61), .B1(new_n973), .B2(new_n1005), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n992), .A2(new_n1002), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n1012));
  XOR2_X1   g587(.A(KEYINPUT58), .B(G1341), .Z(new_n1013));
  NAND3_X1  g588(.A1(new_n997), .A2(new_n998), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n997), .A2(KEYINPUT121), .A3(new_n998), .A4(new_n1013), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n960), .A2(new_n931), .A3(new_n961), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1012), .B1(new_n1019), .B2(new_n552), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1019), .A2(new_n1012), .A3(new_n552), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1009), .B(new_n1011), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n992), .A2(new_n1002), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n595), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n992), .A2(new_n602), .A3(new_n1002), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1006), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT122), .B(G1961), .Z(new_n1029));
  NAND3_X1  g604(.A1(new_n985), .A2(new_n991), .A3(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n994), .B(new_n961), .C1(new_n980), .C2(KEYINPUT45), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(G2078), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n960), .A2(new_n747), .A3(new_n961), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1032), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT123), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(KEYINPUT123), .A3(new_n1032), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1033), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1030), .A2(new_n1039), .A3(G301), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT125), .B(G2078), .Z(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(new_n1032), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n960), .A2(KEYINPUT124), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n960), .A2(KEYINPUT124), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n961), .B(new_n1043), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n989), .B(KEYINPUT120), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1029), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT54), .B(new_n1040), .C1(new_n1049), .C2(new_n885), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  INV_X1    g626(.A(G1981), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n577), .A2(new_n1052), .A3(new_n578), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n577), .B2(new_n578), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n577), .A2(new_n1052), .A3(new_n578), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(KEYINPUT49), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n995), .A2(KEYINPUT115), .A3(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n995), .A2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1059), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1063), .A2(new_n1060), .B1(G1976), .B2(new_n684), .ZN(new_n1065));
  INV_X1    g640(.A(G1976), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(G288), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1064), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1065), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n684), .A2(G1976), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1060), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT115), .B1(new_n995), .B2(G8), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT116), .B1(new_n1075), .B2(KEYINPUT52), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1068), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G8), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n988), .A2(new_n982), .ZN(new_n1079));
  INV_X1    g654(.A(G2090), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n975), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1971), .B1(new_n960), .B2(new_n961), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1078), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT112), .B(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G303), .A2(G8), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1085), .ZN(new_n1089));
  NAND4_X1  g664(.A1(G303), .A2(KEYINPUT55), .A3(G8), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT114), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1084), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1092), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1082), .B1(new_n970), .B2(new_n1080), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1078), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1077), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G2084), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1079), .A2(new_n1100), .A3(new_n975), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1031), .A2(new_n732), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(G168), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G8), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT51), .ZN(new_n1105));
  AOI21_X1  g680(.A(G168), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  OAI211_X1 g682(.A(G8), .B(new_n1103), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1050), .A2(new_n1099), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1047), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1112), .A2(new_n1030), .A3(G301), .ZN(new_n1113));
  AOI21_X1  g688(.A(G301), .B1(new_n1030), .B2(new_n1039), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1028), .A2(new_n1110), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1117));
  NAND2_X1  g692(.A1(G168), .A2(G8), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1117), .B(new_n1119), .C1(new_n1084), .C2(new_n1092), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT63), .B1(new_n1077), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1097), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1094), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1063), .A2(new_n1060), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(new_n1072), .A3(new_n1067), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1058), .B(new_n1055), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1069), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1075), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(G288), .A2(G1976), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1057), .B1(new_n1064), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT117), .B(new_n1057), .C1(new_n1064), .C2(new_n1135), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n1126), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1121), .A2(new_n1133), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1105), .A2(new_n1108), .A3(new_n1142), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1096), .A2(new_n1078), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1084), .A2(new_n1093), .B1(new_n1144), .B2(new_n1095), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1132), .A2(new_n1114), .A3(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1109), .A2(KEYINPUT62), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1141), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g724(.A(KEYINPUT126), .B(new_n959), .C1(new_n1116), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1105), .A2(new_n1108), .A3(new_n1142), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1148), .A2(new_n1114), .A3(new_n1099), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1141), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1005), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n973), .B1(new_n1025), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1021), .A2(new_n1020), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n973), .A2(new_n1005), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n973), .A2(KEYINPUT61), .A3(new_n1005), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1011), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1026), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT60), .B1(new_n1164), .B2(new_n1003), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1156), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1115), .A2(new_n1050), .A3(new_n1099), .A4(new_n1109), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1153), .B(new_n1154), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n959), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1151), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n952), .B1(new_n1150), .B2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g746(.A1(G401), .A2(G229), .A3(new_n459), .A4(G227), .ZN(new_n1173));
  OAI21_X1  g747(.A(new_n1173), .B1(new_n848), .B2(new_n851), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n912), .A2(new_n913), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1175), .ZN(G308));
  AND2_X1   g750(.A1(new_n912), .A2(new_n913), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n836), .A2(new_n842), .A3(new_n841), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n1177), .A2(new_n1178), .A3(new_n1173), .ZN(G225));
endmodule


