//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(G134), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G122), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G116), .ZN(new_n198));
  INV_X1    g012(.A(G116), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G122), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(KEYINPUT14), .A3(G122), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(G107), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n200), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT93), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n198), .A2(new_n200), .A3(KEYINPUT93), .A4(new_n205), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n196), .A2(new_n204), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n198), .A2(new_n200), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT13), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n189), .A2(KEYINPUT13), .A3(G143), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G134), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n216), .A3(new_n195), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT94), .ZN(new_n219));
  XOR2_X1   g033(.A(KEYINPUT9), .B(G234), .Z(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G217), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT94), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n210), .A2(new_n217), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G902), .ZN(new_n226));
  INV_X1    g040(.A(new_n222), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n218), .A2(KEYINPUT94), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G478), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT15), .ZN(new_n231));
  XOR2_X1   g045(.A(new_n229), .B(new_n231), .Z(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G953), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT66), .B(G237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G214), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT88), .A2(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT18), .A2(G131), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n242), .A2(KEYINPUT89), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT88), .A2(G143), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n237), .A2(new_n245), .A3(new_n238), .A4(G214), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n241), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n242), .A2(KEYINPUT89), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G125), .ZN(new_n250));
  INV_X1    g064(.A(G140), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(G125), .A2(G140), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n241), .A2(KEYINPUT89), .A3(new_n242), .A4(new_n246), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n249), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n241), .A2(G131), .A3(new_n246), .ZN(new_n259));
  AOI21_X1  g073(.A(G131), .B1(new_n241), .B2(new_n246), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT17), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT16), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n262), .B1(new_n252), .B2(new_n253), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n251), .A3(G125), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n255), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n253), .ZN(new_n267));
  NOR2_X1   g081(.A1(G125), .A2(G140), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT16), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(G146), .A3(new_n264), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(KEYINPUT74), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n263), .A2(new_n265), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(G146), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT17), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n241), .A2(G131), .A3(new_n246), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n258), .B1(new_n261), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(G113), .B(G122), .Z(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT91), .ZN(new_n281));
  INV_X1    g095(.A(G104), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n283), .B(new_n258), .C1(new_n261), .C2(new_n278), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT92), .B1(new_n287), .B2(new_n226), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT92), .ZN(new_n289));
  AOI211_X1 g103(.A(new_n289), .B(G902), .C1(new_n285), .C2(new_n286), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n233), .B1(new_n291), .B2(G475), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT95), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n270), .B(KEYINPUT75), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n254), .B(KEYINPUT19), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n255), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n294), .B(new_n296), .C1(new_n259), .C2(new_n260), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n258), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n283), .B1(new_n298), .B2(KEYINPUT90), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT90), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n258), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n286), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT20), .ZN(new_n304));
  NOR2_X1   g118(.A1(G475), .A2(G902), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n286), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(new_n299), .B2(new_n301), .ZN(new_n308));
  INV_X1    g122(.A(new_n305), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT20), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G952), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G953), .ZN(new_n313));
  NAND2_X1  g127(.A1(G234), .A2(G237), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n237), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n317), .A2(G902), .A3(new_n314), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT21), .B(G898), .Z(new_n320));
  OAI21_X1  g134(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n292), .A2(new_n293), .A3(new_n311), .A4(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  INV_X1    g137(.A(new_n240), .ZN(new_n324));
  OR2_X1    g138(.A1(KEYINPUT66), .A2(G237), .ZN(new_n325));
  NAND2_X1  g139(.A1(KEYINPUT66), .A2(G237), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n234), .A2(new_n236), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n324), .B1(new_n327), .B2(G214), .ZN(new_n328));
  INV_X1    g142(.A(new_n246), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n323), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n276), .A3(new_n277), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n259), .A2(KEYINPUT17), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n275), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n283), .B1(new_n333), .B2(new_n258), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n226), .B1(new_n307), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n289), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n287), .A2(KEYINPUT92), .A3(new_n226), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(G475), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n232), .A3(new_n321), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n308), .A2(KEYINPUT20), .A3(new_n309), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT95), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n322), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n237), .A2(G221), .A3(G234), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT22), .B(G137), .Z(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n189), .B2(G119), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n353));
  INV_X1    g167(.A(G119), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(G128), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(KEYINPUT73), .A3(G128), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n189), .A2(KEYINPUT72), .A3(G119), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n352), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT24), .B(G110), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n354), .A2(G128), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT23), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT23), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n354), .B2(G128), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n362), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n360), .B1(G110), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n270), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n272), .A2(KEYINPUT75), .A3(G146), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n254), .A2(new_n255), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n366), .A2(new_n368), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n358), .A2(new_n359), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n365), .A2(G110), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n271), .A2(new_n274), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT78), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n371), .B2(new_n374), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n350), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n378), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n349), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G217), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(G234), .B2(new_n226), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G902), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n385), .B(KEYINPUT79), .Z(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT80), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n379), .A2(new_n226), .A3(new_n381), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT25), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT25), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n379), .A2(new_n391), .A3(new_n226), .A4(new_n381), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n384), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n382), .A2(new_n394), .A3(new_n386), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT11), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n194), .B2(G137), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n194), .A2(G137), .ZN(new_n399));
  INV_X1    g213(.A(G137), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT11), .A3(G134), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G131), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n398), .A2(new_n401), .A3(new_n323), .A4(new_n399), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n255), .A2(G143), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n187), .A2(G146), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT0), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n189), .ZN(new_n410));
  NAND2_X1  g224(.A1(KEYINPUT0), .A2(G128), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n406), .A2(new_n407), .A3(new_n411), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n405), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT2), .B(G113), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G116), .B(G119), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(G116), .B(G119), .Z(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n417), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n406), .A3(new_n407), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n189), .A2(new_n255), .A3(G143), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n187), .B(G146), .C1(new_n189), .C2(KEYINPUT1), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT65), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n400), .A3(G134), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n399), .A2(KEYINPUT65), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n194), .A2(G137), .ZN(new_n433));
  OAI211_X1 g247(.A(G131), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n434), .A3(new_n404), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n416), .A2(new_n424), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT28), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n436), .A2(KEYINPUT70), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT70), .B1(new_n436), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT71), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT70), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n429), .A2(new_n434), .A3(new_n404), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n403), .A2(new_n404), .B1(new_n413), .B2(new_n414), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n442), .A2(new_n443), .A3(new_n423), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n444), .B2(KEYINPUT28), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n436), .A2(KEYINPUT70), .A3(new_n437), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n424), .B1(new_n416), .B2(new_n435), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT28), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT29), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n237), .A2(new_n238), .A3(G210), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT26), .B(G101), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n406), .A2(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n406), .A2(new_n407), .A3(new_n411), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT64), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n405), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n424), .B1(new_n463), .B2(new_n435), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT69), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n436), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(KEYINPUT69), .B(new_n424), .C1(new_n463), .C2(new_n435), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT28), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n438), .A2(new_n439), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT29), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n452), .A2(new_n457), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n416), .A2(KEYINPUT30), .A3(new_n435), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n459), .A2(new_n460), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n474), .A2(KEYINPUT64), .B1(new_n403), .B2(new_n404), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n442), .B1(new_n475), .B2(new_n461), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n423), .B(new_n473), .C1(new_n476), .C2(KEYINPUT30), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n477), .A2(new_n436), .ZN(new_n478));
  INV_X1    g292(.A(new_n457), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n470), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n472), .A2(new_n226), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G472), .ZN(new_n484));
  NOR2_X1   g298(.A1(G472), .A2(G902), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n477), .A2(new_n436), .A3(new_n457), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT31), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT31), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n477), .A2(new_n488), .A3(new_n436), .A4(new_n457), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n457), .B1(new_n468), .B2(new_n469), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n485), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT32), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n494), .B(new_n485), .C1(new_n490), .C2(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n396), .B1(new_n484), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n220), .A2(new_n226), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n498), .A2(G221), .ZN(new_n499));
  INV_X1    g313(.A(G469), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(new_n226), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n237), .A2(G227), .ZN(new_n502));
  XNOR2_X1  g316(.A(G110), .B(G140), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT81), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n506), .A2(KEYINPUT3), .B1(new_n282), .B2(G107), .ZN(new_n507));
  OAI22_X1  g321(.A1(new_n506), .A2(KEYINPUT3), .B1(new_n282), .B2(G107), .ZN(new_n508));
  INV_X1    g322(.A(G101), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT3), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(new_n205), .A3(KEYINPUT81), .A4(G104), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n205), .A2(G104), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n282), .A2(G107), .ZN(new_n514));
  OAI21_X1  g328(.A(G101), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n429), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n429), .B1(new_n512), .B2(new_n515), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT12), .B(new_n405), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT84), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n403), .A2(new_n404), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n512), .A2(new_n515), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n521), .B1(new_n524), .B2(new_n516), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT12), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n405), .B1(new_n517), .B2(new_n518), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n520), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n509), .A2(KEYINPUT82), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT4), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(KEYINPUT4), .A3(new_n533), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n512), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n415), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n517), .A2(KEYINPUT10), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT10), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n516), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n405), .A2(KEYINPUT83), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT83), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n403), .B2(new_n404), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n539), .A2(new_n540), .A3(new_n542), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n531), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n547), .A2(new_n504), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n538), .A2(new_n415), .B1(new_n541), .B2(new_n516), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n521), .B1(new_n550), .B2(new_n540), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n505), .A2(new_n548), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n501), .B1(new_n553), .B2(G469), .ZN(new_n554));
  INV_X1    g368(.A(new_n547), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n505), .B1(new_n555), .B2(new_n551), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n531), .A2(new_n547), .A3(new_n504), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n500), .A3(new_n226), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n499), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G214), .B1(G237), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT87), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n474), .A2(G125), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n523), .A2(new_n250), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G224), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n563), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n566), .B(new_n569), .C1(KEYINPUT87), .C2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(KEYINPUT87), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n568), .B1(new_n572), .B2(new_n565), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT5), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n354), .A3(G116), .ZN(new_n576));
  OAI211_X1 g390(.A(G113), .B(new_n576), .C1(new_n421), .C2(new_n575), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n577), .A2(new_n420), .A3(new_n512), .A4(new_n515), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT85), .ZN(new_n579));
  INV_X1    g393(.A(new_n522), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT85), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n420), .A4(new_n577), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n532), .A2(KEYINPUT4), .A3(new_n533), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT4), .B1(new_n532), .B2(new_n533), .ZN(new_n584));
  INV_X1    g398(.A(new_n512), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n579), .B(new_n582), .C1(new_n586), .C2(new_n424), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT6), .ZN(new_n588));
  XOR2_X1   g402(.A(G110), .B(G122), .Z(new_n589));
  NAND4_X1  g403(.A1(new_n587), .A2(KEYINPUT86), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n587), .A2(KEYINPUT86), .A3(new_n589), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n538), .A2(new_n423), .ZN(new_n592));
  INV_X1    g406(.A(new_n589), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n579), .A4(new_n582), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT6), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n574), .B(new_n590), .C1(new_n591), .C2(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n572), .A2(new_n565), .A3(new_n568), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n563), .A2(new_n564), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n569), .A2(KEYINPUT7), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n597), .A2(KEYINPUT7), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n589), .B(KEYINPUT8), .Z(new_n601));
  AOI21_X1  g415(.A(new_n580), .B1(new_n420), .B2(new_n577), .ZN(new_n602));
  INV_X1    g416(.A(new_n578), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n600), .A2(new_n594), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n596), .A2(new_n605), .A3(new_n226), .ZN(new_n606));
  OAI21_X1  g420(.A(G210), .B1(G237), .B2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n596), .A2(new_n605), .A3(new_n226), .A4(new_n607), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n560), .A2(new_n561), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n344), .A2(new_n497), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  INV_X1    g428(.A(new_n499), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n548), .A2(new_n505), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n549), .A2(new_n552), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n500), .B1(new_n618), .B2(new_n226), .ZN(new_n619));
  AOI211_X1 g433(.A(G469), .B(G902), .C1(new_n556), .C2(new_n557), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n396), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n226), .B1(new_n490), .B2(new_n491), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G472), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n624), .A2(new_n492), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n561), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n609), .B2(new_n610), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n628), .A2(new_n321), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT33), .B1(new_n225), .B2(new_n228), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n222), .A2(KEYINPUT96), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n218), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n218), .A2(new_n633), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(G478), .B(new_n226), .C1(new_n631), .C2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT97), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n229), .A2(new_n230), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n311), .A2(new_n338), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n630), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT34), .B(G104), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NAND2_X1  g459(.A1(new_n338), .A2(new_n233), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n311), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n306), .A2(new_n310), .A3(KEYINPUT98), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n626), .A2(new_n629), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT35), .B(G107), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT99), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n651), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n350), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n375), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n386), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n393), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n344), .A2(new_n612), .A3(new_n625), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT37), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(G110), .Z(G12));
  AND2_X1   g475(.A1(new_n393), .A2(new_n657), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n484), .B2(new_n496), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n316), .B1(new_n319), .B2(G900), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT100), .Z(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n663), .A2(new_n612), .A3(new_n650), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XOR2_X1   g482(.A(new_n665), .B(KEYINPUT39), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n560), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT101), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT40), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n611), .B(KEYINPUT38), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n233), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n444), .A2(new_n449), .ZN(new_n676));
  AOI21_X1  g490(.A(G902), .B1(new_n479), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n478), .B2(new_n479), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n678), .A2(G472), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n493), .B2(new_n495), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n675), .A2(new_n680), .A3(new_n658), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n672), .A2(new_n561), .A3(new_n673), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT102), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n187), .ZN(G45));
  NAND2_X1  g498(.A1(new_n639), .A2(new_n640), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n674), .A2(new_n685), .A3(new_n666), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n663), .A2(new_n686), .A3(new_n612), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  AOI21_X1  g502(.A(new_n500), .B1(new_n558), .B2(new_n226), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n620), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n615), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n497), .A2(new_n629), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n642), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT41), .B(G113), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NAND4_X1  g510(.A1(new_n497), .A2(new_n629), .A3(new_n650), .A4(new_n692), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  AND4_X1   g512(.A1(new_n561), .A2(new_n611), .A3(new_n690), .A4(new_n615), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n344), .A2(new_n663), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT103), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n344), .A2(new_n702), .A3(new_n663), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  XOR2_X1   g519(.A(KEYINPUT104), .B(G472), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n623), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n451), .A2(new_n479), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n485), .B1(new_n708), .B2(new_n490), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n691), .A2(new_n710), .A3(new_n396), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n675), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n674), .A2(KEYINPUT105), .A3(new_n233), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n711), .A2(new_n713), .A3(new_n629), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT106), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n197), .ZN(G24));
  NOR2_X1   g531(.A1(new_n710), .A2(new_n662), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n699), .A2(new_n686), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n609), .A2(new_n561), .A3(new_n610), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n621), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n497), .A2(new_n686), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT42), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT42), .B1(new_n724), .B2(new_n725), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n721), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n724), .A2(new_n725), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(KEYINPUT108), .A3(new_n726), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT109), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  INV_X1    g550(.A(new_n722), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n497), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n646), .ZN(new_n739));
  INV_X1    g553(.A(new_n649), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT98), .B1(new_n306), .B2(new_n310), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n739), .B(new_n666), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n560), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n685), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n674), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n311), .A2(KEYINPUT110), .A3(new_n338), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT110), .B1(new_n311), .B2(new_n338), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n685), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n748), .B1(new_n752), .B2(KEYINPUT43), .ZN(new_n753));
  INV_X1    g567(.A(new_n625), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n658), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n618), .B(KEYINPUT45), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(G469), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n759), .B(KEYINPUT46), .C1(new_n500), .C2(new_n226), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n761), .B(G469), .C1(new_n758), .C2(G902), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n559), .A3(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n763), .A2(new_n615), .A3(new_n669), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n755), .A2(new_n756), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n757), .A2(new_n737), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  NAND2_X1  g581(.A1(new_n484), .A2(new_n496), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n763), .A2(new_n769), .A3(new_n615), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n769), .B1(new_n763), .B2(new_n615), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT47), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n770), .B2(new_n771), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n768), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(new_n396), .A3(new_n686), .A4(new_n737), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  INV_X1    g592(.A(new_n690), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n561), .B(new_n615), .C1(new_n779), .C2(KEYINPUT49), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n780), .B(new_n752), .C1(KEYINPUT49), .C2(new_n779), .ZN(new_n781));
  INV_X1    g595(.A(new_n396), .ZN(new_n782));
  INV_X1    g596(.A(new_n673), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .A4(new_n680), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n783), .A2(new_n711), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n747), .A2(new_n674), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n674), .A2(new_n788), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n789), .A2(new_n749), .B1(new_n640), .B2(new_n639), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n315), .B(new_n787), .C1(new_n790), .C2(new_n746), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(KEYINPUT116), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(KEYINPUT116), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n627), .B(new_n786), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n691), .A2(new_n722), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n782), .A3(new_n315), .A4(new_n680), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n674), .A3(new_n685), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n718), .B(new_n797), .C1(new_n792), .C2(new_n793), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n791), .B(KEYINPUT116), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(KEYINPUT117), .A3(new_n718), .A4(new_n797), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n799), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT118), .B1(new_n796), .B2(new_n805), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n782), .A2(new_n803), .A3(new_n709), .A4(new_n707), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n690), .A2(new_n499), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n773), .A2(new_n775), .A3(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n807), .A2(new_n737), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n785), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n803), .A2(new_n497), .A3(new_n797), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n803), .A2(KEYINPUT120), .A3(new_n497), .A4(new_n797), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(KEYINPUT48), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n807), .A2(new_n699), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n313), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n814), .A2(KEYINPUT48), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n342), .A2(new_n646), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n629), .A2(new_n625), .A3(new_n622), .A4(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n659), .A2(new_n613), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n648), .A2(new_n649), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n768), .A2(new_n723), .A3(new_n824), .A4(new_n666), .ZN(new_n825));
  INV_X1    g639(.A(new_n292), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n641), .A2(new_n737), .A3(new_n560), .A4(new_n666), .ZN(new_n827));
  OAI22_X1  g641(.A1(new_n825), .A2(new_n826), .B1(new_n710), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n658), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n674), .A2(new_n685), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n674), .B2(new_n685), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n629), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT113), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n629), .B(new_n835), .C1(new_n831), .C2(new_n832), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n626), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n823), .A2(new_n829), .A3(new_n837), .A4(new_n744), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n667), .A2(new_n687), .A3(new_n719), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n713), .A2(new_n628), .A3(new_n714), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n615), .B(new_n666), .C1(new_n619), .C2(new_n620), .ZN(new_n841));
  OR3_X1    g655(.A1(new_n680), .A2(new_n841), .A3(new_n658), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT114), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n612), .B(new_n663), .C1(new_n743), .C2(new_n686), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n680), .A2(new_n841), .A3(new_n658), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n628), .A3(new_n713), .A4(new_n714), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(new_n846), .A3(new_n719), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n839), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(KEYINPUT52), .A3(new_n848), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n838), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n727), .A2(new_n728), .A3(new_n721), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT108), .B1(new_n732), .B2(new_n726), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n694), .B1(new_n701), .B2(new_n703), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n715), .A2(new_n697), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n854), .A2(new_n855), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n744), .A2(new_n823), .A3(new_n829), .A4(new_n837), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n858), .A2(new_n863), .A3(new_n861), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n844), .A2(new_n850), .A3(new_n849), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n850), .B1(new_n844), .B2(new_n849), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n862), .B(KEYINPUT54), .C1(new_n868), .C2(new_n855), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n855), .B1(new_n864), .B2(new_n867), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n727), .A2(new_n728), .ZN(new_n871));
  AND4_X1   g685(.A1(KEYINPUT53), .A2(new_n871), .A3(new_n860), .A4(new_n859), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n854), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g687(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n811), .A2(new_n820), .A3(new_n869), .A4(new_n876), .ZN(new_n877));
  OR2_X1    g691(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n773), .A2(new_n879), .A3(new_n775), .A4(new_n808), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(KEYINPUT51), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n809), .A2(KEYINPUT119), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n737), .A3(new_n882), .A4(new_n807), .ZN(new_n883));
  AND4_X1   g697(.A1(new_n878), .A2(new_n883), .A3(new_n796), .A4(new_n805), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n798), .A2(new_n642), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n877), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(G952), .A2(G953), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n784), .B1(new_n886), .B2(new_n887), .ZN(G75));
  AOI21_X1  g702(.A(new_n226), .B1(new_n870), .B2(new_n873), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G210), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n590), .B1(new_n591), .B2(new_n595), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(new_n574), .Z(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(KEYINPUT121), .B2(KEYINPUT56), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n890), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n890), .B2(new_n891), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n317), .A2(new_n312), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT122), .Z(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(G51));
  XNOR2_X1  g715(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n501), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n859), .A2(new_n860), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n734), .A2(new_n838), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n844), .A2(new_n849), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT52), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n851), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT53), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n851), .A2(new_n853), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n872), .A2(new_n910), .A3(new_n863), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n909), .A2(new_n911), .A3(new_n874), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n875), .B1(new_n870), .B2(new_n873), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT124), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n916), .B(new_n903), .C1(new_n912), .C2(new_n913), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n558), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n889), .A2(G469), .A3(new_n758), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n900), .B1(new_n918), .B2(new_n919), .ZN(G54));
  NAND3_X1  g734(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(new_n303), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n303), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n900), .B1(new_n922), .B2(new_n923), .ZN(G60));
  NOR2_X1   g738(.A1(new_n631), .A2(new_n636), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n869), .A2(new_n876), .ZN(new_n926));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT59), .Z(new_n928));
  OAI21_X1  g742(.A(new_n925), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n928), .ZN(new_n930));
  OAI221_X1 g744(.A(new_n930), .B1(new_n636), .B2(new_n631), .C1(new_n912), .C2(new_n913), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n929), .A2(new_n931), .A3(new_n899), .ZN(G63));
  NAND2_X1  g746(.A1(new_n870), .A2(new_n873), .ZN(new_n933));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n382), .B(KEYINPUT126), .Z(new_n938));
  AOI21_X1  g752(.A(new_n900), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT61), .B1(new_n939), .B2(KEYINPUT125), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n933), .A2(new_n656), .A3(new_n936), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n939), .B(new_n941), .C1(KEYINPUT125), .C2(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(G66));
  AOI21_X1  g759(.A(new_n221), .B1(new_n320), .B2(G224), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n861), .A2(new_n823), .A3(new_n837), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n237), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n892), .B1(G898), .B2(new_n237), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(G69));
  NAND3_X1  g764(.A1(new_n777), .A2(new_n766), .A3(new_n852), .ZN(new_n951));
  INV_X1    g765(.A(new_n840), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n764), .A2(new_n497), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n858), .A2(new_n744), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n237), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n473), .B1(new_n476), .B2(KEYINPUT30), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n295), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n955), .B(new_n958), .C1(G227), .C2(new_n237), .ZN(new_n959));
  OAI21_X1  g773(.A(G900), .B1(new_n958), .B2(G227), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n317), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n682), .A2(new_n852), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n682), .A2(KEYINPUT62), .A3(new_n852), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OR3_X1    g780(.A1(new_n831), .A2(new_n832), .A3(new_n821), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n968), .A2(new_n671), .A3(new_n738), .A4(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n966), .A2(new_n777), .A3(new_n766), .A4(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n237), .A3(new_n957), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n959), .A2(new_n961), .A3(new_n972), .ZN(G72));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n971), .B2(new_n947), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n478), .A2(new_n479), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n900), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n951), .A2(new_n947), .A3(new_n954), .ZN(new_n979));
  INV_X1    g793(.A(new_n975), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n481), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n862), .B1(new_n868), .B2(new_n855), .ZN(new_n982));
  OR3_X1    g796(.A1(new_n982), .A2(new_n481), .A3(new_n977), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n978), .B(new_n981), .C1(new_n983), .C2(new_n980), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(G57));
endmodule


