//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n473), .A2(new_n475), .A3(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n468), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n472), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(new_n475), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n480), .B1(new_n474), .B2(KEYINPUT3), .ZN(new_n481));
  AND2_X1   g056(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n479), .A2(G137), .A3(new_n481), .A4(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n474), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G101), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n477), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  OAI221_X1 g064(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n484), .C2(G112), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n481), .A2(new_n475), .A3(new_n478), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n468), .ZN(new_n492));
  INV_X1    g067(.A(G124), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n481), .A2(new_n475), .A3(new_n478), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n494), .B1(G136), .B2(new_n496), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n466), .A2(G138), .A3(new_n467), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n473), .A2(new_n475), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT4), .A2(G138), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n484), .A2(new_n507), .B1(G126), .B2(G2105), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n501), .B(new_n505), .C1(new_n508), .C2(new_n495), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(KEYINPUT70), .B1(new_n515), .B2(G62), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n516), .B1(G75), .B2(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(KEYINPUT70), .A3(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n512), .B1(new_n522), .B2(new_n523), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT69), .A3(G50), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n524), .A2(new_n515), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n527), .A2(new_n529), .B1(G88), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n520), .A2(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n513), .A2(new_n514), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n524), .A2(G89), .ZN(new_n538));
  NAND2_X1  g113(.A1(G63), .A2(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n536), .A2(new_n540), .ZN(G168));
  AOI22_X1  g116(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n528), .A2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n530), .A2(G90), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n524), .A2(new_n515), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n542), .A2(new_n543), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT71), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n548), .A2(new_n553), .ZN(G171));
  NAND2_X1  g129(.A1(new_n528), .A2(G43), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT73), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT74), .ZN(G188));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n530), .A2(new_n569), .A3(G91), .ZN(new_n570));
  INV_X1    g145(.A(G91), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT76), .B1(new_n549), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n525), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n528), .A2(new_n573), .A3(new_n576), .A4(G53), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n570), .A2(new_n572), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G65), .ZN(new_n579));
  INV_X1    g154(.A(G78), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n537), .A2(new_n579), .B1(new_n580), .B2(new_n512), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI221_X1 g158(.A(KEYINPUT77), .B1(new_n580), .B2(new_n512), .C1(new_n537), .C2(new_n579), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n583), .A2(G651), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n578), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  INV_X1    g162(.A(G168), .ZN(G286));
  NAND2_X1  g163(.A1(new_n520), .A2(new_n531), .ZN(G303));
  NAND2_X1  g164(.A1(new_n528), .A2(G49), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n530), .A2(G87), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G288));
  AOI22_X1  g169(.A1(new_n530), .A2(G86), .B1(G48), .B2(new_n528), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n537), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n598), .A2(KEYINPUT78), .A3(G651), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n543), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n603), .B1(new_n599), .B2(new_n602), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n595), .B1(new_n604), .B2(new_n605), .ZN(G305));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT80), .B(G47), .Z(new_n608));
  OAI22_X1  g183(.A1(new_n549), .A2(new_n607), .B1(new_n525), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n543), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G290));
  NAND3_X1  g188(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n549), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n537), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g200(.A(new_n624), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(G299), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G297));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G280));
  AND2_X1   g205(.A1(new_n618), .A2(new_n622), .ZN(new_n631));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G860), .ZN(G148));
  NOR2_X1   g208(.A1(new_n560), .A2(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n632), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G868), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n496), .A2(G135), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n484), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n495), .A2(new_n484), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n642), .A2(KEYINPUT82), .A3(G123), .ZN(new_n643));
  AOI21_X1  g218(.A(KEYINPUT82), .B1(new_n642), .B2(G123), .ZN(new_n644));
  OAI221_X1 g219(.A(new_n639), .B1(new_n640), .B2(new_n641), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  INV_X1    g230(.A(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n655), .A2(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT83), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT14), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n655), .B(G2430), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n666), .B1(new_n667), .B2(new_n658), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n669), .A3(new_n660), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2451), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT16), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  AND3_X1   g249(.A1(new_n665), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n665), .B2(new_n670), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n654), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n674), .ZN(new_n678));
  INV_X1    g253(.A(new_n670), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n669), .B1(new_n668), .B2(new_n660), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n665), .A2(new_n670), .A3(new_n674), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n653), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n677), .A2(G14), .A3(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G401));
  XNOR2_X1  g260(.A(KEYINPUT85), .B(G2096), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2084), .B(G2090), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G2072), .A2(G2078), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n443), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT17), .ZN(new_n696));
  INV_X1    g271(.A(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n688), .A3(new_n691), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT18), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n697), .A2(KEYINPUT18), .A3(new_n691), .A4(new_n688), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n693), .A2(new_n696), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G2100), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n688), .B(KEYINPUT84), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(new_n695), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n705), .B(new_n692), .C1(new_n704), .C2(new_n696), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n703), .B1(new_n702), .B2(new_n706), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n687), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n700), .A2(new_n701), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n696), .A2(new_n704), .A3(new_n691), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n705), .A2(new_n692), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n696), .A2(new_n704), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n710), .B(new_n711), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G2100), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n702), .A2(new_n706), .A3(new_n703), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n715), .A2(new_n686), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n709), .A2(new_n717), .ZN(G227));
  XOR2_X1   g293(.A(G1991), .B(G1996), .Z(new_n719));
  XNOR2_X1  g294(.A(G1956), .B(G2474), .ZN(new_n720));
  XNOR2_X1  g295(.A(G1961), .B(G1966), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  INV_X1    g298(.A(G1971), .ZN(new_n724));
  INV_X1    g299(.A(G1976), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(G1971), .A2(G1976), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT19), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n726), .A2(KEYINPUT19), .A3(new_n727), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(new_n722), .B(new_n723), .S(new_n732), .Z(new_n733));
  NOR2_X1   g308(.A1(new_n720), .A2(new_n721), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT20), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT20), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n732), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n733), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n733), .B2(new_n739), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n719), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(G1981), .B(G1986), .ZN(new_n744));
  INV_X1    g319(.A(new_n740), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n736), .A2(new_n738), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n732), .A2(new_n720), .A3(new_n721), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n722), .B2(new_n732), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n719), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n733), .A2(new_n739), .A3(new_n740), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n743), .A2(new_n744), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n744), .B1(new_n743), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(G229));
  INV_X1    g330(.A(G34), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n756), .B2(KEYINPUT24), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(KEYINPUT24), .B2(new_n756), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n488), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT93), .ZN(new_n763));
  INV_X1    g338(.A(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G5), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G171), .B2(new_n764), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n763), .B1(G1961), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n759), .A2(G32), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT26), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n773), .A2(new_n774), .B1(G105), .B2(new_n486), .ZN(new_n775));
  INV_X1    g350(.A(G129), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n492), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n496), .A2(G141), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n770), .B1(new_n779), .B2(new_n759), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT90), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n767), .B1(new_n769), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT94), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT31), .B(G11), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n759), .B1(new_n785), .B2(G28), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(KEYINPUT91), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(G28), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n786), .B2(KEYINPUT91), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G19), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n560), .B2(G16), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n784), .B1(new_n787), .B2(new_n789), .C1(new_n791), .C2(G1341), .ZN(new_n792));
  NOR2_X1   g367(.A1(G168), .A2(new_n764), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n764), .B2(G21), .ZN(new_n794));
  INV_X1    g369(.A(G1966), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n792), .B(new_n796), .C1(G1341), .C2(new_n791), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n795), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(KEYINPUT92), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n759), .A2(G33), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT25), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n496), .A2(G139), .ZN(new_n803));
  NAND2_X1  g378(.A1(G115), .A2(G2104), .ZN(new_n804));
  INV_X1    g379(.A(G127), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n500), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(new_n468), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n802), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n800), .B1(new_n809), .B2(new_n759), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n799), .B1(G2072), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n759), .A2(G35), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT95), .Z(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n759), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT29), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G2090), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n766), .A2(G1961), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n797), .A2(new_n811), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n815), .A2(G2090), .B1(new_n781), .B2(new_n769), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n764), .A2(G20), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT23), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n628), .B2(new_n764), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT96), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1956), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n798), .A2(KEYINPUT92), .ZN(new_n826));
  INV_X1    g401(.A(G1348), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n764), .A2(G4), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n623), .B2(G16), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n826), .B1(new_n759), .B2(new_n645), .C1(new_n827), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(G164), .A2(new_n759), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G27), .B2(new_n759), .ZN(new_n832));
  INV_X1    g407(.A(G2078), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n832), .A2(new_n833), .B1(new_n827), .B2(new_n829), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n834), .B1(new_n833), .B2(new_n832), .C1(new_n810), .C2(G2072), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n760), .A2(new_n761), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT89), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n759), .A2(G26), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT28), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n496), .A2(G140), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n642), .A2(G128), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(G116), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n468), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT88), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI211_X1 g421(.A(KEYINPUT88), .B(new_n842), .C1(new_n468), .C2(new_n843), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n840), .B(new_n841), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n839), .B1(new_n848), .B2(G29), .ZN(new_n849));
  INV_X1    g424(.A(G2067), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NOR4_X1   g426(.A1(new_n830), .A2(new_n835), .A3(new_n837), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n783), .A2(new_n820), .A3(new_n825), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n764), .A2(G23), .ZN(new_n854));
  INV_X1    g429(.A(G288), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n764), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT33), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G1976), .ZN(new_n858));
  MUX2_X1   g433(.A(G6), .B(G305), .S(G16), .Z(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT32), .B(G1981), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  NOR2_X1   g437(.A1(G16), .A2(G22), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G166), .B2(G16), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n724), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n858), .A2(new_n861), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT34), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(KEYINPUT34), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n496), .A2(G131), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n642), .A2(G119), .ZN(new_n870));
  OAI221_X1 g445(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n484), .C2(G107), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT86), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT86), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n869), .A2(new_n870), .A3(new_n874), .A4(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G29), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(G25), .B2(G29), .ZN(new_n879));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G1991), .Z(new_n880));
  AND2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n764), .A2(G24), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n612), .B2(new_n764), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G1986), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n867), .A2(new_n868), .A3(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(KEYINPUT87), .B(KEYINPUT36), .Z(new_n888));
  AOI21_X1  g463(.A(new_n853), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n889), .A2(new_n891), .A3(KEYINPUT97), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT97), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(G311));
  AND3_X1   g469(.A1(new_n889), .A2(new_n891), .A3(KEYINPUT98), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT98), .B1(new_n889), .B2(new_n891), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(G150));
  NAND2_X1  g472(.A1(new_n528), .A2(G55), .ZN(new_n898));
  INV_X1    g473(.A(G93), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n549), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G67), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n513), .B2(new_n514), .ZN(new_n902));
  AND2_X1   g477(.A1(G80), .A2(G543), .ZN(new_n903));
  OAI21_X1  g478(.A(G651), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT99), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n530), .A2(G93), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n904), .A4(new_n898), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n560), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n904), .A3(new_n898), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n911), .B(KEYINPUT99), .C1(new_n559), .C2(new_n557), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(KEYINPUT38), .Z(new_n914));
  NAND2_X1  g489(.A1(new_n631), .A2(G559), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n916), .A2(KEYINPUT39), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(KEYINPUT39), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n917), .A2(new_n918), .A3(G860), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n911), .A2(G860), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT37), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n919), .A2(new_n921), .ZN(G145));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n479), .A2(new_n465), .A3(new_n481), .ZN(new_n925));
  INV_X1    g500(.A(G142), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n496), .A2(KEYINPUT100), .A3(G142), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n930));
  INV_X1    g505(.A(G118), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n468), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n642), .B2(G130), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n649), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n649), .B1(new_n929), .B2(new_n933), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n935), .A2(new_n876), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n929), .A2(new_n933), .ZN(new_n938));
  INV_X1    g513(.A(new_n649), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n940), .A2(new_n934), .B1(new_n873), .B2(new_n875), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n923), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n877), .A2(new_n940), .A3(new_n934), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n876), .B1(new_n935), .B2(new_n936), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT101), .ZN(new_n945));
  INV_X1    g520(.A(new_n779), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n848), .A2(new_n509), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n848), .A2(new_n509), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n848), .A2(new_n509), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n779), .A3(new_n947), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n808), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n808), .B1(new_n950), .B2(new_n952), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n942), .B(new_n945), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(G162), .B(new_n488), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(new_n645), .Z(new_n958));
  INV_X1    g533(.A(new_n955), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT101), .B1(new_n943), .B2(new_n944), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n953), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G37), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n958), .B1(new_n956), .B2(new_n961), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g544(.A(KEYINPUT41), .ZN(new_n970));
  NAND2_X1  g545(.A1(G299), .A2(new_n631), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n623), .A2(new_n585), .A3(new_n578), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(KEYINPUT102), .A3(new_n972), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT102), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n628), .A2(new_n975), .A3(new_n623), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n973), .B1(new_n977), .B2(new_n970), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n913), .B(new_n635), .Z(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(new_n971), .B2(new_n972), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(KEYINPUT103), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n984), .B2(new_n980), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT104), .B1(new_n592), .B2(new_n593), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n592), .A2(KEYINPUT104), .A3(new_n593), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(G290), .A3(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n592), .A2(KEYINPUT104), .A3(new_n593), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n612), .B1(new_n992), .B2(new_n988), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n604), .A2(new_n605), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(G166), .A3(new_n595), .ZN(new_n996));
  NAND2_X1  g571(.A1(G305), .A2(G303), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n987), .B(new_n994), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n994), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n997), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n1000), .B2(KEYINPUT105), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n987), .A3(new_n997), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n986), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n986), .B2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g581(.A(G868), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n911), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1007), .B1(G868), .B2(new_n1008), .ZN(G295));
  OAI21_X1  g584(.A(new_n1007), .B1(G868), .B2(new_n1008), .ZN(G331));
  AND3_X1   g585(.A1(G171), .A2(new_n910), .A3(new_n912), .ZN(new_n1011));
  AOI21_X1  g586(.A(G171), .B1(new_n912), .B2(new_n910), .ZN(new_n1012));
  OAI21_X1  g587(.A(G286), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n913), .A2(G301), .ZN(new_n1014));
  NAND3_X1  g589(.A1(G171), .A2(new_n910), .A3(new_n912), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(G168), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n971), .A2(new_n972), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n978), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1013), .A2(new_n1016), .A3(KEYINPUT106), .A4(new_n1017), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G37), .B1(new_n1024), .B2(new_n1003), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1027));
  INV_X1    g602(.A(new_n998), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT43), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n963), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n977), .A2(KEYINPUT41), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n977), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1021), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1017), .A2(new_n970), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1018), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1003), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1032), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT44), .B1(new_n1031), .B2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1044), .A2(KEYINPUT106), .B1(new_n978), .B2(new_n1021), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1003), .B1(new_n1045), .B2(new_n1020), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT43), .B1(new_n1032), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1039), .A2(new_n1037), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1029), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1045), .A2(new_n1003), .A3(new_n1020), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n1041), .A4(new_n963), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1043), .B1(new_n1053), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g629(.A(G1384), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT45), .B1(new_n509), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n477), .A2(G40), .A3(new_n485), .A4(new_n487), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n877), .A2(new_n880), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n848), .B(new_n850), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n779), .B(G1996), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n877), .A2(new_n880), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(new_n612), .B(G1986), .Z(new_n1065));
  OAI21_X1  g640(.A(new_n1059), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n1055), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1067), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(G1971), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n509), .A2(new_n1055), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1058), .B1(new_n1070), .B2(KEYINPUT50), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G126), .A2(G2105), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n468), .B2(new_n506), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n504), .B1(new_n1073), .B2(new_n491), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1384), .B1(new_n1074), .B2(new_n501), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1071), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(G2090), .ZN(new_n1079));
  OAI21_X1  g654(.A(G8), .B1(new_n1069), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(G303), .A2(G8), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1070), .A2(new_n1058), .ZN(new_n1087));
  INV_X1    g662(.A(G8), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1981), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n595), .C1(new_n604), .C2(new_n605), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n599), .A2(new_n595), .A3(new_n602), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G1981), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT109), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(KEYINPUT109), .A3(G1981), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1092), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n1099));
  AOI21_X1  g674(.A(new_n1090), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1092), .A2(new_n1096), .A3(KEYINPUT49), .A4(new_n1097), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1089), .B(KEYINPUT108), .C1(new_n725), .C2(G288), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n855), .A2(G1976), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(new_n1089), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1106), .B(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1086), .A2(new_n1105), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n469), .B(KEYINPUT67), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n473), .A2(new_n475), .A3(G125), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n484), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n466), .A2(G137), .A3(new_n467), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n495), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G40), .ZN(new_n1117));
  INV_X1    g692(.A(new_n487), .ZN(new_n1118));
  NOR4_X1   g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n509), .A2(new_n1076), .A3(new_n1055), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1120), .A2(G2084), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT45), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1058), .B1(new_n1070), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n1055), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1966), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(G8), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT51), .ZN(new_n1128));
  NOR2_X1   g703(.A1(G168), .A2(new_n1088), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT51), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1071), .A2(new_n761), .A3(new_n1077), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1068), .B2(G1966), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1131), .B1(new_n1137), .B2(G8), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1133), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT118), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1133), .B(new_n1141), .C1(new_n1135), .C2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1111), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1057), .A2(new_n833), .A3(new_n1125), .A4(new_n1119), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(G1961), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1078), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1068), .B2(new_n833), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1124), .A2(new_n1152), .A3(new_n833), .A4(new_n1125), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT53), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1151), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT120), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1146), .A2(KEYINPUT119), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(KEYINPUT53), .A3(new_n1154), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n1151), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1149), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT122), .B1(new_n1162), .B2(G301), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1149), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1159), .A2(new_n1160), .A3(new_n1151), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1160), .B1(new_n1159), .B2(new_n1151), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(G171), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1163), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1145), .A2(new_n1170), .A3(KEYINPUT123), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1140), .A2(KEYINPUT62), .A3(new_n1142), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT123), .B1(new_n1145), .B2(new_n1170), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1092), .B(KEYINPUT112), .Z(new_n1176));
  NOR2_X1   g751(.A1(G288), .A2(G1976), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1176), .B1(new_n1105), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1178), .A2(new_n1090), .B1(new_n1179), .B2(new_n1086), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT113), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT63), .ZN(new_n1182));
  OAI21_X1  g757(.A(G168), .B1(new_n1181), .B2(KEYINPUT63), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n1127), .A2(new_n1183), .ZN(new_n1184));
  OR3_X1    g759(.A1(new_n1111), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1182), .B1(new_n1111), .B2(new_n1184), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1180), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1147), .A2(KEYINPUT53), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1164), .A2(new_n1151), .A3(new_n1188), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1189), .A2(G171), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1163), .A2(new_n1169), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT54), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(KEYINPUT56), .B(G2072), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1068), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(G1956), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1078), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  OR2_X1    g773(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1199));
  NAND2_X1  g774(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1087), .A2(new_n850), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(G1348), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1202), .B1(new_n623), .B2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1195), .A2(new_n1197), .A3(new_n1200), .A4(new_n1199), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1078), .A2(new_n827), .ZN(new_n1210));
  AOI21_X1  g785(.A(KEYINPUT60), .B1(new_n1210), .B2(new_n1203), .ZN(new_n1211));
  OAI21_X1  g786(.A(KEYINPUT116), .B1(new_n1211), .B2(new_n623), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT116), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1213), .B(new_n631), .C1(new_n1206), .C2(KEYINPUT60), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1206), .A2(KEYINPUT60), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1212), .A2(new_n1216), .A3(new_n1214), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT59), .ZN(new_n1221));
  INV_X1    g796(.A(G1996), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1068), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT114), .ZN(new_n1224));
  INV_X1    g799(.A(new_n1087), .ZN(new_n1225));
  XOR2_X1   g800(.A(KEYINPUT58), .B(G1341), .Z(new_n1226));
  AOI22_X1  g801(.A1(new_n1223), .A2(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1068), .A2(KEYINPUT114), .A3(new_n1222), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n560), .A2(KEYINPUT115), .ZN(new_n1230));
  INV_X1    g805(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1221), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  AOI211_X1 g807(.A(KEYINPUT59), .B(new_n1230), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT61), .ZN(new_n1234));
  AND3_X1   g809(.A1(new_n1202), .A2(new_n1234), .A3(new_n1208), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1234), .B1(new_n1202), .B2(new_n1208), .ZN(new_n1236));
  OAI22_X1  g811(.A1(new_n1232), .A2(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1209), .B1(new_n1220), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1192), .B1(new_n1189), .B2(G171), .ZN(new_n1239));
  OAI21_X1  g814(.A(new_n1239), .B1(new_n1167), .B2(G171), .ZN(new_n1240));
  NOR2_X1   g815(.A1(new_n1143), .A2(new_n1111), .ZN(new_n1241));
  NAND3_X1  g816(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1187), .B1(new_n1193), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1066), .B1(new_n1175), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1059), .A2(new_n1222), .ZN(new_n1245));
  XNOR2_X1  g820(.A(new_n1245), .B(KEYINPUT46), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1061), .A2(new_n779), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1247), .A2(new_n1059), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g824(.A(new_n1249), .B(KEYINPUT47), .ZN(new_n1250));
  OR2_X1    g825(.A1(new_n1250), .A2(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1250), .A2(KEYINPUT124), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n1064), .A2(new_n1059), .ZN(new_n1253));
  NOR4_X1   g828(.A1(new_n1057), .A2(G290), .A3(G1986), .A4(new_n1058), .ZN(new_n1254));
  XOR2_X1   g829(.A(new_n1254), .B(KEYINPUT48), .Z(new_n1255));
  NAND2_X1  g830(.A1(new_n1062), .A2(new_n1061), .ZN(new_n1256));
  OAI22_X1  g831(.A1(new_n1256), .A2(new_n1063), .B1(G2067), .B2(new_n848), .ZN(new_n1257));
  AOI22_X1  g832(.A1(new_n1253), .A2(new_n1255), .B1(new_n1059), .B2(new_n1257), .ZN(new_n1258));
  AND3_X1   g833(.A1(new_n1251), .A2(new_n1252), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1244), .A2(new_n1259), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g835(.A(KEYINPUT125), .ZN(new_n1262));
  AOI21_X1  g836(.A(new_n462), .B1(new_n709), .B2(new_n717), .ZN(new_n1263));
  NAND2_X1  g837(.A1(new_n684), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g838(.A(new_n1262), .B1(G229), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g839(.A(new_n744), .ZN(new_n1266));
  NOR3_X1   g840(.A1(new_n741), .A2(new_n742), .A3(new_n719), .ZN(new_n1267));
  AOI21_X1  g841(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(new_n1268));
  OAI21_X1  g842(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g843(.A1(new_n743), .A2(new_n744), .A3(new_n752), .ZN(new_n1270));
  NAND2_X1  g844(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g845(.A1(new_n1271), .A2(KEYINPUT125), .A3(new_n684), .A4(new_n1263), .ZN(new_n1272));
  NAND2_X1  g846(.A1(new_n1265), .A2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g847(.A(new_n1273), .B1(new_n964), .B2(new_n966), .ZN(new_n1274));
  INV_X1    g848(.A(new_n1274), .ZN(new_n1275));
  AOI21_X1  g849(.A(new_n1041), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1276));
  NOR3_X1   g850(.A1(new_n1032), .A2(new_n1040), .A3(KEYINPUT43), .ZN(new_n1277));
  OAI21_X1  g851(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g852(.A1(new_n1278), .A2(KEYINPUT126), .ZN(new_n1279));
  INV_X1    g853(.A(KEYINPUT126), .ZN(new_n1280));
  NAND3_X1  g854(.A1(new_n1052), .A2(new_n1280), .A3(new_n1275), .ZN(new_n1281));
  NAND3_X1  g855(.A1(new_n1279), .A2(KEYINPUT127), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g856(.A(KEYINPUT127), .ZN(new_n1283));
  AOI21_X1  g857(.A(new_n1280), .B1(new_n1052), .B2(new_n1275), .ZN(new_n1284));
  AOI211_X1 g858(.A(KEYINPUT126), .B(new_n1274), .C1(new_n1047), .C2(new_n1051), .ZN(new_n1285));
  OAI21_X1  g859(.A(new_n1283), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g860(.A1(new_n1282), .A2(new_n1286), .ZN(G308));
  NAND2_X1  g861(.A1(new_n1279), .A2(new_n1281), .ZN(G225));
endmodule


