//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n458), .B1(new_n448), .B2(new_n455), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  XOR2_X1   g038(.A(KEYINPUT67), .B(G2105), .Z(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n466), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n465), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n471), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n462), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n462), .A2(new_n466), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n480), .A2(G124), .B1(new_n482), .B2(G136), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n464), .C2(G112), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NOR2_X1   g061(.A1(new_n472), .A2(new_n473), .ZN(new_n487));
  NAND2_X1  g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n466), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n474), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n464), .A2(new_n494), .A3(G138), .A4(new_n462), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n499), .A2(KEYINPUT68), .A3(G651), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT68), .B1(new_n499), .B2(G651), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G88), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n507), .A2(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  XOR2_X1   g087(.A(new_n512), .B(KEYINPUT69), .Z(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n515), .B1(new_n497), .B2(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n499), .A2(KEYINPUT68), .A3(G651), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(new_n517), .B1(KEYINPUT6), .B2(new_n497), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(G50), .A3(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n510), .A2(new_n514), .A3(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  AND3_X1   g096(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT71), .Z(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(G543), .B1(new_n518), .B2(KEYINPUT70), .ZN(new_n528));
  OAI211_X1 g103(.A(KEYINPUT70), .B(new_n498), .C1(new_n500), .C2(new_n501), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n509), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n527), .A2(new_n532), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(new_n531), .A2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n508), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n509), .A2(G90), .B1(new_n539), .B2(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  XNOR2_X1  g117(.A(KEYINPUT72), .B(G43), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n531), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n508), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n509), .A2(G81), .B1(new_n547), .B2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n502), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n557), .A2(G53), .A3(G543), .A4(new_n529), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n504), .B1(new_n502), .B2(new_n556), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n560), .A2(new_n561), .A3(G53), .A4(new_n529), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  XOR2_X1   g139(.A(KEYINPUT73), .B(G65), .Z(new_n565));
  AND2_X1   g140(.A1(new_n565), .A2(new_n507), .ZN(new_n566));
  AND2_X1   g141(.A1(G78), .A2(G543), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n564), .B(G651), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n565), .A2(new_n507), .B1(G78), .B2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT74), .B1(new_n569), .B2(new_n497), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n568), .A2(new_n570), .B1(G91), .B2(new_n509), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n563), .A2(new_n571), .ZN(G299));
  OR2_X1    g147(.A1(new_n507), .A2(G74), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n509), .A2(G87), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n560), .A2(G49), .A3(new_n529), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  AND2_X1   g151(.A1(G48), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n505), .B2(new_n506), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n518), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n505), .B2(new_n506), .ZN(new_n582));
  AND2_X1   g157(.A1(G73), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n531), .A2(G47), .ZN(new_n586));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n508), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n509), .A2(G85), .B1(new_n589), .B2(G651), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G290));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(G301), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n509), .A2(G92), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT75), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G651), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n596), .A2(KEYINPUT75), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G54), .ZN(new_n601));
  NOR3_X1   g176(.A1(new_n528), .A2(new_n530), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT76), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n497), .B1(new_n596), .B2(KEYINPUT75), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(KEYINPUT75), .B2(new_n596), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT76), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n560), .A2(new_n529), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n601), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n595), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n593), .B1(new_n611), .B2(new_n592), .ZN(G321));
  XNOR2_X1  g187(.A(G321), .B(KEYINPUT78), .ZN(G284));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n462), .A2(new_n467), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n480), .A2(G123), .ZN(new_n630));
  OAI221_X1 g205(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n482), .A2(G135), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2096), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n628), .A2(new_n629), .A3(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  OR2_X1    g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(new_n627), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(G2096), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT81), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT80), .B(KEYINPUT20), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n674), .A2(KEYINPUT81), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(KEYINPUT81), .ZN(new_n679));
  INV_X1    g254(.A(new_n676), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n671), .A2(new_n672), .ZN(new_n682));
  OR3_X1    g257(.A1(new_n670), .A2(new_n673), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n670), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n677), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G1981), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n685), .B1(new_n675), .B2(new_n676), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(KEYINPUT82), .A3(new_n681), .ZN(new_n692));
  AND3_X1   g267(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n690), .B1(new_n689), .B2(new_n692), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n667), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n689), .A2(new_n692), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G1981), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n697), .A2(G1986), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT83), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AND3_X1   g277(.A1(new_n695), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n695), .B2(new_n699), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n666), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n693), .A2(new_n694), .A3(new_n667), .ZN(new_n706));
  AOI21_X1  g281(.A(G1986), .B1(new_n697), .B2(new_n698), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n701), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n695), .A2(new_n699), .A3(new_n702), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n708), .A2(new_n665), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(new_n710), .ZN(G229));
  INV_X1    g286(.A(KEYINPUT95), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  INV_X1    g290(.A(G129), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n479), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n467), .A2(G105), .ZN(new_n718));
  INV_X1    g293(.A(G141), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n481), .B2(new_n719), .ZN(new_n720));
  OR3_X1    g295(.A1(new_n717), .A2(KEYINPUT89), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT89), .B1(new_n717), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n721), .A2(KEYINPUT90), .A3(new_n722), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n725), .A2(G29), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G32), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(G29), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT91), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n729), .B(new_n731), .Z(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  NAND2_X1  g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  INV_X1    g313(.A(G127), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n487), .B2(new_n739), .ZN(new_n740));
  AOI22_X1  g315(.A1(G139), .A2(new_n482), .B1(new_n740), .B2(new_n478), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n735), .B1(new_n743), .B2(new_n734), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(G2072), .ZN(new_n745));
  NOR2_X1   g320(.A1(G27), .A2(G29), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G164), .B2(G29), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n744), .A2(G2072), .B1(G2078), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n734), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n734), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT29), .B(G2090), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n745), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G5), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G171), .B2(new_n754), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1961), .Z(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n758), .B2(new_n759), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G160), .B2(new_n734), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G2084), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(G2084), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n633), .A2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT30), .B(G28), .ZN(new_n766));
  OR2_X1    g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT31), .A2(G11), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n766), .A2(new_n734), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND4_X1   g344(.A1(new_n763), .A2(new_n764), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n734), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n480), .A2(G128), .B1(new_n482), .B2(G140), .ZN(new_n774));
  OAI221_X1 g349(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n773), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT88), .B(G2067), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G2078), .ZN(new_n780));
  INV_X1    g355(.A(new_n747), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n753), .A2(new_n757), .A3(new_n770), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n733), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n754), .A2(G4), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n611), .B2(new_n754), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G1348), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT93), .B(KEYINPUT23), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n754), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G299), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1956), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n754), .A2(G21), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G286), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1966), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G1341), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n550), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G16), .B2(G19), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n797), .B2(new_n799), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n794), .A2(new_n795), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT92), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT92), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n784), .A2(new_n787), .A3(new_n792), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n786), .A2(G1348), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n713), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n783), .ZN(new_n809));
  AND4_X1   g384(.A1(new_n792), .A2(new_n809), .A3(new_n805), .A4(new_n732), .ZN(new_n810));
  INV_X1    g385(.A(new_n807), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n810), .A2(KEYINPUT94), .A3(new_n811), .A4(new_n787), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n754), .A2(G6), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n580), .A2(new_n584), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n754), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT32), .B(G1981), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G1971), .ZN(new_n819));
  NAND2_X1  g394(.A1(G166), .A2(G16), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G16), .B2(G22), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n819), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n754), .A2(G23), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n574), .A2(new_n575), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(new_n754), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT33), .B(G1976), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT86), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n829), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n822), .A2(new_n823), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT34), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n754), .A2(G24), .ZN(new_n834));
  INV_X1    g409(.A(G290), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n754), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT85), .B(G1986), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n734), .A2(G25), .ZN(new_n839));
  OAI221_X1 g414(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT84), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n480), .A2(G119), .B1(new_n482), .B2(G131), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n839), .B1(new_n843), .B2(G29), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G1991), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n838), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n833), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT36), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n832), .A2(KEYINPUT34), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n848), .B2(new_n850), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n712), .B1(new_n813), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g430(.A(KEYINPUT95), .B(new_n853), .C1(new_n808), .C2(new_n812), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(G311));
  NAND2_X1  g432(.A1(new_n813), .A2(new_n854), .ZN(G150));
  NAND2_X1  g433(.A1(new_n611), .A2(G559), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n549), .A2(KEYINPUT99), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n544), .A2(new_n861), .A3(new_n548), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(new_n497), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(KEYINPUT97), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(KEYINPUT97), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n866), .A2(new_n867), .B1(G93), .B2(new_n509), .ZN(new_n868));
  XNOR2_X1  g443(.A(KEYINPUT98), .B(G55), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n607), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n860), .A2(new_n862), .B1(new_n868), .B2(new_n870), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n859), .B(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n878));
  AOI21_X1  g453(.A(G860), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n871), .A2(G860), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT37), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(G145));
  INV_X1    g458(.A(new_n625), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n843), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n841), .A2(new_n625), .A3(new_n842), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n482), .A2(G142), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT101), .Z(new_n889));
  NOR2_X1   g464(.A1(new_n464), .A2(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n891));
  INV_X1    g466(.A(G130), .ZN(new_n892));
  OAI22_X1  g467(.A1(new_n890), .A2(new_n891), .B1(new_n892), .B2(new_n479), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n887), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n889), .A2(new_n893), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n885), .A2(new_n896), .A3(new_n886), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n895), .B1(new_n894), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n493), .A2(new_n495), .ZN(new_n901));
  INV_X1    g476(.A(new_n491), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n742), .B1(new_n725), .B2(new_n726), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n723), .A2(new_n742), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n726), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT90), .B1(new_n721), .B2(new_n722), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n743), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(G164), .A3(new_n905), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n776), .B(KEYINPUT100), .Z(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n907), .B2(new_n911), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n900), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n633), .B(G160), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n485), .ZN(new_n919));
  INV_X1    g494(.A(new_n916), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(new_n899), .A3(new_n914), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n919), .B1(new_n917), .B2(new_n921), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n926), .B(KEYINPUT40), .Z(G395));
  XOR2_X1   g502(.A(new_n620), .B(new_n874), .Z(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n603), .A2(new_n608), .ZN(new_n930));
  INV_X1    g505(.A(new_n595), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n615), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n609), .A2(G299), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n929), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT41), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n933), .A2(new_n939), .A3(new_n934), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n928), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n934), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n609), .A2(G299), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT103), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n936), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n928), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(G288), .B(G305), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(G303), .B(KEYINPUT104), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(G290), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(G290), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n953), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n951), .A3(new_n948), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(KEYINPUT105), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n957), .B(new_n958), .Z(new_n959));
  AND3_X1   g534(.A1(new_n942), .A2(new_n947), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n942), .B2(new_n947), .ZN(new_n961));
  OAI21_X1  g536(.A(G868), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n868), .A2(new_n870), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n962), .B1(G868), .B2(new_n963), .ZN(G295));
  OAI21_X1  g539(.A(new_n962), .B1(G868), .B2(new_n963), .ZN(G331));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n954), .A2(new_n956), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n860), .A3(new_n862), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n863), .A2(new_n871), .ZN(new_n969));
  NAND2_X1  g544(.A1(G286), .A2(G301), .ZN(new_n970));
  NAND2_X1  g545(.A1(G168), .A2(G171), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n970), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n872), .B2(new_n873), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n938), .B2(new_n940), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n974), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n946), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n967), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n954), .A2(new_n956), .A3(KEYINPUT107), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT107), .B1(new_n954), .B2(new_n956), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n977), .B(KEYINPUT41), .C1(new_n943), .C2(new_n944), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n975), .A2(new_n939), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n982), .B(new_n983), .C1(new_n984), .C2(new_n946), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n979), .A2(new_n985), .A3(new_n923), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n966), .B1(new_n986), .B2(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n941), .A2(new_n977), .ZN(new_n988));
  INV_X1    g563(.A(new_n978), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n989), .A3(new_n982), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(new_n979), .A3(new_n923), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n987), .B1(KEYINPUT43), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n979), .A2(new_n985), .A3(new_n994), .A4(new_n923), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT108), .B1(new_n996), .B2(new_n966), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n998), .B(KEYINPUT44), .C1(new_n993), .C2(new_n995), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n992), .B1(new_n997), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(G164), .B2(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G40), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n465), .A2(new_n1004), .A3(new_n476), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OR3_X1    g581(.A1(new_n1006), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT46), .B1(new_n1006), .B2(G1996), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n776), .A2(G2067), .ZN(new_n1009));
  INV_X1    g584(.A(G2067), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n774), .A2(new_n1010), .A3(new_n775), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(new_n723), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1006), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1007), .A2(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1015), .B(KEYINPUT47), .Z(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n667), .A3(new_n835), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT48), .ZN(new_n1018));
  INV_X1    g593(.A(G1996), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n908), .B2(new_n909), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n843), .B(new_n845), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1012), .B1(G1996), .B2(new_n723), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1018), .B1(new_n1024), .B2(new_n1006), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n841), .A2(new_n845), .A3(new_n842), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1011), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1014), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1016), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n563), .A2(new_n1031), .A3(new_n571), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n563), .B2(new_n571), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n903), .A2(KEYINPUT45), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(KEYINPUT109), .A3(new_n1002), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1384), .B1(new_n901), .B2(new_n902), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT56), .B(G2072), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1005), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1956), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1005), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1034), .B1(new_n1043), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT61), .B1(new_n1050), .B2(KEYINPUT120), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G160), .A2(G40), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1042), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n1053), .B(new_n1054), .C1(new_n1037), .C2(new_n1040), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1049), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1043), .A2(new_n1034), .A3(new_n1049), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1051), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(KEYINPUT61), .A3(new_n1059), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1053), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1064), .A2(new_n1019), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1038), .A2(new_n1005), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1067), .B(new_n797), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1063), .B(new_n550), .C1(new_n1065), .C2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1064), .B2(new_n1019), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT59), .B1(new_n1071), .B2(new_n549), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1348), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1066), .A2(new_n1010), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1077), .A2(KEYINPUT60), .A3(new_n932), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n609), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n932), .A2(new_n1076), .A3(new_n1075), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1081), .B2(KEYINPUT60), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1061), .A2(new_n1062), .A3(new_n1073), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n932), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1059), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n1057), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1085), .B2(new_n1057), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1048), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1961), .B1(new_n1092), .B2(new_n1046), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1002), .A2(KEYINPUT117), .A3(new_n1005), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1036), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1096), .A2(G2078), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n1036), .A3(new_n1095), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT121), .B1(new_n1104), .B2(G2078), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1093), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g681(.A(G2078), .B(new_n1053), .C1(new_n1037), .C2(new_n1040), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT122), .B1(new_n1107), .B2(KEYINPUT53), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1064), .A2(new_n780), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n1094), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(G301), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(new_n476), .B(KEYINPUT123), .Z(new_n1114));
  NAND3_X1  g689(.A1(new_n780), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1114), .A2(new_n465), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1093), .B1(new_n1041), .B2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1112), .A2(G301), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1091), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1106), .A2(new_n1112), .A3(G301), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1120), .B(KEYINPUT54), .C1(new_n1121), .C2(G301), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1092), .A2(new_n1046), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT110), .B(G2090), .Z(new_n1124));
  OAI22_X1  g699(.A1(new_n1064), .A2(G1971), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(G303), .A2(G8), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT55), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(G8), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1038), .B2(new_n1005), .ZN(new_n1131));
  INV_X1    g706(.A(G1976), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(G288), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT52), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n825), .A2(G1976), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1135), .A2(new_n1131), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(G288), .B2(new_n1132), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1134), .A2(KEYINPUT111), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1135), .A2(new_n1137), .A3(KEYINPUT111), .A4(new_n1131), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT112), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n815), .A2(new_n1140), .A3(new_n690), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT112), .B1(G305), .B2(G1981), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT113), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n580), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n518), .B(KEYINPUT113), .C1(new_n577), .C2(new_n579), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n584), .A3(new_n1145), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1141), .A2(new_n1142), .B1(new_n1146), .B2(G1981), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1131), .B1(new_n1147), .B2(KEYINPUT49), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1146), .A2(G1981), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1149), .A2(KEYINPUT49), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1139), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1138), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1128), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1125), .A2(G8), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1129), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1123), .A2(G2084), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1104), .A2(new_n795), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(G168), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(G8), .ZN(new_n1160));
  AOI21_X1  g735(.A(G168), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT51), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT51), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1163), .A3(G8), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1156), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1090), .A2(new_n1119), .A3(new_n1122), .A4(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1132), .B(new_n825), .C1(new_n1148), .C2(new_n1151), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT115), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n1149), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1167), .B2(new_n1149), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT114), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1131), .B(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1138), .A2(new_n1152), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1155), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT116), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1174), .A2(new_n1155), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1170), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1167), .A2(new_n1168), .A3(new_n1149), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1172), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT116), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1177), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n1184));
  AOI211_X1 g759(.A(new_n1130), .B(G286), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1156), .B2(new_n1186), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1188), .A2(KEYINPUT63), .A3(new_n1129), .A4(new_n1185), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1176), .A2(new_n1183), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1166), .A2(new_n1190), .A3(KEYINPUT124), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT124), .B1(new_n1166), .B2(new_n1190), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1162), .A2(new_n1193), .A3(new_n1164), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1194), .A2(new_n1113), .A3(new_n1129), .A4(new_n1188), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1196), .B1(new_n1197), .B2(KEYINPUT62), .ZN(new_n1198));
  AOI211_X1 g773(.A(KEYINPUT125), .B(new_n1193), .C1(new_n1162), .C2(new_n1164), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1195), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1191), .A2(new_n1192), .A3(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(G290), .B(new_n667), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1006), .B1(new_n1024), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1030), .B1(new_n1201), .B2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g779(.A1(new_n460), .A2(G227), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1206), .A2(new_n651), .ZN(new_n1207));
  XNOR2_X1  g781(.A(new_n1207), .B(KEYINPUT126), .ZN(new_n1208));
  NAND3_X1  g782(.A1(new_n705), .A2(new_n710), .A3(new_n1208), .ZN(new_n1209));
  NOR2_X1   g783(.A1(new_n926), .A2(new_n1209), .ZN(new_n1210));
  AND3_X1   g784(.A1(new_n996), .A2(new_n1210), .A3(KEYINPUT127), .ZN(new_n1211));
  AOI21_X1  g785(.A(KEYINPUT127), .B1(new_n996), .B2(new_n1210), .ZN(new_n1212));
  NOR2_X1   g786(.A1(new_n1211), .A2(new_n1212), .ZN(G308));
  NAND2_X1  g787(.A1(new_n996), .A2(new_n1210), .ZN(G225));
endmodule


