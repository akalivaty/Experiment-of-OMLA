//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1294, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1349, new_n1350, new_n1351;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(new_n204), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT64), .Z(new_n213));
  AOI21_X1  g0013(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT65), .B(G238), .Z(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n214), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT66), .Z(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n210), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT70), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n244), .A2(KEYINPUT70), .A3(new_n210), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G13), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT71), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(new_n204), .B2(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n203), .A2(KEYINPUT71), .A3(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n254), .A2(G50), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G150), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n261), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G58), .A2(G68), .ZN(new_n267));
  INV_X1    g0067(.A(G50), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n204), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n249), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n259), .B(new_n270), .C1(G50), .C2(new_n252), .ZN(new_n271));
  XOR2_X1   g0071(.A(new_n271), .B(KEYINPUT9), .Z(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT68), .B(G45), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n210), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n279), .A2(new_n280), .B1(new_n282), .B2(new_n203), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n278), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G222), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  INV_X1    g0093(.A(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G1698), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT69), .B(G223), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n292), .B1(new_n293), .B2(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n279), .A2(new_n280), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n286), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G190), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n300), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n272), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n301), .B(KEYINPUT75), .C1(new_n302), .C2(new_n300), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n306), .B(new_n305), .C1(new_n272), .C2(new_n303), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G244), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n278), .B1(new_n284), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n291), .A2(G232), .ZN(new_n313));
  INV_X1    g0113(.A(G107), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n313), .B1(new_n314), .B2(new_n294), .C1(new_n215), .C2(new_n295), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n315), .B2(new_n299), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n316), .A2(G169), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n262), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT73), .B1(new_n322), .B2(new_n265), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n322), .A2(new_n265), .A3(KEYINPUT73), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n245), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n253), .A2(new_n245), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n293), .B1(new_n256), .B2(new_n257), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n327), .A2(new_n328), .B1(new_n293), .B2(new_n253), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n317), .A2(new_n319), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n316), .B2(G190), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n302), .B2(new_n316), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT74), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT72), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n300), .A2(new_n318), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n271), .B1(new_n300), .B2(G169), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n300), .A2(G169), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n341), .A2(KEYINPUT72), .A3(new_n271), .A4(new_n337), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n334), .B1(new_n331), .B2(new_n333), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n275), .A2(KEYINPUT76), .A3(new_n277), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n283), .A2(G238), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT76), .B1(new_n275), .B2(new_n277), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n287), .A2(new_n289), .A3(G232), .A4(G1698), .ZN(new_n353));
  INV_X1    g0153(.A(G1698), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n287), .A2(new_n289), .A3(G226), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G97), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n353), .B(new_n355), .C1(new_n263), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n299), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n347), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n278), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n348), .A3(new_n349), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n357), .A2(new_n299), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT13), .ZN(new_n364));
  OAI21_X1  g0164(.A(G169), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT14), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n348), .A2(new_n349), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n367), .A2(new_n347), .A3(new_n358), .A4(new_n361), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT77), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT77), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n352), .A2(new_n370), .A3(new_n347), .A4(new_n358), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT13), .B1(new_n362), .B2(new_n363), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n369), .A2(G179), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(G169), .C1(new_n359), .C2(new_n364), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n366), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n265), .B2(new_n293), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n249), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT11), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT78), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n249), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n253), .A2(new_n216), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT12), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n327), .A2(G68), .A3(new_n258), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n381), .B1(new_n380), .B2(new_n383), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n384), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n376), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n369), .A2(G190), .A3(new_n371), .A4(new_n372), .ZN(new_n393));
  OAI21_X1  g0193(.A(G200), .B1(new_n359), .B2(new_n364), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(new_n390), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n310), .A2(new_n346), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n281), .A2(G1), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT84), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(KEYINPUT5), .C2(new_n274), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n203), .B(G45), .C1(new_n274), .C2(KEYINPUT5), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT84), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT5), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(G41), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(new_n276), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n400), .A2(new_n402), .A3(new_n298), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G270), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n298), .B1(new_n401), .B2(new_n404), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(G257), .A2(G1698), .ZN(new_n410));
  INV_X1    g0210(.A(G264), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n411), .B2(G1698), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n288), .A2(KEYINPUT79), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT79), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT3), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n416), .A3(G33), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT80), .B1(new_n288), .B2(G33), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT80), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n414), .A2(new_n416), .A3(new_n421), .A4(G33), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n413), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G303), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n294), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT86), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n418), .B1(new_n427), .B2(G33), .ZN(new_n428));
  AND4_X1   g0228(.A1(new_n421), .A2(new_n414), .A3(new_n416), .A4(G33), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n412), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n425), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT86), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n426), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n409), .B1(new_n434), .B2(new_n299), .ZN(new_n435));
  INV_X1    g0235(.A(G169), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G283), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n204), .C1(G33), .C2(new_n356), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n204), .A2(G116), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n440), .A3(new_n245), .ZN(new_n441));
  XOR2_X1   g0241(.A(new_n441), .B(KEYINPUT20), .Z(new_n442));
  INV_X1    g0242(.A(G116), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n203), .B2(G33), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n327), .A2(new_n444), .B1(new_n439), .B2(new_n251), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n436), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT21), .B1(new_n435), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT21), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n298), .B1(new_n426), .B2(new_n433), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n446), .B(new_n449), .C1(new_n450), .C2(new_n409), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n434), .A2(new_n299), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n442), .A2(new_n445), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n409), .A2(new_n318), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n454), .ZN(new_n457));
  OAI21_X1  g0257(.A(G200), .B1(new_n450), .B2(new_n409), .ZN(new_n458));
  INV_X1    g0258(.A(new_n409), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G190), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n457), .B(new_n458), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n452), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G238), .A2(G1698), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n311), .B2(G1698), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n428), .B2(new_n429), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n263), .A2(new_n443), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n298), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT85), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n398), .A2(G250), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n398), .A2(new_n276), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n298), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n465), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n420), .B2(new_n422), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n299), .B1(new_n477), .B2(new_n467), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT85), .B1(new_n478), .B2(new_n473), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n436), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(G20), .B1(new_n420), .B2(new_n422), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G68), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT19), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n264), .A2(new_n483), .A3(G97), .ZN(new_n484));
  AOI21_X1  g0284(.A(G20), .B1(G33), .B2(G97), .ZN(new_n485));
  INV_X1    g0285(.A(G87), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G97), .A2(G107), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n484), .B1(new_n488), .B2(new_n483), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n245), .ZN(new_n491));
  INV_X1    g0291(.A(new_n322), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n252), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n203), .A2(G33), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n247), .A2(new_n252), .A3(new_n495), .A4(new_n248), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n491), .B(new_n494), .C1(new_n496), .C2(new_n322), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n470), .B1(new_n469), .B2(new_n474), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n478), .A2(KEYINPUT85), .A3(new_n473), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n318), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n480), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(G200), .B1(new_n475), .B2(new_n479), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n498), .A2(G190), .A3(new_n499), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n496), .A2(new_n486), .ZN(new_n504));
  AOI211_X1 g0304(.A(new_n493), .B(new_n504), .C1(new_n490), .C2(new_n245), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n496), .A2(G97), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n252), .A2(new_n356), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT83), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT83), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT6), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n356), .A2(new_n314), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n515), .B2(new_n487), .ZN(new_n516));
  NAND2_X1  g0316(.A1(KEYINPUT6), .A2(G97), .ZN(new_n517));
  OR3_X1    g0317(.A1(new_n517), .A2(KEYINPUT82), .A3(G107), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT82), .B1(new_n517), .B2(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G20), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n260), .A2(G77), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n289), .B1(new_n427), .B2(G33), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT7), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(G20), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n290), .A2(new_n204), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n523), .A2(new_n525), .B1(new_n526), .B2(new_n524), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n521), .B(new_n522), .C1(new_n527), .C2(new_n314), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n245), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n513), .A2(new_n529), .ZN(new_n530));
  AND4_X1   g0330(.A1(new_n400), .A2(new_n402), .A3(new_n298), .A4(new_n405), .ZN(new_n531));
  INV_X1    g0331(.A(new_n408), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(G257), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n311), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(new_n354), .A3(new_n287), .A4(new_n289), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n287), .A2(new_n289), .A3(G250), .A4(G1698), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n437), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n311), .A2(G1698), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n428), .B2(new_n429), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n538), .B1(new_n540), .B2(new_n534), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n533), .B1(new_n541), .B2(new_n298), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n436), .ZN(new_n543));
  INV_X1    g0343(.A(new_n539), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n420), .B2(new_n422), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(KEYINPUT4), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n299), .B1(new_n546), .B2(new_n538), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(new_n318), .A3(new_n533), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n530), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n542), .A2(G200), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n510), .A2(new_n512), .B1(new_n528), .B2(new_n245), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(G190), .A3(new_n533), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AND4_X1   g0353(.A1(new_n501), .A2(new_n506), .A3(new_n549), .A4(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(G250), .B(new_n354), .C1(new_n428), .C2(new_n429), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT90), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n420), .A2(new_n422), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT90), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(G250), .A4(new_n354), .ZN(new_n559));
  AND2_X1   g0359(.A1(G257), .A2(G1698), .ZN(new_n560));
  XOR2_X1   g0360(.A(KEYINPUT91), .B(G294), .Z(new_n561));
  AOI22_X1  g0361(.A1(new_n557), .A2(new_n560), .B1(G33), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n556), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n299), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n532), .A2(G264), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n564), .A2(new_n318), .A3(new_n406), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n565), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n563), .B2(new_n299), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n406), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n436), .ZN(new_n570));
  INV_X1    g0370(.A(new_n245), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT22), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n486), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n481), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT24), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n204), .A2(G87), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n572), .B1(new_n290), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT23), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n204), .B2(G107), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n314), .A2(KEYINPUT23), .A3(G20), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n579), .A2(new_n580), .B1(new_n467), .B2(new_n204), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n574), .A2(new_n575), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT87), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n582), .B1(new_n481), .B2(new_n573), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(KEYINPUT87), .A3(new_n575), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n574), .A2(new_n583), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT88), .B1(new_n590), .B2(KEYINPUT24), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT88), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n587), .A2(new_n592), .A3(new_n575), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n571), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n252), .A2(G107), .ZN(new_n596));
  XNOR2_X1  g0396(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n596), .B(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n314), .B2(new_n496), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n566), .B(new_n570), .C1(new_n595), .C2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n564), .A2(new_n461), .A3(new_n406), .A4(new_n565), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n531), .B(new_n567), .C1(new_n563), .C2(new_n299), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(G200), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n590), .A2(KEYINPUT88), .A3(KEYINPUT24), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n592), .B1(new_n587), .B2(new_n575), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n586), .A3(new_n605), .A4(new_n588), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n599), .B1(new_n606), .B2(new_n245), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n463), .A2(new_n554), .A3(new_n600), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n320), .A2(new_n258), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n254), .A2(new_n611), .B1(new_n253), .B2(new_n262), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g0413(.A(G58), .B(G68), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n614), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n527), .B2(new_n216), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT16), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n571), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n420), .A2(new_n204), .A3(new_n422), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n619), .A2(KEYINPUT7), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n420), .A2(new_n524), .A3(new_n204), .A4(new_n422), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G68), .ZN(new_n622));
  OAI211_X1 g0422(.A(KEYINPUT16), .B(new_n615), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n613), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n285), .A2(G1698), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(G223), .B2(G1698), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n420), .B2(new_n422), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n263), .A2(new_n486), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n299), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n283), .A2(G232), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n278), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n461), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n626), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n428), .B2(new_n429), .ZN(new_n635));
  INV_X1    g0435(.A(new_n628), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n631), .B1(new_n637), .B2(new_n299), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n633), .B1(new_n638), .B2(G200), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n624), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT17), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n624), .A2(KEYINPUT17), .A3(new_n639), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT18), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n618), .A2(new_n623), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n612), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n436), .B1(new_n629), .B2(new_n632), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n638), .A2(G179), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n645), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n629), .A2(G179), .A3(new_n632), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n648), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n624), .A2(new_n654), .A3(KEYINPUT18), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT81), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n647), .A2(new_n645), .A3(new_n651), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT81), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT18), .B1(new_n624), .B2(new_n654), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n644), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n397), .A2(new_n609), .A3(new_n661), .ZN(G372));
  NOR2_X1   g0462(.A1(new_n397), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n478), .A2(new_n473), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n436), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n497), .A2(new_n500), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n566), .B1(new_n602), .B2(G169), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n607), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n452), .A2(new_n456), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n549), .A2(new_n553), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n664), .A2(G200), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n503), .A2(new_n505), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n608), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n666), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n530), .A2(new_n543), .A3(new_n548), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n501), .A2(new_n676), .A3(new_n506), .A4(KEYINPUT26), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(KEYINPUT92), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(new_n666), .A3(new_n673), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT92), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n678), .B1(new_n683), .B2(new_n677), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n663), .B1(new_n675), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n652), .A2(new_n655), .ZN(new_n686));
  INV_X1    g0486(.A(new_n331), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n391), .A2(new_n376), .B1(new_n687), .B2(new_n395), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n642), .A2(new_n643), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n690), .A2(new_n310), .B1(new_n340), .B2(new_n342), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(G369));
  INV_X1    g0492(.A(new_n251), .ZN(new_n693));
  OR3_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .A3(G20), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT27), .B1(new_n693), .B2(G20), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n457), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n669), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n452), .A2(new_n456), .A3(new_n462), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n603), .A2(new_n607), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n668), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n607), .B2(new_n699), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n668), .A2(new_n698), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n698), .B1(new_n452), .B2(new_n456), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n668), .A2(new_n699), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n716), .ZN(G399));
  NAND2_X1  g0517(.A1(new_n207), .A2(new_n274), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT93), .Z(new_n719));
  NAND3_X1  g0519(.A1(new_n487), .A2(new_n486), .A3(new_n443), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n719), .A2(new_n203), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n213), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  INV_X1    g0523(.A(new_n666), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n673), .A2(new_n549), .A3(new_n553), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n607), .B2(new_n603), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n452), .B(new_n456), .C1(new_n667), .C2(new_n607), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n501), .A2(new_n676), .A3(new_n506), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n680), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n680), .B2(new_n679), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n698), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n501), .A2(new_n506), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(new_n682), .A3(KEYINPUT26), .A4(new_n676), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT92), .B1(new_n679), .B2(new_n680), .ZN(new_n736));
  INV_X1    g0536(.A(new_n677), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n698), .B1(new_n738), .B2(new_n728), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n733), .B1(KEYINPUT29), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n564), .A2(new_n565), .A3(new_n498), .A4(new_n499), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n453), .A2(new_n455), .A3(new_n547), .A4(new_n533), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n455), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n542), .A2(new_n450), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n475), .A2(new_n479), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n746), .A2(KEYINPUT30), .A3(new_n568), .A4(new_n747), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n542), .A2(new_n318), .A3(new_n664), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n569), .A2(new_n749), .A3(new_n460), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n744), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n698), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(new_n609), .C2(new_n698), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n740), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n723), .B1(new_n759), .B2(G1), .ZN(G364));
  NOR2_X1   g0560(.A1(new_n250), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n203), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n719), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n705), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G330), .B2(new_n703), .ZN(new_n766));
  NAND2_X1  g0566(.A1(G355), .A2(KEYINPUT94), .ZN(new_n767));
  OR2_X1    g0567(.A1(G355), .A2(KEYINPUT94), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n207), .A2(new_n294), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n557), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n207), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n213), .A2(new_n273), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n242), .B2(new_n281), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n769), .B1(G116), .B2(new_n207), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n210), .B1(G20), .B2(new_n436), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n764), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n204), .A2(G179), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT96), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(KEYINPUT96), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT97), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT32), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT32), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n204), .A2(new_n318), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n796), .A2(new_n461), .A3(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n785), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n797), .A2(G58), .B1(G77), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n796), .A2(new_n302), .A3(G190), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n800), .B1(new_n216), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n784), .A2(new_n461), .A3(G200), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G107), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n796), .A2(new_n461), .A3(new_n302), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n294), .B(new_n806), .C1(new_n808), .C2(new_n268), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n486), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n461), .A2(G179), .A3(G200), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n204), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n356), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n803), .A2(new_n809), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n793), .A2(new_n794), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n789), .B(KEYINPUT98), .Z(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G329), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n807), .A2(G326), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n797), .A2(G322), .B1(G311), .B2(new_n799), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n821), .A2(new_n804), .B1(new_n810), .B2(new_n424), .ZN(new_n822));
  XOR2_X1   g0622(.A(KEYINPUT33), .B(G317), .Z(new_n823));
  OAI21_X1  g0623(.A(new_n290), .B1(new_n802), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n813), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n822), .B(new_n824), .C1(new_n561), .C2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT99), .B1(new_n816), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n780), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n816), .A2(KEYINPUT99), .A3(new_n827), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n782), .B(new_n783), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n779), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n703), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n766), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G396));
  OAI22_X1  g0636(.A1(new_n802), .A2(new_n821), .B1(new_n798), .B2(new_n443), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G294), .B2(new_n797), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n290), .B1(new_n808), .B2(new_n424), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n805), .A2(G87), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n314), .B2(new_n810), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n839), .A2(new_n814), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n817), .ZN(new_n843));
  INV_X1    g0643(.A(G311), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n838), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n817), .A2(G132), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n801), .A2(G150), .B1(new_n807), .B2(G137), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n797), .A2(G143), .B1(G159), .B2(new_n799), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n850));
  INV_X1    g0650(.A(G58), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n557), .B1(new_n851), .B2(new_n813), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n849), .B2(KEYINPUT34), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n805), .A2(G68), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n268), .B2(new_n810), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT100), .Z(new_n856));
  NAND4_X1  g0656(.A1(new_n846), .A2(new_n850), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n829), .B1(new_n845), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n780), .A2(new_n777), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n783), .B(new_n858), .C1(new_n293), .C2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n330), .A2(new_n698), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n333), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n331), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n687), .A2(new_n699), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n861), .B1(new_n777), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n331), .A2(new_n333), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n869), .B(new_n699), .C1(new_n684), .C2(new_n675), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n739), .B2(new_n866), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n871), .A2(new_n757), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n764), .B1(new_n871), .B2(new_n757), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(G384));
  NAND4_X1  g0675(.A1(new_n707), .A2(new_n463), .A3(new_n554), .A4(new_n699), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n755), .A2(KEYINPUT105), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT105), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n751), .A2(new_n878), .A3(KEYINPUT31), .A4(new_n698), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n876), .A2(new_n754), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n390), .A2(new_n699), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n392), .A2(new_n395), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT102), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n395), .A2(new_n373), .A3(new_n375), .A4(new_n366), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n884), .B1(new_n885), .B2(new_n881), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n884), .A3(new_n881), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n887), .A2(new_n866), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n623), .A2(new_n249), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n619), .A2(KEYINPUT7), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(G68), .A3(new_n621), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT16), .B1(new_n895), .B2(new_n615), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n612), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n696), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n658), .B1(new_n657), .B2(new_n659), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n689), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n901), .B2(new_n660), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n647), .A2(new_n651), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n647), .A2(new_n898), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .A4(new_n640), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT103), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n646), .A2(new_n639), .A3(new_n612), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n646), .A2(new_n612), .B1(new_n649), .B2(new_n650), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(KEYINPUT103), .A3(new_n905), .A4(new_n904), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n897), .A2(new_n651), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n899), .A2(new_n913), .A3(new_n640), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n908), .A2(new_n912), .B1(KEYINPUT37), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n892), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n696), .B1(new_n646), .B2(new_n612), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n909), .A2(new_n910), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT103), .B1(new_n919), .B2(new_n905), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n906), .A2(new_n907), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n899), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n661), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n922), .A2(new_n924), .A3(KEYINPUT38), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT104), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n916), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n916), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n891), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n911), .A2(new_n904), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n908), .A2(new_n912), .B1(KEYINPUT37), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n904), .B1(new_n644), .B2(new_n686), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n892), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n925), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n880), .A2(new_n889), .A3(KEYINPUT40), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n929), .A2(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n663), .A2(new_n880), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  INV_X1    g0740(.A(G330), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n870), .A2(new_n865), .ZN(new_n943));
  INV_X1    g0743(.A(new_n888), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n883), .B2(new_n886), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n943), .B(new_n945), .C1(new_n927), .C2(new_n928), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n935), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n392), .A2(new_n698), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n916), .A2(new_n925), .A3(KEYINPUT39), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n696), .B1(new_n652), .B2(new_n655), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n946), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n733), .B(new_n663), .C1(KEYINPUT29), .C2(new_n739), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n691), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n953), .B(new_n955), .Z(new_n956));
  OAI22_X1  g0756(.A1(new_n942), .A2(new_n956), .B1(new_n203), .B2(new_n761), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n956), .B2(new_n942), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n959), .A2(G116), .A3(new_n211), .A4(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT36), .Z(new_n962));
  OAI211_X1 g0762(.A(new_n213), .B(G77), .C1(new_n851), .C2(new_n216), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n268), .A2(G68), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n203), .B(G13), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n958), .A2(new_n962), .A3(new_n965), .ZN(G367));
  OAI221_X1 g0766(.A(new_n781), .B1(new_n207), .B2(new_n322), .C1(new_n773), .C2(new_n235), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(new_n764), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n666), .A2(new_n505), .A3(new_n699), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n666), .B(new_n673), .C1(new_n505), .C2(new_n699), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n804), .A2(new_n293), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n294), .B1(new_n268), .B2(new_n798), .C1(new_n802), .C2(new_n790), .ZN(new_n973));
  INV_X1    g0773(.A(new_n810), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n972), .B(new_n973), .C1(G58), .C2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(KEYINPUT113), .B(G137), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n789), .B2(new_n976), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n797), .A2(G150), .B1(new_n807), .B2(G143), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n216), .B2(new_n813), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT112), .Z(new_n980));
  NOR2_X1   g0780(.A1(new_n810), .A2(new_n443), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n770), .B1(KEYINPUT46), .B2(new_n981), .C1(new_n789), .C2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n797), .ZN(new_n984));
  INV_X1    g0784(.A(new_n561), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n424), .A2(new_n984), .B1(new_n802), .B2(new_n985), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n808), .A2(new_n844), .B1(new_n798), .B2(new_n821), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n805), .A2(G97), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n314), .B2(new_n813), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n981), .A2(KEYINPUT46), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(KEYINPUT111), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(KEYINPUT111), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n977), .A2(new_n980), .B1(new_n983), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT114), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  OAI221_X1 g0797(.A(new_n968), .B1(new_n833), .B2(new_n971), .C1(new_n997), .C2(new_n829), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n530), .A2(new_n698), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n671), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n676), .A2(new_n698), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n999), .B1(new_n715), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n713), .A2(KEYINPUT45), .A3(new_n714), .A4(new_n1003), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT44), .B1(new_n715), .B2(new_n1004), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n715), .A2(KEYINPUT44), .A3(new_n1004), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1007), .B(new_n711), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1008), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1013), .A2(new_n1009), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT110), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n1015), .A3(new_n711), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n713), .B1(new_n710), .B2(new_n712), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1019), .B(new_n713), .C1(new_n710), .C2(new_n712), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(new_n758), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1014), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n711), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1017), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n759), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n719), .B(KEYINPUT41), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n763), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT108), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n668), .A2(new_n671), .A3(new_n1000), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n698), .B1(new_n1034), .B2(new_n549), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT42), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n707), .A2(new_n1003), .A3(new_n712), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT106), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(KEYINPUT42), .A3(new_n1039), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1035), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n971), .B(KEYINPUT43), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1033), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1035), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1040), .A2(new_n1041), .A3(new_n1036), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT42), .B1(new_n1043), .B2(new_n1039), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1046), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(KEYINPUT108), .A3(new_n1052), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT107), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1045), .A2(KEYINPUT107), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1054), .A2(new_n1060), .B1(new_n711), .B2(new_n1004), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n711), .A2(new_n1004), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1062), .A2(new_n1063), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n998), .B1(new_n1032), .B2(new_n1065), .ZN(G387));
  NAND3_X1  g0866(.A1(new_n1024), .A2(KEYINPUT118), .A3(new_n758), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n719), .C1(new_n758), .C2(new_n1024), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT118), .B1(new_n1024), .B2(new_n758), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OR3_X1    g0870(.A1(new_n1024), .A2(KEYINPUT115), .A3(new_n762), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT115), .B1(new_n1024), .B2(new_n762), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n708), .A2(new_n709), .A3(new_n779), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n801), .A2(new_n320), .B1(G68), .B2(new_n799), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT116), .Z(new_n1075));
  OAI221_X1 g0875(.A(new_n988), .B1(new_n808), .B2(new_n790), .C1(new_n268), .C2(new_n984), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n813), .A2(new_n322), .B1(new_n810), .B2(new_n293), .ZN(new_n1077));
  INV_X1    g0877(.A(G150), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n557), .B1(new_n789), .B2(new_n1078), .ZN(new_n1079));
  OR4_X1    g0879(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n789), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(G326), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n557), .B1(G116), .B2(new_n805), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n985), .A2(new_n810), .B1(new_n813), .B2(new_n821), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n801), .A2(G311), .B1(new_n807), .B2(G322), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n424), .B2(new_n798), .C1(new_n982), .C2(new_n984), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT49), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1082), .B(new_n1083), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1080), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1093), .A2(KEYINPUT117), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n829), .B1(new_n1093), .B2(KEYINPUT117), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n207), .A2(new_n294), .A3(new_n720), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n231), .A2(new_n273), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1097), .B1(new_n773), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(G45), .B(new_n720), .C1(G68), .C2(G77), .ZN(new_n1100));
  OR3_X1    g0900(.A1(new_n262), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT50), .B1(new_n262), .B2(G50), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(G107), .B2(new_n207), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n783), .B(new_n1096), .C1(new_n781), .C2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1071), .A2(new_n1072), .B1(new_n1073), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1070), .A2(new_n1107), .ZN(G393));
  OR3_X1    g0908(.A1(new_n1014), .A2(KEYINPUT119), .A3(new_n711), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT119), .B1(new_n1014), .B2(new_n711), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(new_n1110), .B1(new_n1016), .B2(new_n1012), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1029), .B(new_n719), .C1(new_n1111), .C2(new_n1025), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1004), .A2(new_n779), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n781), .B1(new_n356), .B2(new_n207), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n772), .B2(new_n239), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n797), .A2(G311), .B1(new_n807), .B2(G317), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT121), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT120), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1118), .A2(KEYINPUT52), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(KEYINPUT52), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n806), .B1(new_n821), .B2(new_n810), .C1(new_n443), .C2(new_n813), .ZN(new_n1121));
  INV_X1    g0921(.A(G294), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n290), .B1(new_n1122), .B2(new_n798), .C1(new_n802), .C2(new_n424), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1121), .B(new_n1123), .C1(G322), .C2(new_n1081), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1119), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n813), .A2(new_n293), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n840), .B1(new_n262), .B2(new_n798), .C1(new_n802), .C2(new_n268), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(G68), .C2(new_n974), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n797), .A2(G159), .B1(new_n807), .B2(G150), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT51), .Z(new_n1130));
  AOI21_X1  g0930(.A(new_n770), .B1(new_n1081), .B2(G143), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT122), .Z(new_n1134));
  AOI211_X1 g0934(.A(new_n783), .B(new_n1115), .C1(new_n1134), .C2(new_n780), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1111), .A2(new_n763), .B1(new_n1113), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1112), .A2(new_n1136), .ZN(G390));
  AOI21_X1  g0937(.A(new_n949), .B1(new_n925), .B2(new_n934), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n945), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n865), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n732), .B2(new_n864), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1138), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n756), .A2(new_n945), .A3(G330), .A4(new_n866), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n916), .A2(new_n925), .A3(KEYINPUT39), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT39), .B1(new_n925), .B2(new_n934), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n949), .B1(new_n943), .B2(new_n945), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1142), .B(new_n1143), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n948), .A2(new_n950), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1140), .B1(new_n739), .B2(new_n869), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1150), .A2(new_n1139), .B1(new_n392), .B2(new_n698), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n732), .A2(new_n864), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n945), .B1(new_n1152), .B2(new_n1140), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1149), .A2(new_n1151), .B1(new_n1153), .B2(new_n1138), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n880), .A2(new_n889), .A3(G330), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1148), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(new_n762), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1149), .A2(new_n777), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n859), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n764), .B1(new_n320), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n843), .A2(new_n1122), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n802), .A2(new_n314), .B1(new_n798), .B2(new_n356), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G283), .B2(new_n807), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1126), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n294), .B(new_n811), .C1(G116), .C2(new_n797), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1163), .A2(new_n854), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n974), .A2(G150), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT53), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n797), .A2(G132), .ZN(new_n1169));
  INV_X1    g0969(.A(G128), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1169), .B1(new_n808), .B2(new_n1170), .C1(new_n802), .C2(new_n976), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n813), .A2(new_n790), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT54), .B(G143), .Z(new_n1173));
  AOI21_X1  g0973(.A(new_n290), .B1(new_n799), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n268), .B2(new_n804), .ZN(new_n1175));
  OR4_X1    g0975(.A1(new_n1168), .A2(new_n1171), .A3(new_n1172), .A4(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n817), .A2(G125), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1161), .A2(new_n1166), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1160), .B1(new_n1178), .B2(new_n780), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1157), .B1(new_n1158), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n663), .A2(new_n880), .A3(G330), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n954), .A2(new_n691), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n756), .A2(G330), .A3(new_n866), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1139), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n1155), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n943), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n754), .B1(new_n609), .B2(new_n698), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n877), .A2(new_n879), .ZN(new_n1188));
  OAI211_X1 g0988(.A(G330), .B(new_n866), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1139), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1182), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n1148), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(KEYINPUT123), .A3(new_n719), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1192), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1156), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT123), .B1(new_n1193), .B2(new_n719), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1180), .B1(new_n1197), .B2(new_n1198), .ZN(G378));
  INV_X1    g0999(.A(new_n1182), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1156), .B2(new_n1195), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n941), .B1(new_n936), .B2(new_n935), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n902), .A2(new_n915), .A3(new_n892), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT38), .B1(new_n922), .B2(new_n924), .ZN(new_n1204));
  OAI21_X1  g1004(.A(KEYINPUT104), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n916), .A2(new_n925), .A3(new_n926), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n890), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1202), .B1(new_n1207), .B2(KEYINPUT40), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n308), .A2(new_n309), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n338), .A2(new_n339), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n271), .A2(new_n898), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1211), .B(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1213), .B(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1208), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n953), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1216), .B(new_n1202), .C1(new_n1207), .C2(KEYINPUT40), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1219), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1222));
  OAI211_X1 g1022(.A(KEYINPUT57), .B(new_n1201), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1220), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n929), .A2(new_n930), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1216), .B1(new_n1225), .B2(new_n1202), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n953), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1227), .A2(new_n1228), .B1(new_n1200), .B2(new_n1193), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1223), .B(new_n719), .C1(new_n1229), .C2(KEYINPUT57), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n763), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n770), .A2(new_n274), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n851), .A2(new_n804), .B1(new_n810), .B2(new_n293), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n817), .C2(G283), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT124), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n984), .A2(new_n314), .B1(new_n322), .B2(new_n798), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n802), .A2(new_n356), .B1(new_n808), .B2(new_n443), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(G68), .C2(new_n825), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1235), .A2(KEYINPUT58), .A3(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(G33), .A2(G41), .ZN(new_n1240));
  INV_X1    g1040(.A(G124), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1240), .B1(new_n790), .B2(new_n804), .C1(new_n789), .C2(new_n1241), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n801), .A2(G132), .B1(new_n807), .B2(G125), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n797), .A2(G128), .B1(G137), .B2(new_n799), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n825), .A2(G150), .B1(new_n974), .B2(new_n1173), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1242), .B1(KEYINPUT59), .B2(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1240), .A2(G50), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1247), .A2(new_n1248), .B1(new_n1232), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1239), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT58), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n780), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1253), .B(new_n764), .C1(G50), .C2(new_n1159), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1217), .B2(new_n777), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1231), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1230), .A2(new_n1257), .ZN(G375));
  AND2_X1   g1058(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n943), .A2(new_n1185), .B1(new_n1259), .B2(new_n1190), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT125), .B1(new_n1260), .B2(new_n762), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1186), .A2(new_n1191), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n763), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n764), .B1(G68), .B2(new_n1159), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n843), .A2(new_n424), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n443), .A2(new_n802), .B1(new_n984), .B2(new_n821), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G294), .B2(new_n807), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n294), .B(new_n972), .C1(G107), .C2(new_n799), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n825), .A2(new_n492), .B1(new_n974), .B2(G97), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n843), .A2(new_n1170), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n851), .A2(new_n804), .B1(new_n810), .B2(new_n790), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G50), .B2(new_n825), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1173), .A2(new_n801), .B1(new_n807), .B2(G132), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n976), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n797), .A2(new_n1276), .B1(G150), .B2(new_n799), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1274), .A2(new_n1275), .A3(new_n557), .A4(new_n1277), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1266), .A2(new_n1271), .B1(new_n1272), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1265), .B1(new_n1279), .B2(new_n780), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n945), .B2(new_n778), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1261), .A2(new_n1264), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1186), .A2(new_n1191), .A3(new_n1182), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1195), .A2(new_n1031), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(G381));
  INV_X1    g1086(.A(G390), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1070), .A2(new_n835), .A3(new_n1107), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n874), .A3(new_n1289), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1290), .A2(G387), .A3(G381), .ZN(new_n1291));
  INV_X1    g1091(.A(G378), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1257), .A4(new_n1230), .ZN(G407));
  NAND2_X1  g1093(.A1(new_n697), .A2(G213), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G407), .B(G213), .C1(G375), .C2(new_n1296), .ZN(G409));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G387), .A2(new_n1287), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(G393), .B(new_n835), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G390), .B(new_n998), .C1(new_n1032), .C2(new_n1065), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1300), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1230), .A2(G378), .A3(new_n1257), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1031), .B(new_n1201), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(new_n1231), .A3(new_n1256), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1198), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(new_n1196), .A3(new_n1194), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(new_n1310), .A3(new_n1180), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1295), .B1(new_n1306), .B2(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1186), .A2(new_n1182), .A3(KEYINPUT60), .A4(new_n1191), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n719), .ZN(new_n1314));
  OAI21_X1  g1114(.A(KEYINPUT60), .B1(new_n1260), .B2(new_n1182), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1284), .B2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT126), .B1(new_n1316), .B2(new_n1282), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT60), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1284), .B1(new_n1192), .B2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(new_n719), .A3(new_n1313), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1283), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1317), .A2(new_n1322), .A3(G384), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1283), .A2(new_n1320), .A3(new_n1321), .A4(new_n874), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1295), .A2(G2897), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1323), .A2(G2897), .A3(new_n1295), .A4(new_n1324), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1305), .B1(new_n1312), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT62), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(new_n1312), .B2(new_n1325), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1312), .A2(new_n1331), .A3(new_n1325), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1304), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1304), .B(new_n1305), .C1(new_n1312), .C2(new_n1329), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT63), .B1(new_n1312), .B2(new_n1325), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1325), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1298), .B1(new_n1335), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1330), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1337), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1325), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1341), .A2(new_n1342), .A3(new_n1304), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1334), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1345), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1344), .B(KEYINPUT127), .C1(new_n1346), .C2(new_n1304), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1340), .A2(new_n1347), .ZN(G405));
  NAND2_X1  g1148(.A1(G375), .A2(new_n1292), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1306), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1350), .B(new_n1325), .ZN(new_n1351));
  XOR2_X1   g1151(.A(new_n1351), .B(new_n1304), .Z(G402));
endmodule


