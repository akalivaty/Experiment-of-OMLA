//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986;
  NAND2_X1  g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  OR2_X1    g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT9), .ZN(new_n205));
  OAI211_X1 g004(.A(new_n202), .B(new_n203), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n203), .A2(new_n202), .ZN(new_n207));
  INV_X1    g006(.A(G57gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G64gat), .ZN(new_n209));
  INV_X1    g008(.A(G64gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G57gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n202), .A2(new_n205), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n207), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT91), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n206), .A2(KEYINPUT91), .A3(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT21), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G231gat), .ZN(new_n222));
  INV_X1    g021(.A(G233gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n221), .B(new_n224), .Z(new_n225));
  INV_X1    g024(.A(G127gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G183gat), .B(G211gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n225), .A2(new_n226), .ZN(new_n230));
  OR3_X1    g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n228), .B2(new_n230), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n206), .A2(KEYINPUT91), .A3(new_n214), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT91), .B1(new_n206), .B2(new_n214), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G1gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT16), .ZN(new_n238));
  INV_X1    g037(.A(G15gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G22gat), .ZN(new_n240));
  INV_X1    g039(.A(G22gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G15gat), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n238), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(G1gat), .B1(new_n240), .B2(new_n242), .ZN(new_n244));
  OAI21_X1  g043(.A(G8gat), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n241), .A2(G15gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n239), .A2(G22gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n237), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G8gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n238), .A2(new_n240), .A3(new_n242), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n251), .A3(KEYINPUT85), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT85), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n243), .A2(new_n244), .A3(G8gat), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n249), .B1(new_n248), .B2(new_n250), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n236), .A2(KEYINPUT21), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT92), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G155gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n258), .B(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n233), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G190gat), .B(G218gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT7), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT7), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(KEYINPUT93), .A3(G85gat), .A4(G92gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G99gat), .ZN(new_n271));
  INV_X1    g070(.A(G106gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT94), .ZN(new_n274));
  NAND2_X1  g073(.A1(G99gat), .A2(G106gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G85gat), .ZN(new_n277));
  INV_X1    g076(.A(G92gat), .ZN(new_n278));
  AOI22_X1  g077(.A1(KEYINPUT8), .A2(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n270), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n274), .B1(new_n273), .B2(new_n275), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n280), .A2(new_n281), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G29gat), .ZN(new_n285));
  INV_X1    g084(.A(G36gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT14), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT14), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(G29gat), .B2(G36gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT83), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT83), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n287), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G29gat), .A2(G36gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(KEYINPUT84), .A2(G29gat), .A3(G36gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n291), .A2(new_n293), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT15), .ZN(new_n301));
  OR2_X1    g100(.A1(G43gat), .A2(G50gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(G43gat), .A2(G50gat), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n301), .A3(new_n303), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n305), .A2(new_n289), .A3(new_n287), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n304), .A2(new_n298), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n300), .A2(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n284), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(G232gat), .A2(G233gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(KEYINPUT41), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n312));
  INV_X1    g111(.A(new_n304), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n292), .B1(new_n287), .B2(new_n289), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(new_n298), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n315), .B2(new_n293), .ZN(new_n316));
  INV_X1    g115(.A(new_n290), .ZN(new_n317));
  AND4_X1   g116(.A1(new_n313), .A2(new_n317), .A3(new_n299), .A4(new_n305), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n312), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n307), .A2(new_n317), .A3(new_n305), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n287), .A2(new_n289), .A3(new_n292), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n321), .A2(new_n314), .A3(new_n298), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n320), .B(KEYINPUT17), .C1(new_n322), .C2(new_n313), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n323), .A3(new_n284), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n265), .B1(new_n311), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n265), .A3(new_n324), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n310), .A2(KEYINPUT41), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(G134gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n325), .B2(KEYINPUT95), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n328), .B(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n231), .A2(new_n232), .A3(new_n261), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n263), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G120gat), .B(G148gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G176gat), .B(G204gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT99), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n236), .A2(new_n284), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n280), .A2(new_n281), .ZN(new_n342));
  INV_X1    g141(.A(new_n281), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n343), .A2(new_n270), .A3(new_n276), .A4(new_n279), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n342), .A2(new_n344), .B1(new_n206), .B2(new_n214), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G230gat), .A2(G233gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT98), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT10), .B1(new_n282), .B2(new_n283), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT96), .B1(new_n351), .B2(new_n219), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT96), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT10), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n342), .B2(new_n344), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n236), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n345), .B1(new_n236), .B2(new_n284), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n352), .B(new_n356), .C1(new_n357), .C2(KEYINPUT10), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n348), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n340), .B1(new_n350), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT98), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n349), .B(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n354), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n365), .A2(KEYINPUT97), .A3(new_n352), .A4(new_n356), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT97), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n358), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n368), .A3(new_n348), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n369), .A3(new_n339), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n336), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G113gat), .B(G141gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G169gat), .B(G197gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT12), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n320), .B1(new_n322), .B2(new_n313), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n252), .A3(new_n256), .ZN(new_n381));
  NAND2_X1  g180(.A1(G229gat), .A2(G233gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n254), .A2(new_n255), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n319), .A2(new_n323), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT18), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT88), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n379), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n245), .A2(new_n251), .A3(KEYINPUT85), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT85), .B1(new_n245), .B2(new_n251), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n308), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n381), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n382), .B(KEYINPUT13), .Z(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(KEYINPUT86), .A3(new_n394), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n386), .A2(KEYINPUT18), .A3(new_n382), .A4(new_n381), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT18), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n319), .A2(new_n323), .A3(new_n385), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(new_n383), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT88), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n399), .A3(new_n400), .A4(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n397), .A2(new_n403), .A3(new_n400), .A4(new_n398), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n406), .A2(new_n407), .A3(new_n379), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n406), .B2(new_n379), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT89), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT89), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n412), .B(new_n405), .C1(new_n408), .C2(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT72), .ZN(new_n415));
  INV_X1    g214(.A(G169gat), .ZN(new_n416));
  INV_X1    g215(.A(G176gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT23), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT23), .ZN(new_n421));
  NAND2_X1  g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT24), .ZN(new_n424));
  INV_X1    g223(.A(G183gat), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n424), .A2(new_n425), .A3(G190gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  INV_X1    g226(.A(G190gat), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n420), .A2(KEYINPUT64), .A3(new_n421), .A4(new_n422), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT25), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n423), .A2(new_n430), .A3(KEYINPUT25), .A4(new_n432), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT28), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT27), .B(G183gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT65), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n425), .A2(KEYINPUT27), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n428), .B1(new_n441), .B2(KEYINPUT65), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n437), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(KEYINPUT28), .A3(new_n428), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n422), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(KEYINPUT26), .B2(new_n418), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n418), .A2(KEYINPUT26), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n447), .A2(new_n448), .B1(G183gat), .B2(G190gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n436), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n434), .A2(new_n435), .B1(new_n445), .B2(new_n449), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT68), .ZN(new_n455));
  INV_X1    g254(.A(G120gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G113gat), .ZN(new_n457));
  INV_X1    g256(.A(G113gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G120gat), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT1), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G134gat), .ZN(new_n464));
  OAI211_X1 g263(.A(G127gat), .B(new_n464), .C1(new_n460), .C2(KEYINPUT66), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n226), .A2(G134gat), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n455), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G227gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n223), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n465), .A2(new_n466), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n461), .A3(new_n462), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n476), .A3(KEYINPUT68), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT32), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G43gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT69), .ZN(new_n483));
  INV_X1    g282(.A(G71gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(new_n271), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n479), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n486), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n478), .B(KEYINPUT32), .C1(new_n480), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT71), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n436), .A2(new_n450), .A3(KEYINPUT68), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT68), .B1(new_n436), .B2(new_n450), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n492), .A2(new_n493), .A3(new_n476), .ZN(new_n494));
  INV_X1    g293(.A(new_n477), .ZN(new_n495));
  OAI22_X1  g294(.A1(new_n494), .A2(new_n495), .B1(new_n471), .B2(new_n223), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT70), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(KEYINPUT34), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n491), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n472), .B1(new_n470), .B2(new_n477), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n501), .A2(KEYINPUT71), .A3(new_n498), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n490), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT34), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(KEYINPUT70), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n496), .A2(new_n491), .A3(new_n499), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT71), .B1(new_n501), .B2(new_n498), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(new_n487), .A3(new_n489), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n504), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n506), .B1(new_n504), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n415), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G197gat), .B(G204gat), .ZN(new_n516));
  INV_X1    g315(.A(G211gat), .ZN(new_n517));
  INV_X1    g316(.A(G218gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n516), .B1(KEYINPUT22), .B2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G211gat), .B(G218gat), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G226gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(new_n223), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n454), .B2(KEYINPUT29), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT73), .B1(new_n451), .B2(new_n524), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528));
  AOI211_X1 g327(.A(new_n528), .B(new_n525), .C1(new_n436), .C2(new_n450), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n522), .B(new_n526), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n522), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT29), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n524), .B1(new_n451), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n454), .A2(new_n525), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n535), .A3(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(KEYINPUT73), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n528), .B1(new_n454), .B2(new_n525), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT74), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n539), .A2(new_n540), .A3(new_n522), .A4(new_n526), .ZN(new_n541));
  XOR2_X1   g340(.A(G8gat), .B(G36gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT75), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT76), .ZN(new_n544));
  XNOR2_X1  g343(.A(G64gat), .B(G92gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(KEYINPUT37), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n536), .A2(new_n541), .A3(KEYINPUT37), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT38), .ZN(new_n552));
  XNOR2_X1  g351(.A(G1gat), .B(G29gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT0), .ZN(new_n554));
  XNOR2_X1  g353(.A(G57gat), .B(G85gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n554), .B(new_n555), .Z(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT78), .ZN(new_n559));
  INV_X1    g358(.A(G141gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G148gat), .ZN(new_n561));
  INV_X1    g360(.A(G148gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G141gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G155gat), .A2(G162gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT2), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n559), .B1(new_n567), .B2(KEYINPUT79), .ZN(new_n568));
  XNOR2_X1  g367(.A(G155gat), .B(G162gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n561), .A2(new_n563), .B1(KEYINPUT2), .B2(new_n565), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n559), .B(new_n569), .C1(new_n567), .C2(KEYINPUT79), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT3), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(KEYINPUT3), .A3(new_n573), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n476), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n474), .A2(new_n574), .A3(new_n475), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G225gat), .A2(G233gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n469), .A2(KEYINPUT4), .A3(new_n574), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n578), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT5), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT5), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n572), .A2(new_n573), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n476), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n579), .ZN(new_n590));
  INV_X1    g389(.A(new_n582), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n584), .ZN(new_n593));
  AOI211_X1 g392(.A(new_n556), .B(new_n558), .C1(new_n586), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n586), .A2(new_n593), .ZN(new_n595));
  INV_X1    g394(.A(new_n556), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n557), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n586), .A2(new_n556), .A3(new_n593), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n536), .A2(new_n541), .ZN(new_n600));
  INV_X1    g399(.A(new_n546), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT38), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n539), .A2(new_n531), .A3(new_n526), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n522), .B1(new_n533), .B2(new_n534), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(KEYINPUT37), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n549), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n552), .A2(new_n599), .A3(new_n602), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n522), .B1(new_n576), .B2(new_n532), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n575), .B1(new_n531), .B2(KEYINPUT29), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n588), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G78gat), .B(G106gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G228gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n241), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT31), .B(G50gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n613), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT30), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n600), .A2(KEYINPUT30), .A3(new_n601), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n547), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n624), .A3(new_n591), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n625), .A2(new_n556), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT81), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n623), .A2(new_n591), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT39), .B1(new_n590), .B2(new_n591), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n626), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n592), .A2(new_n584), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n596), .B1(new_n633), .B2(new_n585), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n631), .B1(new_n591), .B2(new_n623), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n625), .A2(new_n556), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n627), .B(new_n628), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n632), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n618), .B1(new_n622), .B2(new_n638), .ZN(new_n639));
  AOI211_X1 g438(.A(new_n619), .B(new_n546), .C1(new_n536), .C2(new_n541), .ZN(new_n640));
  INV_X1    g439(.A(new_n547), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT77), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n634), .A2(new_n598), .A3(new_n558), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n595), .A2(new_n596), .A3(new_n557), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT77), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n621), .A2(new_n646), .A3(new_n547), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n642), .A2(new_n645), .A3(new_n647), .A4(new_n620), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n608), .A2(new_n639), .B1(new_n648), .B2(new_n618), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n415), .B(KEYINPUT36), .C1(new_n511), .C2(new_n512), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n515), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n511), .A2(new_n512), .ZN(new_n652));
  INV_X1    g451(.A(new_n648), .ZN(new_n653));
  INV_X1    g452(.A(new_n618), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n511), .A2(new_n512), .A3(new_n618), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n622), .A2(new_n599), .A3(KEYINPUT35), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n655), .A2(KEYINPUT35), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n414), .B1(new_n651), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT90), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n504), .A2(new_n510), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n497), .A2(KEYINPUT34), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n504), .A2(new_n506), .A3(new_n510), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n665), .A3(new_n654), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT35), .B1(new_n666), .B2(new_n648), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n656), .A2(new_n657), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n515), .A2(new_n649), .A3(new_n650), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(KEYINPUT90), .A3(new_n414), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n373), .B1(new_n661), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n599), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT100), .B(G1gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1324gat));
  AOI21_X1  g475(.A(KEYINPUT90), .B1(new_n671), .B2(new_n414), .ZN(new_n677));
  INV_X1    g476(.A(new_n414), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n660), .B(new_n678), .C1(new_n669), .C2(new_n670), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n622), .B(new_n372), .C1(new_n677), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G8gat), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT104), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685));
  INV_X1    g484(.A(new_n683), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n673), .A2(new_n685), .A3(new_n622), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n682), .B(KEYINPUT102), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(KEYINPUT103), .B(new_n689), .C1(new_n680), .C2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n661), .A2(new_n672), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n694), .A2(new_n622), .A3(new_n372), .A4(new_n690), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT103), .B1(new_n695), .B2(new_n689), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n681), .B(new_n688), .C1(new_n693), .C2(new_n696), .ZN(G1325gat));
  NAND2_X1  g496(.A1(new_n673), .A2(new_n652), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n239), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n515), .A2(new_n650), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G15gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n673), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n699), .A2(new_n700), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n704), .ZN(new_n706));
  AOI21_X1  g505(.A(G15gat), .B1(new_n673), .B2(new_n652), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT106), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(G1326gat));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n673), .A2(new_n710), .A3(new_n618), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n618), .B(new_n372), .C1(new_n677), .C2(new_n679), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT107), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n711), .A2(new_n713), .A3(new_n715), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1327gat));
  NAND2_X1  g518(.A1(new_n263), .A2(new_n335), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n371), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n334), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n694), .A2(new_n285), .A3(new_n599), .A4(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n334), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n671), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n334), .B1(new_n669), .B2(new_n670), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n410), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n723), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n645), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n725), .A2(new_n726), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n727), .A2(new_n738), .A3(new_n739), .ZN(G1328gat));
  NAND4_X1  g539(.A1(new_n694), .A2(new_n286), .A3(new_n622), .A4(new_n724), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  INV_X1    g541(.A(new_n622), .ZN(new_n743));
  OAI21_X1  g542(.A(G36gat), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(G1329gat));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n701), .A3(new_n733), .A4(new_n736), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G43gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT108), .ZN(new_n749));
  INV_X1    g548(.A(new_n652), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(G43gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n694), .A2(new_n724), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n749), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n748), .B(new_n752), .C1(KEYINPUT108), .C2(KEYINPUT47), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1330gat));
  NOR2_X1   g556(.A1(new_n654), .A2(G50gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n694), .A2(new_n724), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT48), .B1(new_n759), .B2(KEYINPUT109), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n731), .A2(new_n618), .A3(new_n733), .A4(new_n736), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G50gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n762), .B(new_n759), .C1(KEYINPUT109), .C2(KEYINPUT48), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1331gat));
  AOI211_X1 g565(.A(new_n410), .B(new_n336), .C1(new_n669), .C2(new_n670), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(new_n371), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n599), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g569(.A(new_n743), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n371), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT110), .ZN(new_n773));
  OR2_X1    g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1333gat));
  AOI21_X1  g574(.A(new_n484), .B1(new_n768), .B2(new_n701), .ZN(new_n776));
  INV_X1    g575(.A(new_n371), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n750), .A2(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n767), .A2(new_n484), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n776), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n776), .B2(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1334gat));
  NOR2_X1   g583(.A1(new_n654), .A2(new_n777), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g586(.A1(new_n720), .A2(new_n735), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n777), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n734), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n645), .ZN(new_n792));
  INV_X1    g591(.A(new_n788), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n671), .A2(new_n728), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n732), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n599), .A2(new_n277), .A3(new_n371), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n792), .B1(new_n799), .B2(new_n800), .ZN(G1336gat));
  NAND4_X1  g600(.A1(new_n731), .A2(new_n622), .A3(new_n733), .A4(new_n790), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n743), .A2(G92gat), .A3(new_n777), .ZN(new_n803));
  AOI22_X1  g602(.A1(G92gat), .A2(new_n802), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n804), .B(new_n805), .ZN(G1337gat));
  INV_X1    g605(.A(new_n701), .ZN(new_n807));
  OAI21_X1  g606(.A(G99gat), .B1(new_n791), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n798), .A2(new_n271), .A3(new_n778), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1338gat));
  AND3_X1   g609(.A1(new_n732), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT51), .B1(new_n732), .B2(new_n793), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n785), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n272), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(KEYINPUT113), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(KEYINPUT113), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n654), .A2(new_n272), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n731), .A2(new_n733), .A3(new_n790), .A4(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n814), .A2(new_n817), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(G106gat), .B1(new_n798), .B2(new_n785), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n818), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n816), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n821), .A2(new_n824), .ZN(G1339gat));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n358), .A2(new_n826), .A3(new_n348), .ZN(new_n827));
  INV_X1    g626(.A(new_n339), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n826), .B1(new_n359), .B2(new_n360), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n369), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(KEYINPUT55), .ZN(new_n832));
  INV_X1    g631(.A(new_n370), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n369), .A2(new_n830), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n827), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n834), .A2(new_n841), .A3(new_n410), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n393), .A2(new_n394), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n382), .B1(new_n386), .B2(new_n381), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n405), .B1(new_n378), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n777), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n728), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n334), .A2(new_n846), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n841), .A3(new_n834), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n720), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n372), .A2(new_n735), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n618), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n622), .A2(new_n645), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n652), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(new_n458), .A3(new_n678), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n645), .B1(new_n853), .B2(new_n854), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n860), .A2(new_n743), .A3(new_n656), .ZN(new_n861));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n410), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n859), .A2(new_n862), .ZN(G1340gat));
  AOI21_X1  g662(.A(G120gat), .B1(new_n861), .B2(new_n371), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n750), .A2(new_n456), .A3(new_n777), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n857), .B2(new_n865), .ZN(G1341gat));
  OAI21_X1  g665(.A(G127gat), .B1(new_n858), .B2(new_n720), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n861), .A2(new_n226), .A3(new_n721), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1342gat));
  NAND3_X1  g668(.A1(new_n861), .A2(new_n464), .A3(new_n728), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n858), .B2(new_n334), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(G1343gat));
  NOR3_X1   g673(.A1(new_n701), .A2(new_n654), .A3(new_n622), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n860), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n414), .A2(new_n560), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n856), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n701), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  XOR2_X1   g680(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n882));
  OAI21_X1  g681(.A(new_n370), .B1(new_n831), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n838), .B2(new_n840), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n847), .B1(new_n414), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n851), .B1(new_n885), .B2(new_n728), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n720), .ZN(new_n887));
  AOI211_X1 g686(.A(new_n881), .B(new_n654), .C1(new_n887), .C2(new_n854), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n654), .B1(new_n853), .B2(new_n854), .ZN(new_n889));
  XNOR2_X1  g688(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n880), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n410), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n878), .B1(new_n895), .B2(G141gat), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n560), .B1(new_n894), .B2(new_n414), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n876), .B2(new_n877), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n896), .A2(new_n897), .B1(new_n898), .B2(new_n899), .ZN(G1344gat));
  NOR3_X1   g699(.A1(new_n336), .A2(new_n414), .A3(new_n371), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n654), .B1(new_n903), .B2(KEYINPUT118), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT118), .B(new_n901), .C1(new_n886), .C2(new_n720), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n889), .A2(new_n891), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n777), .B1(new_n880), .B2(KEYINPUT117), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(KEYINPUT117), .B2(new_n880), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT59), .B(G148gat), .C1(new_n910), .C2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n876), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n562), .A3(new_n371), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n562), .B1(new_n894), .B2(new_n371), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n913), .B(new_n915), .C1(new_n916), .C2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g716(.A(G155gat), .B1(new_n914), .B2(new_n721), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n721), .A2(G155gat), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT119), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n918), .B1(new_n894), .B2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n893), .B2(new_n334), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n331), .A3(new_n728), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1347gat));
  NAND2_X1  g723(.A1(new_n853), .A2(new_n854), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n743), .A2(new_n599), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n656), .A3(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n410), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n926), .B(KEYINPUT120), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(new_n750), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n855), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(new_n416), .A3(new_n678), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n929), .A2(new_n933), .ZN(G1348gat));
  NOR3_X1   g733(.A1(new_n932), .A2(new_n417), .A3(new_n777), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT122), .Z(new_n936));
  AOI211_X1 g735(.A(KEYINPUT121), .B(G176gat), .C1(new_n928), .C2(new_n371), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n928), .A2(new_n371), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n417), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n936), .A2(new_n937), .A3(new_n940), .ZN(G1349gat));
  OAI21_X1  g740(.A(G183gat), .B1(new_n932), .B2(new_n720), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n721), .A2(new_n438), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n927), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(KEYINPUT123), .B2(KEYINPUT60), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n942), .A2(new_n944), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n948), .B1(new_n945), .B2(KEYINPUT60), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n947), .B1(new_n949), .B2(new_n946), .ZN(G1350gat));
  NAND3_X1  g749(.A1(new_n928), .A2(new_n428), .A3(new_n728), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n931), .A2(new_n855), .A3(new_n728), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  AND4_X1   g752(.A1(KEYINPUT125), .A2(new_n952), .A3(new_n953), .A4(G190gat), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n428), .B1(new_n955), .B2(KEYINPUT61), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n952), .A2(new_n956), .B1(KEYINPUT125), .B2(new_n953), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n951), .B1(new_n954), .B2(new_n957), .ZN(G1351gat));
  NAND4_X1  g757(.A1(new_n925), .A2(new_n807), .A3(new_n618), .A4(new_n926), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT126), .Z(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n410), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n930), .A2(new_n701), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n901), .B1(new_n886), .B2(new_n720), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT118), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n618), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n881), .B1(new_n966), .B2(new_n905), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n963), .B1(new_n967), .B2(new_n908), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n414), .A2(G197gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n961), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  NOR3_X1   g769(.A1(new_n959), .A2(G204gat), .A3(new_n777), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT62), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n968), .A2(new_n371), .ZN(new_n973));
  INV_X1    g772(.A(G204gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n517), .A3(new_n721), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT63), .ZN(new_n977));
  AOI211_X1 g776(.A(new_n977), .B(new_n517), .C1(new_n968), .C2(new_n721), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n721), .B(new_n962), .C1(new_n907), .C2(new_n909), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n976), .B1(new_n978), .B2(new_n980), .ZN(G1354gat));
  OAI21_X1  g780(.A(new_n728), .B1(new_n968), .B2(KEYINPUT127), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n983));
  AOI211_X1 g782(.A(new_n983), .B(new_n963), .C1(new_n967), .C2(new_n908), .ZN(new_n984));
  OAI21_X1  g783(.A(G218gat), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n960), .A2(new_n518), .A3(new_n728), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


