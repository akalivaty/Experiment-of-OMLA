

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U553 ( .A1(n663), .A2(G8), .ZN(n702) );
  NOR2_X1 U554 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X2 U555 ( .A1(G164), .A2(G1384), .ZN(n728) );
  INV_X1 U556 ( .A(KEYINPUT97), .ZN(n610) );
  NOR2_X1 U557 ( .A1(n702), .A2(n687), .ZN(n518) );
  INV_X1 U558 ( .A(KEYINPUT95), .ZN(n598) );
  INV_X1 U559 ( .A(KEYINPUT96), .ZN(n603) );
  INV_X1 U560 ( .A(KEYINPUT29), .ZN(n654) );
  XNOR2_X1 U561 ( .A(n655), .B(n654), .ZN(n658) );
  INV_X1 U562 ( .A(KEYINPUT99), .ZN(n661) );
  XNOR2_X1 U563 ( .A(n671), .B(KEYINPUT101), .ZN(n672) );
  NAND2_X1 U564 ( .A1(n793), .A2(G54), .ZN(n634) );
  INV_X1 U565 ( .A(KEYINPUT65), .ZN(n525) );
  XNOR2_X1 U566 ( .A(n639), .B(KEYINPUT15), .ZN(n986) );
  INV_X1 U567 ( .A(KEYINPUT40), .ZN(n764) );
  NOR2_X1 U568 ( .A1(G543), .A2(G651), .ZN(n797) );
  NAND2_X1 U569 ( .A1(G89), .A2(n797), .ZN(n519) );
  XOR2_X1 U570 ( .A(KEYINPUT4), .B(n519), .Z(n520) );
  XNOR2_X1 U571 ( .A(n520), .B(KEYINPUT73), .ZN(n523) );
  INV_X1 U572 ( .A(G651), .ZN(n528) );
  XOR2_X1 U573 ( .A(KEYINPUT0), .B(G543), .Z(n572) );
  OR2_X1 U574 ( .A1(n528), .A2(n572), .ZN(n521) );
  XNOR2_X1 U575 ( .A(KEYINPUT67), .B(n521), .ZN(n798) );
  NAND2_X1 U576 ( .A1(G76), .A2(n798), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U578 ( .A(n524), .B(KEYINPUT5), .ZN(n534) );
  NOR2_X1 U579 ( .A1(n572), .A2(G651), .ZN(n526) );
  XNOR2_X2 U580 ( .A(n526), .B(n525), .ZN(n793) );
  NAND2_X1 U581 ( .A1(n793), .A2(G51), .ZN(n527) );
  XNOR2_X1 U582 ( .A(n527), .B(KEYINPUT74), .ZN(n531) );
  NOR2_X1 U583 ( .A1(G543), .A2(n528), .ZN(n529) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n529), .Z(n792) );
  NAND2_X1 U585 ( .A1(G63), .A2(n792), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U587 ( .A(KEYINPUT6), .B(n532), .Z(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U589 ( .A(n535), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U590 ( .A(G2105), .ZN(n542) );
  NOR2_X1 U591 ( .A1(n542), .A2(G2104), .ZN(n536) );
  XNOR2_X1 U592 ( .A(n536), .B(KEYINPUT66), .ZN(n591) );
  NAND2_X1 U593 ( .A1(n591), .A2(G126), .ZN(n538) );
  INV_X1 U594 ( .A(KEYINPUT85), .ZN(n537) );
  XNOR2_X1 U595 ( .A(n538), .B(n537), .ZN(n540) );
  AND2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U597 ( .A1(n890), .A2(G114), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n541), .B(KEYINPUT86), .ZN(n547) );
  AND2_X1 U600 ( .A1(n542), .A2(G2104), .ZN(n886) );
  NAND2_X1 U601 ( .A1(G102), .A2(n886), .ZN(n545) );
  NOR2_X1 U602 ( .A1(G2104), .A2(G2105), .ZN(n543) );
  XOR2_X1 U603 ( .A(KEYINPUT17), .B(n543), .Z(n712) );
  NAND2_X1 U604 ( .A1(G138), .A2(n712), .ZN(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X2 U606 ( .A1(n547), .A2(n546), .ZN(G164) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U608 ( .A1(G64), .A2(n792), .ZN(n549) );
  NAND2_X1 U609 ( .A1(G52), .A2(n793), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n797), .A2(G90), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n550), .B(KEYINPUT68), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G77), .A2(n798), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U616 ( .A1(n555), .A2(n554), .ZN(G171) );
  INV_X1 U617 ( .A(G171), .ZN(G301) );
  NAND2_X1 U618 ( .A1(G91), .A2(n797), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G78), .A2(n798), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G65), .A2(n792), .ZN(n558) );
  XNOR2_X1 U622 ( .A(KEYINPUT69), .B(n558), .ZN(n559) );
  NOR2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n793), .A2(G53), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(G299) );
  NAND2_X1 U626 ( .A1(G88), .A2(n797), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G75), .A2(n798), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U629 ( .A1(G62), .A2(n792), .ZN(n566) );
  NAND2_X1 U630 ( .A1(G50), .A2(n793), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U632 ( .A1(n568), .A2(n567), .ZN(G166) );
  INV_X1 U633 ( .A(G166), .ZN(G303) );
  NAND2_X1 U634 ( .A1(G49), .A2(n793), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U637 ( .A1(n792), .A2(n571), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(G87), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(G288) );
  NAND2_X1 U640 ( .A1(G86), .A2(n797), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G61), .A2(n792), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n798), .A2(G73), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT2), .B(n577), .Z(n578) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n793), .A2(G48), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(G305) );
  AND2_X1 U648 ( .A1(n798), .A2(G72), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G85), .A2(n797), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G47), .A2(n793), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n792), .A2(G60), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(G290) );
  NAND2_X1 U655 ( .A1(n890), .A2(G113), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G101), .A2(n886), .ZN(n588) );
  XOR2_X1 U657 ( .A(KEYINPUT23), .B(n588), .Z(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n832) );
  NAND2_X1 U659 ( .A1(n712), .A2(G137), .ZN(n594) );
  INV_X1 U660 ( .A(n591), .ZN(n592) );
  INV_X1 U661 ( .A(n592), .ZN(n891) );
  NAND2_X1 U662 ( .A1(G125), .A2(n891), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n831) );
  INV_X1 U664 ( .A(G40), .ZN(n595) );
  OR2_X1 U665 ( .A1(n831), .A2(n595), .ZN(n596) );
  OR2_X1 U666 ( .A1(n832), .A2(n596), .ZN(n729) );
  INV_X1 U667 ( .A(n729), .ZN(n597) );
  NAND2_X2 U668 ( .A1(n728), .A2(n597), .ZN(n663) );
  NOR2_X1 U669 ( .A1(G2084), .A2(n663), .ZN(n678) );
  NOR2_X1 U670 ( .A1(G1966), .A2(n702), .ZN(n676) );
  NOR2_X1 U671 ( .A1(n678), .A2(n676), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n599), .B(n598), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n600), .A2(G8), .ZN(n601) );
  XNOR2_X1 U674 ( .A(KEYINPUT30), .B(n601), .ZN(n602) );
  NOR2_X2 U675 ( .A1(n602), .A2(G168), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(n608) );
  NAND2_X1 U677 ( .A1(G1961), .A2(n663), .ZN(n606) );
  INV_X1 U678 ( .A(n663), .ZN(n642) );
  XOR2_X1 U679 ( .A(G2078), .B(KEYINPUT25), .Z(n924) );
  NAND2_X1 U680 ( .A1(n642), .A2(n924), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n656) );
  NAND2_X1 U682 ( .A1(G301), .A2(n656), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U684 ( .A(n609), .B(KEYINPUT31), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(n610), .ZN(n660) );
  INV_X1 U686 ( .A(G299), .ZN(n971) );
  NAND2_X1 U687 ( .A1(n642), .A2(G2072), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT27), .ZN(n614) );
  INV_X1 U689 ( .A(G1956), .ZN(n972) );
  NOR2_X1 U690 ( .A1(n972), .A2(n642), .ZN(n613) );
  NOR2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n649) );
  NOR2_X1 U692 ( .A1(n971), .A2(n649), .ZN(n616) );
  XNOR2_X1 U693 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n616), .B(n615), .ZN(n653) );
  NAND2_X1 U695 ( .A1(n797), .A2(G81), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n617), .B(KEYINPUT12), .ZN(n619) );
  NAND2_X1 U697 ( .A1(G68), .A2(n798), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n621) );
  XOR2_X1 U699 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n620) );
  XNOR2_X1 U700 ( .A(n621), .B(n620), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n792), .A2(G56), .ZN(n622) );
  XOR2_X1 U702 ( .A(KEYINPUT14), .B(n622), .Z(n623) );
  NOR2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n793), .A2(G43), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n983) );
  INV_X1 U706 ( .A(G1996), .ZN(n717) );
  NOR2_X1 U707 ( .A1(n663), .A2(n717), .ZN(n628) );
  XOR2_X1 U708 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n627) );
  XNOR2_X1 U709 ( .A(n628), .B(n627), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n663), .A2(G1341), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U712 ( .A1(n983), .A2(n631), .ZN(n641) );
  NAND2_X1 U713 ( .A1(G66), .A2(n792), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G92), .A2(n797), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G79), .A2(n798), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT72), .B(n634), .Z(n635) );
  NOR2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U720 ( .A1(n641), .A2(n986), .ZN(n640) );
  XOR2_X1 U721 ( .A(n640), .B(KEYINPUT94), .Z(n648) );
  NAND2_X1 U722 ( .A1(n641), .A2(n986), .ZN(n646) );
  NOR2_X1 U723 ( .A1(n642), .A2(G1348), .ZN(n644) );
  NOR2_X1 U724 ( .A1(G2067), .A2(n663), .ZN(n643) );
  NOR2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n971), .A2(n649), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n655) );
  OR2_X1 U731 ( .A1(G301), .A2(n656), .ZN(n657) );
  NAND2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n674) );
  NAND2_X1 U734 ( .A1(n674), .A2(G286), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n662), .B(n661), .ZN(n669) );
  NOR2_X1 U736 ( .A1(G1971), .A2(n702), .ZN(n665) );
  NOR2_X1 U737 ( .A1(G2090), .A2(n663), .ZN(n664) );
  NOR2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U739 ( .A1(n666), .A2(G303), .ZN(n667) );
  XNOR2_X1 U740 ( .A(KEYINPUT100), .B(n667), .ZN(n668) );
  NAND2_X1 U741 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n670), .A2(G8), .ZN(n673) );
  XOR2_X1 U743 ( .A(KEYINPUT32), .B(KEYINPUT102), .Z(n671) );
  XNOR2_X1 U744 ( .A(n673), .B(n672), .ZN(n682) );
  INV_X1 U745 ( .A(n674), .ZN(n675) );
  NOR2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n677), .B(KEYINPUT98), .ZN(n680) );
  NAND2_X1 U748 ( .A1(n678), .A2(G8), .ZN(n679) );
  NAND2_X1 U749 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n696) );
  NOR2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n683) );
  XOR2_X1 U752 ( .A(KEYINPUT103), .B(n683), .Z(n974) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n684) );
  NOR2_X1 U754 ( .A1(n974), .A2(n684), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n696), .A2(n685), .ZN(n686) );
  XNOR2_X1 U756 ( .A(n686), .B(KEYINPUT104), .ZN(n688) );
  NAND2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n975) );
  INV_X1 U758 ( .A(n975), .ZN(n687) );
  AND2_X1 U759 ( .A1(n688), .A2(n518), .ZN(n689) );
  NOR2_X1 U760 ( .A1(n689), .A2(KEYINPUT33), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n974), .A2(KEYINPUT33), .ZN(n690) );
  NOR2_X1 U762 ( .A1(n690), .A2(n702), .ZN(n691) );
  XOR2_X1 U763 ( .A(G1981), .B(G305), .Z(n989) );
  NAND2_X1 U764 ( .A1(n693), .A2(n989), .ZN(n752) );
  INV_X1 U765 ( .A(KEYINPUT105), .ZN(n698) );
  NOR2_X1 U766 ( .A1(G2090), .A2(G303), .ZN(n694) );
  NAND2_X1 U767 ( .A1(G8), .A2(n694), .ZN(n695) );
  NAND2_X1 U768 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(n699) );
  AND2_X1 U770 ( .A1(n699), .A2(n702), .ZN(n704) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XOR2_X1 U772 ( .A(n700), .B(KEYINPUT24), .Z(n701) );
  NOR2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U774 ( .A1(n704), .A2(n703), .ZN(n750) );
  NAND2_X1 U775 ( .A1(G117), .A2(n890), .ZN(n705) );
  XOR2_X1 U776 ( .A(KEYINPUT90), .B(n705), .Z(n708) );
  NAND2_X1 U777 ( .A1(n886), .A2(G105), .ZN(n706) );
  XOR2_X1 U778 ( .A(KEYINPUT38), .B(n706), .Z(n707) );
  NOR2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U780 ( .A1(G129), .A2(n891), .ZN(n709) );
  NAND2_X1 U781 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U782 ( .A(n711), .B(KEYINPUT91), .ZN(n714) );
  BUF_X1 U783 ( .A(n712), .Z(n887) );
  NAND2_X1 U784 ( .A1(G141), .A2(n887), .ZN(n713) );
  NAND2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U786 ( .A(KEYINPUT92), .B(n715), .ZN(n908) );
  NOR2_X1 U787 ( .A1(G1996), .A2(n908), .ZN(n950) );
  INV_X1 U788 ( .A(n908), .ZN(n716) );
  NOR2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n727) );
  NAND2_X1 U790 ( .A1(n890), .A2(G107), .ZN(n719) );
  NAND2_X1 U791 ( .A1(G119), .A2(n891), .ZN(n718) );
  NAND2_X1 U792 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U793 ( .A(KEYINPUT88), .B(n720), .Z(n722) );
  NAND2_X1 U794 ( .A1(n886), .A2(G95), .ZN(n721) );
  NAND2_X1 U795 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U796 ( .A1(G131), .A2(n887), .ZN(n723) );
  XNOR2_X1 U797 ( .A(KEYINPUT89), .B(n723), .ZN(n724) );
  OR2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n898) );
  AND2_X1 U799 ( .A1(n898), .A2(G1991), .ZN(n726) );
  NOR2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n947) );
  NOR2_X1 U801 ( .A1(n728), .A2(n729), .ZN(n757) );
  INV_X1 U802 ( .A(n757), .ZN(n730) );
  NOR2_X1 U803 ( .A1(n947), .A2(n730), .ZN(n754) );
  NOR2_X1 U804 ( .A1(G1991), .A2(n898), .ZN(n959) );
  NOR2_X1 U805 ( .A1(G1986), .A2(G290), .ZN(n731) );
  XNOR2_X1 U806 ( .A(KEYINPUT106), .B(n731), .ZN(n732) );
  NOR2_X1 U807 ( .A1(n959), .A2(n732), .ZN(n733) );
  NOR2_X1 U808 ( .A1(n754), .A2(n733), .ZN(n734) );
  NOR2_X1 U809 ( .A1(n950), .A2(n734), .ZN(n735) );
  XNOR2_X1 U810 ( .A(KEYINPUT39), .B(n735), .ZN(n746) );
  NAND2_X1 U811 ( .A1(G104), .A2(n886), .ZN(n737) );
  NAND2_X1 U812 ( .A1(G140), .A2(n887), .ZN(n736) );
  NAND2_X1 U813 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U814 ( .A(KEYINPUT34), .B(n738), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n890), .A2(G116), .ZN(n740) );
  NAND2_X1 U816 ( .A1(G128), .A2(n891), .ZN(n739) );
  NAND2_X1 U817 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U818 ( .A(n741), .B(KEYINPUT35), .Z(n742) );
  NOR2_X1 U819 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U820 ( .A(KEYINPUT36), .B(n744), .Z(n745) );
  XNOR2_X1 U821 ( .A(KEYINPUT87), .B(n745), .ZN(n901) );
  XNOR2_X1 U822 ( .A(G2067), .B(KEYINPUT37), .ZN(n747) );
  NOR2_X1 U823 ( .A1(n901), .A2(n747), .ZN(n963) );
  NAND2_X1 U824 ( .A1(n757), .A2(n963), .ZN(n756) );
  NAND2_X1 U825 ( .A1(n746), .A2(n756), .ZN(n748) );
  NAND2_X1 U826 ( .A1(n901), .A2(n747), .ZN(n956) );
  NAND2_X1 U827 ( .A1(n748), .A2(n956), .ZN(n749) );
  NAND2_X1 U828 ( .A1(n749), .A2(n757), .ZN(n753) );
  AND2_X1 U829 ( .A1(n750), .A2(n753), .ZN(n751) );
  NAND2_X1 U830 ( .A1(n752), .A2(n751), .ZN(n763) );
  INV_X1 U831 ( .A(n753), .ZN(n761) );
  INV_X1 U832 ( .A(n754), .ZN(n755) );
  NAND2_X1 U833 ( .A1(n756), .A2(n755), .ZN(n759) );
  XNOR2_X1 U834 ( .A(G1986), .B(G290), .ZN(n985) );
  AND2_X1 U835 ( .A1(n985), .A2(n757), .ZN(n758) );
  NOR2_X1 U836 ( .A1(n759), .A2(n758), .ZN(n760) );
  OR2_X1 U837 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U838 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U839 ( .A(n765), .B(n764), .ZN(G329) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U841 ( .A(G57), .ZN(G237) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n766) );
  XNOR2_X1 U843 ( .A(n766), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U844 ( .A(G223), .ZN(n833) );
  NAND2_X1 U845 ( .A1(n833), .A2(G567), .ZN(n767) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  XNOR2_X1 U847 ( .A(G860), .B(KEYINPUT71), .ZN(n773) );
  OR2_X1 U848 ( .A1(n983), .A2(n773), .ZN(G153) );
  NAND2_X1 U849 ( .A1(G868), .A2(G301), .ZN(n769) );
  OR2_X1 U850 ( .A1(n986), .A2(G868), .ZN(n768) );
  NAND2_X1 U851 ( .A1(n769), .A2(n768), .ZN(G284) );
  INV_X1 U852 ( .A(G868), .ZN(n813) );
  NOR2_X1 U853 ( .A1(G286), .A2(n813), .ZN(n770) );
  XOR2_X1 U854 ( .A(KEYINPUT75), .B(n770), .Z(n772) );
  NOR2_X1 U855 ( .A1(G868), .A2(G299), .ZN(n771) );
  NOR2_X1 U856 ( .A1(n772), .A2(n771), .ZN(G297) );
  NAND2_X1 U857 ( .A1(n773), .A2(G559), .ZN(n774) );
  NAND2_X1 U858 ( .A1(n774), .A2(n986), .ZN(n775) );
  XNOR2_X1 U859 ( .A(n775), .B(KEYINPUT76), .ZN(n776) );
  XNOR2_X1 U860 ( .A(KEYINPUT16), .B(n776), .ZN(G148) );
  NOR2_X1 U861 ( .A1(G868), .A2(n983), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G868), .A2(n986), .ZN(n777) );
  NOR2_X1 U863 ( .A1(G559), .A2(n777), .ZN(n778) );
  NOR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(G282) );
  XNOR2_X1 U865 ( .A(G2100), .B(KEYINPUT79), .ZN(n790) );
  NAND2_X1 U866 ( .A1(G111), .A2(n890), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G99), .A2(n886), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U869 ( .A(n782), .B(KEYINPUT77), .ZN(n784) );
  NAND2_X1 U870 ( .A1(G135), .A2(n887), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U872 ( .A1(n891), .A2(G123), .ZN(n785) );
  XOR2_X1 U873 ( .A(KEYINPUT18), .B(n785), .Z(n786) );
  NOR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n955) );
  XNOR2_X1 U875 ( .A(n955), .B(G2096), .ZN(n788) );
  XNOR2_X1 U876 ( .A(n788), .B(KEYINPUT78), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G559), .A2(n986), .ZN(n791) );
  XNOR2_X1 U879 ( .A(n983), .B(n791), .ZN(n810) );
  NOR2_X1 U880 ( .A1(n810), .A2(G860), .ZN(n803) );
  NAND2_X1 U881 ( .A1(G67), .A2(n792), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G55), .A2(n793), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U884 ( .A(KEYINPUT80), .B(n796), .ZN(n802) );
  NAND2_X1 U885 ( .A1(G93), .A2(n797), .ZN(n800) );
  NAND2_X1 U886 ( .A1(G80), .A2(n798), .ZN(n799) );
  NAND2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U888 ( .A1(n802), .A2(n801), .ZN(n812) );
  XOR2_X1 U889 ( .A(n803), .B(n812), .Z(G145) );
  XNOR2_X1 U890 ( .A(n971), .B(G166), .ZN(n809) );
  XOR2_X1 U891 ( .A(n812), .B(G290), .Z(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(G305), .ZN(n805) );
  XNOR2_X1 U893 ( .A(KEYINPUT81), .B(n805), .ZN(n807) );
  XNOR2_X1 U894 ( .A(G288), .B(KEYINPUT19), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n807), .B(n806), .ZN(n808) );
  XNOR2_X1 U896 ( .A(n809), .B(n808), .ZN(n911) );
  XOR2_X1 U897 ( .A(n810), .B(n911), .Z(n811) );
  NAND2_X1 U898 ( .A1(n811), .A2(G868), .ZN(n815) );
  NAND2_X1 U899 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U900 ( .A1(n815), .A2(n814), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n816) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n816), .Z(n817) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U907 ( .A1(G120), .A2(G69), .ZN(n820) );
  NOR2_X1 U908 ( .A1(G237), .A2(n820), .ZN(n821) );
  NAND2_X1 U909 ( .A1(G108), .A2(n821), .ZN(n837) );
  NAND2_X1 U910 ( .A1(G567), .A2(n837), .ZN(n822) );
  XNOR2_X1 U911 ( .A(KEYINPUT84), .B(n822), .ZN(n829) );
  XOR2_X1 U912 ( .A(KEYINPUT82), .B(KEYINPUT22), .Z(n824) );
  NAND2_X1 U913 ( .A1(G132), .A2(G82), .ZN(n823) );
  XNOR2_X1 U914 ( .A(n824), .B(n823), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n825), .A2(G96), .ZN(n826) );
  NOR2_X1 U916 ( .A1(n826), .A2(G218), .ZN(n827) );
  XNOR2_X1 U917 ( .A(n827), .B(KEYINPUT83), .ZN(n838) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n838), .ZN(n828) );
  NAND2_X1 U919 ( .A1(n829), .A2(n828), .ZN(n921) );
  NAND2_X1 U920 ( .A1(G483), .A2(G661), .ZN(n830) );
  NOR2_X1 U921 ( .A1(n921), .A2(n830), .ZN(n836) );
  NAND2_X1 U922 ( .A1(n836), .A2(G36), .ZN(G176) );
  NOR2_X1 U923 ( .A1(n832), .A2(n831), .ZN(G160) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U926 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(G188) );
  XOR2_X1 U929 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U931 ( .A(G132), .ZN(G219) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G82), .ZN(G220) );
  NOR2_X1 U935 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U937 ( .A(G1341), .B(G2454), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n839), .B(G2430), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n840), .B(G1348), .ZN(n846) );
  XOR2_X1 U940 ( .A(G2443), .B(G2427), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2438), .B(G2446), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n844) );
  XOR2_X1 U943 ( .A(G2451), .B(G2435), .Z(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  NAND2_X1 U946 ( .A1(n847), .A2(G14), .ZN(n848) );
  XNOR2_X1 U947 ( .A(KEYINPUT107), .B(n848), .ZN(G401) );
  XOR2_X1 U948 ( .A(G2096), .B(G2100), .Z(n850) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U951 ( .A(KEYINPUT43), .B(G2090), .Z(n852) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U954 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2078), .B(G2084), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(G227) );
  XOR2_X1 U957 ( .A(G1981), .B(G1971), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1966), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n859), .B(G2474), .Z(n861) );
  XNOR2_X1 U961 ( .A(G1956), .B(G1976), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U963 ( .A(KEYINPUT41), .B(G1961), .Z(n863) );
  XNOR2_X1 U964 ( .A(G1996), .B(G1991), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(G229) );
  NAND2_X1 U967 ( .A1(n891), .A2(G124), .ZN(n866) );
  XOR2_X1 U968 ( .A(KEYINPUT109), .B(n866), .Z(n867) );
  XNOR2_X1 U969 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G136), .A2(n887), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U972 ( .A(KEYINPUT110), .B(n870), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G112), .A2(n890), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G100), .A2(n886), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U976 ( .A1(n874), .A2(n873), .ZN(G162) );
  NAND2_X1 U977 ( .A1(G118), .A2(n890), .ZN(n884) );
  NAND2_X1 U978 ( .A1(G130), .A2(n891), .ZN(n875) );
  XNOR2_X1 U979 ( .A(KEYINPUT111), .B(n875), .ZN(n882) );
  NAND2_X1 U980 ( .A1(n887), .A2(G142), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n876), .B(KEYINPUT112), .ZN(n878) );
  NAND2_X1 U982 ( .A1(G106), .A2(n886), .ZN(n877) );
  NAND2_X1 U983 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U984 ( .A(KEYINPUT113), .B(n879), .ZN(n880) );
  XNOR2_X1 U985 ( .A(KEYINPUT45), .B(n880), .ZN(n881) );
  NOR2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n885), .B(G162), .ZN(n897) );
  NAND2_X1 U989 ( .A1(G103), .A2(n886), .ZN(n889) );
  NAND2_X1 U990 ( .A1(G139), .A2(n887), .ZN(n888) );
  NAND2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U992 ( .A1(n890), .A2(G115), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G127), .A2(n891), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n943) );
  XOR2_X1 U997 ( .A(n897), .B(n943), .Z(n900) );
  XOR2_X1 U998 ( .A(G164), .B(n898), .Z(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n901), .B(KEYINPUT46), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1003 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G160), .B(n955), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1008 ( .A(n983), .B(n911), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(G171), .B(n986), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n914), .B(G286), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n915), .ZN(G397) );
  OR2_X1 U1013 ( .A1(n921), .A2(G401), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n921), .ZN(G319) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1022 ( .A(G2084), .B(G34), .Z(n922) );
  XNOR2_X1 U1023 ( .A(KEYINPUT54), .B(n922), .ZN(n938) );
  XNOR2_X1 U1024 ( .A(G2090), .B(G35), .ZN(n936) );
  XOR2_X1 U1025 ( .A(G25), .B(G1991), .Z(n923) );
  NAND2_X1 U1026 ( .A1(n923), .A2(G28), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(G1996), .B(G32), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(n924), .B(G27), .ZN(n925) );
  NOR2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1030 ( .A(KEYINPUT116), .B(n927), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(G2067), .B(G26), .ZN(n929) );
  XNOR2_X1 U1032 ( .A(G33), .B(G2072), .ZN(n928) );
  NOR2_X1 U1033 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1036 ( .A(KEYINPUT53), .B(n934), .ZN(n935) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(n939), .B(KEYINPUT117), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT55), .B(n940), .ZN(n941) );
  INV_X1 U1041 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n968), .ZN(n942) );
  NAND2_X1 U1043 ( .A1(n942), .A2(G11), .ZN(n970) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(KEYINPUT115), .ZN(n965) );
  XOR2_X1 U1045 ( .A(G2072), .B(n943), .Z(n945) );
  XOR2_X1 U1046 ( .A(G164), .B(G2078), .Z(n944) );
  NOR2_X1 U1047 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(KEYINPUT50), .B(n946), .ZN(n948) );
  NAND2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n953) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(n951), .B(KEYINPUT51), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n961) );
  XOR2_X1 U1054 ( .A(G2084), .B(G160), .Z(n954) );
  NOR2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n957) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n965), .B(n964), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n966), .A2(KEYINPUT55), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n1030) );
  XOR2_X1 U1064 ( .A(KEYINPUT56), .B(G16), .Z(n1000) );
  XNOR2_X1 U1065 ( .A(G166), .B(G1971), .ZN(n981) );
  XNOR2_X1 U1066 ( .A(n971), .B(KEYINPUT118), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(n972), .ZN(n979) );
  INV_X1 U1068 ( .A(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1070 ( .A(KEYINPUT119), .B(n977), .Z(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n982), .B(KEYINPUT120), .ZN(n997) );
  XNOR2_X1 U1074 ( .A(G1341), .B(n983), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n995) );
  XNOR2_X1 U1076 ( .A(G1348), .B(n986), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(G171), .B(G1961), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n993) );
  XNOR2_X1 U1079 ( .A(G168), .B(G1966), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1081 ( .A(KEYINPUT57), .B(n991), .Z(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1085 ( .A(KEYINPUT121), .B(n998), .Z(n999) );
  NOR2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1028) );
  XNOR2_X1 U1087 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G1981), .B(G6), .ZN(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(KEYINPUT122), .B(n1003), .Z(n1005) );
  XNOR2_X1 U1091 ( .A(G1956), .B(G20), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(KEYINPUT123), .B(n1006), .Z(n1010) );
  XNOR2_X1 U1094 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1007), .B(G4), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1348), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1098 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n1011) );
  XNOR2_X1 U1099 ( .A(n1012), .B(n1011), .ZN(n1019) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G1986), .B(G24), .Z(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(G1966), .B(G21), .Z(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT126), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(G5), .B(G1961), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1025), .Z(n1026) );
  NOR2_X1 U1113 ( .A1(G16), .A2(n1026), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1116 ( .A(KEYINPUT127), .B(n1031), .ZN(n1032) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1032), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

