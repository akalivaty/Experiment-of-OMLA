

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747;

  XNOR2_X1 U367 ( .A(n373), .B(n358), .ZN(n404) );
  NAND2_X1 U368 ( .A1(n601), .A2(n578), .ZN(n373) );
  INV_X1 U369 ( .A(G953), .ZN(n737) );
  AND2_X1 U370 ( .A1(n374), .A2(n377), .ZN(n345) );
  XNOR2_X2 U371 ( .A(n486), .B(n726), .ZN(n672) );
  NAND2_X2 U372 ( .A1(n500), .A2(n438), .ZN(n501) );
  XNOR2_X2 U373 ( .A(n426), .B(n354), .ZN(n500) );
  INV_X2 U374 ( .A(KEYINPUT69), .ZN(n365) );
  XNOR2_X2 U375 ( .A(n485), .B(n484), .ZN(n726) );
  NOR2_X1 U376 ( .A1(n526), .A2(n625), .ZN(n368) );
  XNOR2_X2 U377 ( .A(n382), .B(KEYINPUT84), .ZN(n703) );
  AND2_X2 U378 ( .A1(n590), .A2(n500), .ZN(n382) );
  XOR2_X2 U379 ( .A(n576), .B(n595), .Z(n642) );
  INV_X1 U380 ( .A(n573), .ZN(n581) );
  INV_X2 U381 ( .A(G128), .ZN(n389) );
  XNOR2_X1 U382 ( .A(n446), .B(n445), .ZN(n573) );
  XNOR2_X1 U383 ( .A(n428), .B(n427), .ZN(n363) );
  XNOR2_X1 U384 ( .A(n365), .B(G101), .ZN(n364) );
  XNOR2_X1 U385 ( .A(G119), .B(G113), .ZN(n428) );
  AND2_X2 U386 ( .A1(n614), .A2(n613), .ZN(n735) );
  XNOR2_X1 U387 ( .A(n417), .B(KEYINPUT32), .ZN(n690) );
  XNOR2_X1 U388 ( .A(n543), .B(n542), .ZN(n705) );
  AND2_X1 U389 ( .A1(n533), .A2(n532), .ZN(n417) );
  BUF_X1 U390 ( .A(n570), .Z(n595) );
  XNOR2_X1 U391 ( .A(n492), .B(n491), .ZN(n570) );
  AND2_X1 U392 ( .A1(n693), .A2(n488), .ZN(n446) );
  XNOR2_X1 U393 ( .A(n724), .B(n364), .ZN(n477) );
  NOR2_X2 U394 ( .A1(n668), .A2(n618), .ZN(n619) );
  XNOR2_X2 U395 ( .A(n503), .B(n439), .ZN(n732) );
  INV_X1 U396 ( .A(G237), .ZN(n487) );
  XNOR2_X1 U397 ( .A(KEYINPUT4), .B(G131), .ZN(n439) );
  AND2_X1 U398 ( .A1(n539), .A2(n350), .ZN(n530) );
  INV_X1 U399 ( .A(n628), .ZN(n419) );
  NAND2_X2 U400 ( .A1(n393), .A2(n390), .ZN(n585) );
  OR2_X1 U401 ( .A1(n681), .A2(n391), .ZN(n390) );
  AND2_X1 U402 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U403 ( .A1(n392), .A2(n488), .ZN(n391) );
  XNOR2_X1 U404 ( .A(n579), .B(n376), .ZN(n620) );
  INV_X1 U405 ( .A(KEYINPUT41), .ZN(n376) );
  NAND2_X1 U406 ( .A1(n402), .A2(n592), .ZN(n401) );
  NAND2_X1 U407 ( .A1(n370), .A2(n369), .ZN(n550) );
  NAND2_X1 U408 ( .A1(n371), .A2(n351), .ZN(n369) );
  NAND2_X1 U409 ( .A1(n705), .A2(n429), .ZN(n370) );
  XNOR2_X1 U410 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U411 ( .A(G137), .B(KEYINPUT77), .ZN(n441) );
  XOR2_X1 U412 ( .A(KEYINPUT101), .B(KEYINPUT5), .Z(n442) );
  XNOR2_X1 U413 ( .A(KEYINPUT48), .B(KEYINPUT89), .ZN(n599) );
  XNOR2_X1 U414 ( .A(G113), .B(G122), .ZN(n415) );
  XNOR2_X1 U415 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n416) );
  XNOR2_X1 U416 ( .A(G143), .B(G131), .ZN(n512) );
  XOR2_X1 U417 ( .A(G140), .B(G104), .Z(n513) );
  XOR2_X1 U418 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n518) );
  XNOR2_X1 U419 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U420 ( .A(KEYINPUT80), .B(G107), .Z(n448) );
  XOR2_X1 U421 ( .A(G137), .B(G140), .Z(n464) );
  INV_X1 U422 ( .A(G146), .ZN(n433) );
  XNOR2_X1 U423 ( .A(n385), .B(G116), .ZN(n505) );
  XNOR2_X1 U424 ( .A(G122), .B(G107), .ZN(n385) );
  NAND2_X1 U425 ( .A1(n573), .A2(n641), .ZN(n411) );
  INV_X1 U426 ( .A(KEYINPUT30), .ZN(n410) );
  XNOR2_X1 U427 ( .A(n524), .B(n423), .ZN(n538) );
  XNOR2_X1 U428 ( .A(n523), .B(n424), .ZN(n423) );
  INV_X1 U429 ( .A(G475), .ZN(n424) );
  NAND2_X1 U430 ( .A1(n414), .A2(n413), .ZN(n575) );
  INV_X1 U431 ( .A(n585), .ZN(n413) );
  XNOR2_X1 U432 ( .A(n585), .B(KEYINPUT1), .ZN(n526) );
  INV_X1 U433 ( .A(n641), .ZN(n388) );
  NAND2_X1 U434 ( .A1(n420), .A2(n383), .ZN(n539) );
  AND2_X1 U435 ( .A1(n384), .A2(n422), .ZN(n383) );
  NAND2_X1 U436 ( .A1(n511), .A2(n488), .ZN(n421) );
  AND2_X1 U437 ( .A1(n539), .A2(n540), .ZN(n578) );
  BUF_X1 U438 ( .A(n526), .Z(n624) );
  NOR2_X1 U439 ( .A1(G953), .A2(G237), .ZN(n516) );
  OR2_X1 U440 ( .A1(n567), .A2(n628), .ZN(n625) );
  NAND2_X1 U441 ( .A1(G234), .A2(G237), .ZN(n494) );
  NAND2_X1 U442 ( .A1(n539), .A2(n538), .ZN(n644) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n580) );
  INV_X1 U444 ( .A(KEYINPUT71), .ZN(n380) );
  NAND2_X1 U445 ( .A1(n567), .A2(n568), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n368), .B(KEYINPUT76), .ZN(n541) );
  NAND2_X1 U447 ( .A1(n425), .A2(G902), .ZN(n422) );
  XNOR2_X1 U448 ( .A(n407), .B(n406), .ZN(n405) );
  XNOR2_X1 U449 ( .A(n444), .B(n443), .ZN(n407) );
  XNOR2_X1 U450 ( .A(G128), .B(G119), .ZN(n453) );
  XOR2_X1 U451 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n454) );
  XNOR2_X1 U452 ( .A(n476), .B(G134), .ZN(n503) );
  XNOR2_X1 U453 ( .A(n386), .B(n505), .ZN(n507) );
  XNOR2_X1 U454 ( .A(n506), .B(KEYINPUT9), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n522), .B(n521), .ZN(n679) );
  XNOR2_X1 U456 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U457 ( .A(n416), .B(n415), .ZN(n519) );
  XNOR2_X1 U458 ( .A(n432), .B(n431), .ZN(n430) );
  XNOR2_X1 U459 ( .A(n464), .B(n450), .ZN(n431) );
  XNOR2_X1 U460 ( .A(n363), .B(KEYINPUT16), .ZN(n485) );
  XNOR2_X1 U461 ( .A(n418), .B(n356), .ZN(n532) );
  XNOR2_X1 U462 ( .A(n372), .B(KEYINPUT102), .ZN(n637) );
  AND2_X1 U463 ( .A1(n541), .A2(n634), .ZN(n372) );
  XNOR2_X1 U464 ( .A(n408), .B(KEYINPUT79), .ZN(n593) );
  NOR2_X1 U465 ( .A1(n575), .A2(n574), .ZN(n412) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n409) );
  NAND2_X1 U467 ( .A1(n570), .A2(n641), .ZN(n426) );
  XNOR2_X1 U468 ( .A(n545), .B(KEYINPUT100), .ZN(n371) );
  NOR2_X1 U469 ( .A1(n603), .A2(n606), .ZN(n571) );
  NAND2_X1 U470 ( .A1(n398), .A2(n397), .ZN(n396) );
  INV_X1 U471 ( .A(G143), .ZN(n687) );
  INV_X1 U472 ( .A(n646), .ZN(n429) );
  BUF_X1 U473 ( .A(n573), .Z(n634) );
  XNOR2_X1 U474 ( .A(KEYINPUT69), .B(G101), .ZN(n346) );
  AND2_X1 U475 ( .A1(n379), .A2(n377), .ZN(n347) );
  AND2_X1 U476 ( .A1(n378), .A2(n377), .ZN(n348) );
  XOR2_X1 U477 ( .A(n530), .B(KEYINPUT109), .Z(n349) );
  AND2_X1 U478 ( .A1(n538), .A2(n419), .ZN(n350) );
  AND2_X1 U479 ( .A1(n429), .A2(n581), .ZN(n351) );
  XOR2_X1 U480 ( .A(KEYINPUT24), .B(G110), .Z(n352) );
  AND2_X1 U481 ( .A1(n569), .A2(n387), .ZN(n353) );
  XOR2_X1 U482 ( .A(KEYINPUT67), .B(KEYINPUT19), .Z(n354) );
  AND2_X1 U483 ( .A1(n371), .A2(n581), .ZN(n355) );
  XOR2_X1 U484 ( .A(n531), .B(KEYINPUT22), .Z(n356) );
  XOR2_X1 U485 ( .A(KEYINPUT68), .B(KEYINPUT0), .Z(n357) );
  XOR2_X1 U486 ( .A(KEYINPUT113), .B(KEYINPUT40), .Z(n358) );
  XOR2_X1 U487 ( .A(n693), .B(n692), .Z(n359) );
  XOR2_X1 U488 ( .A(n679), .B(n678), .Z(n360) );
  XOR2_X1 U489 ( .A(n683), .B(n682), .Z(n361) );
  XNOR2_X1 U490 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n362) );
  AND2_X1 U491 ( .A1(n675), .A2(G953), .ZN(n718) );
  INV_X1 U492 ( .A(n718), .ZN(n377) );
  XNOR2_X1 U493 ( .A(n363), .B(n346), .ZN(n406) );
  XNOR2_X2 U494 ( .A(G110), .B(G104), .ZN(n724) );
  NAND2_X1 U495 ( .A1(n366), .A2(n349), .ZN(n418) );
  XNOR2_X1 U496 ( .A(n366), .B(KEYINPUT97), .ZN(n544) );
  AND2_X1 U497 ( .A1(n637), .A2(n366), .ZN(n543) );
  XNOR2_X2 U498 ( .A(n501), .B(n357), .ZN(n366) );
  XNOR2_X2 U499 ( .A(n430), .B(n367), .ZN(n681) );
  XNOR2_X1 U500 ( .A(n367), .B(n405), .ZN(n693) );
  XNOR2_X2 U501 ( .A(n732), .B(n433), .ZN(n367) );
  INV_X1 U502 ( .A(n625), .ZN(n414) );
  XNOR2_X1 U503 ( .A(n586), .B(KEYINPUT112), .ZN(n590) );
  NAND2_X1 U504 ( .A1(n593), .A2(n642), .ZN(n577) );
  OR2_X2 U505 ( .A1(n715), .A2(G902), .ZN(n470) );
  NAND2_X1 U506 ( .A1(n412), .A2(n409), .ZN(n408) );
  NOR2_X2 U507 ( .A1(n400), .A2(n401), .ZN(n399) );
  XNOR2_X2 U508 ( .A(n581), .B(KEYINPUT6), .ZN(n569) );
  XNOR2_X2 U509 ( .A(n474), .B(n473), .ZN(n621) );
  AND2_X2 U510 ( .A1(n621), .A2(n502), .ZN(n400) );
  NOR2_X1 U511 ( .A1(n544), .A2(n502), .ZN(n397) );
  XNOR2_X1 U512 ( .A(n680), .B(n360), .ZN(n374) );
  XNOR2_X1 U513 ( .A(n375), .B(n553), .ZN(n561) );
  NAND2_X1 U514 ( .A1(n552), .A2(n551), .ZN(n375) );
  NOR2_X1 U515 ( .A1(n589), .A2(n710), .ZN(n598) );
  NAND2_X1 U516 ( .A1(n620), .A2(n590), .ZN(n587) );
  XNOR2_X1 U517 ( .A(n694), .B(n359), .ZN(n378) );
  XNOR2_X1 U518 ( .A(n684), .B(n361), .ZN(n379) );
  XNOR2_X1 U519 ( .A(n463), .B(n462), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n713), .A2(n425), .ZN(n384) );
  NAND2_X1 U521 ( .A1(n706), .A2(n353), .ZN(n603) );
  NOR2_X1 U522 ( .A1(n580), .A2(n388), .ZN(n387) );
  XNOR2_X2 U523 ( .A(n389), .B(G143), .ZN(n476) );
  NAND2_X1 U524 ( .A1(n681), .A2(n437), .ZN(n395) );
  INV_X1 U525 ( .A(n437), .ZN(n392) );
  NAND2_X1 U526 ( .A1(n437), .A2(G902), .ZN(n394) );
  NAND2_X1 U527 ( .A1(n399), .A2(n396), .ZN(n403) );
  INV_X1 U528 ( .A(n621), .ZN(n398) );
  NAND2_X1 U529 ( .A1(n544), .A2(n502), .ZN(n402) );
  XNOR2_X2 U530 ( .A(n403), .B(n525), .ZN(n744) );
  NAND2_X1 U531 ( .A1(n404), .A2(n745), .ZN(n588) );
  XNOR2_X1 U532 ( .A(n404), .B(G131), .ZN(G33) );
  OR2_X1 U533 ( .A1(n713), .A2(n421), .ZN(n420) );
  INV_X1 U534 ( .A(n511), .ZN(n425) );
  XNOR2_X2 U535 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n427) );
  XNOR2_X1 U536 ( .A(n477), .B(n449), .ZN(n432) );
  INV_X1 U537 ( .A(n532), .ZN(n548) );
  AND2_X1 U538 ( .A1(n434), .A2(n377), .ZN(G63) );
  XNOR2_X1 U539 ( .A(n436), .B(n435), .ZN(n434) );
  XNOR2_X1 U540 ( .A(n713), .B(n362), .ZN(n435) );
  NAND2_X1 U541 ( .A1(n714), .A2(G478), .ZN(n436) );
  XNOR2_X2 U542 ( .A(KEYINPUT78), .B(n612), .ZN(n668) );
  XOR2_X1 U543 ( .A(n452), .B(n451), .Z(n437) );
  OR2_X1 U544 ( .A1(n566), .A2(n499), .ZN(n438) );
  INV_X1 U545 ( .A(KEYINPUT91), .ZN(n555) );
  INV_X1 U546 ( .A(KEYINPUT72), .ZN(n451) );
  XNOR2_X1 U547 ( .A(n468), .B(KEYINPUT25), .ZN(n469) );
  XNOR2_X1 U548 ( .A(n455), .B(n454), .ZN(n463) );
  BUF_X1 U549 ( .A(n621), .Z(n651) );
  INV_X1 U550 ( .A(KEYINPUT53), .ZN(n661) );
  NAND2_X1 U551 ( .A1(n516), .A2(G210), .ZN(n440) );
  XNOR2_X1 U552 ( .A(n440), .B(G116), .ZN(n444) );
  INV_X1 U553 ( .A(G902), .ZN(n488) );
  INV_X1 U554 ( .A(G472), .ZN(n445) );
  INV_X1 U555 ( .A(KEYINPUT98), .ZN(n447) );
  NAND2_X1 U556 ( .A1(G227), .A2(n737), .ZN(n450) );
  INV_X1 U557 ( .A(G469), .ZN(n452) );
  XNOR2_X1 U558 ( .A(n352), .B(n453), .ZN(n455) );
  NAND2_X1 U559 ( .A1(G234), .A2(n737), .ZN(n461) );
  INV_X1 U560 ( .A(KEYINPUT8), .ZN(n456) );
  NAND2_X1 U561 ( .A1(KEYINPUT70), .A2(n456), .ZN(n459) );
  INV_X1 U562 ( .A(KEYINPUT70), .ZN(n457) );
  NAND2_X1 U563 ( .A1(n457), .A2(KEYINPUT8), .ZN(n458) );
  NAND2_X1 U564 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U565 ( .A(n461), .B(n460), .ZN(n504) );
  NAND2_X1 U566 ( .A1(n504), .A2(G221), .ZN(n462) );
  XNOR2_X1 U567 ( .A(G146), .B(G125), .ZN(n475) );
  XNOR2_X1 U568 ( .A(KEYINPUT10), .B(n475), .ZN(n515) );
  XNOR2_X1 U569 ( .A(n464), .B(n515), .ZN(n734) );
  XNOR2_X1 U570 ( .A(n465), .B(n734), .ZN(n715) );
  XOR2_X1 U571 ( .A(KEYINPUT20), .B(KEYINPUT99), .Z(n467) );
  XNOR2_X1 U572 ( .A(KEYINPUT15), .B(G902), .ZN(n664) );
  NAND2_X1 U573 ( .A1(G234), .A2(n664), .ZN(n466) );
  XNOR2_X1 U574 ( .A(n467), .B(n466), .ZN(n471) );
  NAND2_X1 U575 ( .A1(n471), .A2(G217), .ZN(n468) );
  XNOR2_X2 U576 ( .A(n470), .B(n469), .ZN(n567) );
  NAND2_X1 U577 ( .A1(n471), .A2(G221), .ZN(n472) );
  XNOR2_X1 U578 ( .A(n472), .B(KEYINPUT21), .ZN(n628) );
  NAND2_X1 U579 ( .A1(n569), .A2(n541), .ZN(n474) );
  XOR2_X1 U580 ( .A(KEYINPUT110), .B(KEYINPUT33), .Z(n473) );
  XNOR2_X1 U581 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U582 ( .A(n478), .B(n477), .ZN(n483) );
  NAND2_X1 U583 ( .A1(n737), .A2(G224), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n479), .B(KEYINPUT4), .ZN(n481) );
  XNOR2_X1 U585 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n480) );
  XNOR2_X1 U586 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U587 ( .A(n483), .B(n482), .ZN(n486) );
  INV_X1 U588 ( .A(n505), .ZN(n484) );
  NAND2_X1 U589 ( .A1(n672), .A2(n664), .ZN(n492) );
  NAND2_X1 U590 ( .A1(n488), .A2(n487), .ZN(n493) );
  NAND2_X1 U591 ( .A1(n493), .A2(G210), .ZN(n490) );
  XNOR2_X1 U592 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n489) );
  XNOR2_X1 U593 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U594 ( .A1(n493), .A2(G214), .ZN(n641) );
  XOR2_X1 U595 ( .A(KEYINPUT14), .B(KEYINPUT95), .Z(n495) );
  XNOR2_X1 U596 ( .A(n495), .B(n494), .ZN(n496) );
  NAND2_X1 U597 ( .A1(G952), .A2(n496), .ZN(n657) );
  NOR2_X1 U598 ( .A1(n657), .A2(G953), .ZN(n566) );
  AND2_X1 U599 ( .A1(G902), .A2(n496), .ZN(n563) );
  NOR2_X1 U600 ( .A1(G898), .A2(n737), .ZN(n729) );
  NAND2_X1 U601 ( .A1(n563), .A2(n729), .ZN(n498) );
  INV_X1 U602 ( .A(KEYINPUT96), .ZN(n497) );
  XNOR2_X1 U603 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U604 ( .A(KEYINPUT34), .B(KEYINPUT82), .ZN(n502) );
  INV_X1 U605 ( .A(n503), .ZN(n510) );
  NAND2_X1 U606 ( .A1(G217), .A2(n504), .ZN(n508) );
  XOR2_X1 U607 ( .A(KEYINPUT7), .B(KEYINPUT107), .Z(n506) );
  XNOR2_X1 U608 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U609 ( .A(n510), .B(n509), .ZN(n713) );
  XNOR2_X1 U610 ( .A(KEYINPUT108), .B(G478), .ZN(n511) );
  XNOR2_X1 U611 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U612 ( .A(n515), .B(n514), .ZN(n522) );
  NAND2_X1 U613 ( .A1(G214), .A2(n516), .ZN(n517) );
  XNOR2_X1 U614 ( .A(n518), .B(n517), .ZN(n520) );
  NOR2_X1 U615 ( .A1(G902), .A2(n679), .ZN(n524) );
  XNOR2_X1 U616 ( .A(KEYINPUT106), .B(KEYINPUT13), .ZN(n523) );
  NOR2_X1 U617 ( .A1(n539), .A2(n538), .ZN(n592) );
  XNOR2_X1 U618 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n525) );
  INV_X1 U619 ( .A(n624), .ZN(n527) );
  INV_X1 U620 ( .A(n567), .ZN(n534) );
  INV_X1 U621 ( .A(n534), .ZN(n627) );
  NAND2_X1 U622 ( .A1(n527), .A2(n627), .ZN(n529) );
  XOR2_X1 U623 ( .A(KEYINPUT83), .B(n569), .Z(n528) );
  NOR2_X1 U624 ( .A1(n529), .A2(n528), .ZN(n533) );
  INV_X1 U625 ( .A(KEYINPUT65), .ZN(n531) );
  NOR2_X1 U626 ( .A1(n634), .A2(n534), .ZN(n535) );
  NAND2_X1 U627 ( .A1(n624), .A2(n535), .ZN(n536) );
  NOR2_X1 U628 ( .A1(n548), .A2(n536), .ZN(n686) );
  NOR2_X2 U629 ( .A1(n690), .A2(n686), .ZN(n556) );
  NAND2_X1 U630 ( .A1(n744), .A2(n556), .ZN(n537) );
  NAND2_X1 U631 ( .A1(n537), .A2(KEYINPUT44), .ZN(n552) );
  INV_X1 U632 ( .A(n538), .ZN(n540) );
  NOR2_X1 U633 ( .A1(n540), .A2(n539), .ZN(n708) );
  NOR2_X1 U634 ( .A1(n578), .A2(n708), .ZN(n646) );
  XNOR2_X1 U635 ( .A(KEYINPUT31), .B(KEYINPUT103), .ZN(n542) );
  NOR2_X1 U636 ( .A1(n544), .A2(n575), .ZN(n545) );
  NOR2_X1 U637 ( .A1(n569), .A2(n627), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n624), .A2(n546), .ZN(n547) );
  OR2_X1 U639 ( .A1(n548), .A2(n547), .ZN(n696) );
  INV_X1 U640 ( .A(n696), .ZN(n549) );
  NOR2_X1 U641 ( .A1(n550), .A2(n549), .ZN(n551) );
  INV_X1 U642 ( .A(KEYINPUT90), .ZN(n553) );
  INV_X1 U643 ( .A(KEYINPUT44), .ZN(n554) );
  AND2_X1 U644 ( .A1(n744), .A2(n554), .ZN(n558) );
  XNOR2_X1 U645 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U646 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U647 ( .A(n559), .B(KEYINPUT74), .ZN(n560) );
  NAND2_X1 U648 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X2 U649 ( .A(n562), .B(KEYINPUT45), .ZN(n719) );
  NAND2_X1 U650 ( .A1(G953), .A2(n563), .ZN(n564) );
  NOR2_X1 U651 ( .A1(G900), .A2(n564), .ZN(n565) );
  NOR2_X1 U652 ( .A1(n566), .A2(n565), .ZN(n574) );
  NOR2_X1 U653 ( .A1(n628), .A2(n574), .ZN(n568) );
  XOR2_X1 U654 ( .A(KEYINPUT111), .B(n578), .Z(n706) );
  INV_X1 U655 ( .A(n595), .ZN(n606) );
  XOR2_X1 U656 ( .A(KEYINPUT36), .B(n571), .Z(n572) );
  NOR2_X1 U657 ( .A1(n624), .A2(n572), .ZN(n710) );
  XOR2_X1 U658 ( .A(KEYINPUT38), .B(KEYINPUT75), .Z(n576) );
  XNOR2_X2 U659 ( .A(n577), .B(KEYINPUT39), .ZN(n601) );
  NAND2_X1 U660 ( .A1(n642), .A2(n641), .ZN(n647) );
  NOR2_X1 U661 ( .A1(n644), .A2(n647), .ZN(n579) );
  INV_X1 U662 ( .A(KEYINPUT28), .ZN(n583) );
  NOR2_X1 U663 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U664 ( .A(n583), .B(n582), .ZN(n584) );
  NOR2_X1 U665 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U666 ( .A(KEYINPUT42), .B(n587), .ZN(n745) );
  XNOR2_X1 U667 ( .A(n588), .B(KEYINPUT46), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n703), .A2(n429), .ZN(n591) );
  XNOR2_X1 U669 ( .A(n591), .B(KEYINPUT47), .ZN(n596) );
  AND2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n594) );
  AND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n688) );
  NOR2_X1 U672 ( .A1(n596), .A2(n688), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n600) );
  XNOR2_X2 U674 ( .A(n600), .B(n599), .ZN(n614) );
  INV_X1 U675 ( .A(n614), .ZN(n610) );
  NAND2_X1 U676 ( .A1(n601), .A2(n708), .ZN(n712) );
  NAND2_X1 U677 ( .A1(KEYINPUT2), .A2(n712), .ZN(n602) );
  XNOR2_X1 U678 ( .A(KEYINPUT85), .B(n602), .ZN(n608) );
  INV_X1 U679 ( .A(n603), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n604), .A2(n624), .ZN(n605) );
  XNOR2_X1 U681 ( .A(KEYINPUT43), .B(n605), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n689) );
  NAND2_X1 U683 ( .A1(n608), .A2(n689), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  AND2_X1 U685 ( .A1(n719), .A2(n611), .ZN(n612) );
  AND2_X1 U686 ( .A1(n712), .A2(n689), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n719), .A2(n735), .ZN(n616) );
  INV_X1 U688 ( .A(KEYINPUT2), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n666) );
  BUF_X1 U690 ( .A(n666), .Z(n617) );
  XOR2_X1 U691 ( .A(KEYINPUT86), .B(n617), .Z(n618) );
  XNOR2_X1 U692 ( .A(n619), .B(KEYINPUT88), .ZN(n623) );
  INV_X1 U693 ( .A(n620), .ZN(n640) );
  NOR2_X1 U694 ( .A1(n640), .A2(n651), .ZN(n622) );
  NOR2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n660) );
  NAND2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U697 ( .A(KEYINPUT50), .B(n626), .ZN(n632) );
  XOR2_X1 U698 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n630) );
  NAND2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U702 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U703 ( .A(KEYINPUT117), .B(n635), .Z(n636) );
  NOR2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U705 ( .A(KEYINPUT51), .B(n638), .Z(n639) );
  NOR2_X1 U706 ( .A1(n640), .A2(n639), .ZN(n653) );
  NOR2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U708 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U709 ( .A(n645), .B(KEYINPUT118), .ZN(n649) );
  NOR2_X1 U710 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U711 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U712 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U713 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U714 ( .A(n654), .B(KEYINPUT52), .Z(n655) );
  XNOR2_X1 U715 ( .A(KEYINPUT119), .B(n655), .ZN(n656) );
  NOR2_X1 U716 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U717 ( .A1(G953), .A2(n658), .ZN(n659) );
  NAND2_X1 U718 ( .A1(n660), .A2(n659), .ZN(n663) );
  XNOR2_X1 U719 ( .A(n661), .B(KEYINPUT120), .ZN(n662) );
  XNOR2_X1 U720 ( .A(n663), .B(n662), .ZN(G75) );
  INV_X1 U721 ( .A(n664), .ZN(n665) );
  NAND2_X1 U722 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X2 U723 ( .A(n667), .B(KEYINPUT64), .ZN(n669) );
  NOR2_X4 U724 ( .A1(n669), .A2(n668), .ZN(n714) );
  NAND2_X1 U725 ( .A1(n714), .A2(G210), .ZN(n674) );
  XNOR2_X1 U726 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n670) );
  XOR2_X1 U727 ( .A(n670), .B(KEYINPUT55), .Z(n671) );
  XNOR2_X1 U728 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U729 ( .A(n674), .B(n673), .ZN(n676) );
  INV_X1 U730 ( .A(G952), .ZN(n675) );
  NOR2_X2 U731 ( .A1(n676), .A2(n718), .ZN(n677) );
  XNOR2_X1 U732 ( .A(n677), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U733 ( .A1(n714), .A2(G475), .ZN(n680) );
  XOR2_X1 U734 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n678) );
  XNOR2_X1 U735 ( .A(n345), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U736 ( .A1(n714), .A2(G469), .ZN(n684) );
  XOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n683) );
  XNOR2_X1 U738 ( .A(n681), .B(KEYINPUT122), .ZN(n682) );
  INV_X1 U739 ( .A(KEYINPUT123), .ZN(n685) );
  XNOR2_X1 U740 ( .A(n347), .B(n685), .ZN(G54) );
  XOR2_X1 U741 ( .A(G110), .B(n686), .Z(G12) );
  XNOR2_X1 U742 ( .A(n688), .B(n687), .ZN(G45) );
  XNOR2_X1 U743 ( .A(n689), .B(G140), .ZN(G42) );
  XOR2_X1 U744 ( .A(n690), .B(G119), .Z(G21) );
  NAND2_X1 U745 ( .A1(n714), .A2(G472), .ZN(n694) );
  XOR2_X1 U746 ( .A(KEYINPUT92), .B(KEYINPUT114), .Z(n691) );
  XNOR2_X1 U747 ( .A(n691), .B(KEYINPUT62), .ZN(n692) );
  XNOR2_X1 U748 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n348), .B(n695), .ZN(G57) );
  XNOR2_X1 U750 ( .A(G101), .B(n696), .ZN(G3) );
  NAND2_X1 U751 ( .A1(n355), .A2(n706), .ZN(n697) );
  XNOR2_X1 U752 ( .A(n697), .B(G104), .ZN(G6) );
  XOR2_X1 U753 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n699) );
  NAND2_X1 U754 ( .A1(n355), .A2(n708), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U756 ( .A(G107), .B(n700), .ZN(G9) );
  XOR2_X1 U757 ( .A(G128), .B(KEYINPUT29), .Z(n702) );
  NAND2_X1 U758 ( .A1(n708), .A2(n703), .ZN(n701) );
  XNOR2_X1 U759 ( .A(n702), .B(n701), .ZN(G30) );
  NAND2_X1 U760 ( .A1(n703), .A2(n706), .ZN(n704) );
  XNOR2_X1 U761 ( .A(n704), .B(G146), .ZN(G48) );
  NAND2_X1 U762 ( .A1(n705), .A2(n706), .ZN(n707) );
  XNOR2_X1 U763 ( .A(n707), .B(G113), .ZN(G15) );
  NAND2_X1 U764 ( .A1(n705), .A2(n708), .ZN(n709) );
  XNOR2_X1 U765 ( .A(n709), .B(G116), .ZN(G18) );
  XNOR2_X1 U766 ( .A(G125), .B(n710), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U768 ( .A(G134), .B(n712), .ZN(G36) );
  NAND2_X1 U769 ( .A1(n714), .A2(G217), .ZN(n716) );
  XNOR2_X1 U770 ( .A(n715), .B(n716), .ZN(n717) );
  NOR2_X1 U771 ( .A1(n718), .A2(n717), .ZN(G66) );
  NAND2_X1 U772 ( .A1(n719), .A2(n737), .ZN(n723) );
  NAND2_X1 U773 ( .A1(G953), .A2(G224), .ZN(n720) );
  XNOR2_X1 U774 ( .A(KEYINPUT61), .B(n720), .ZN(n721) );
  NAND2_X1 U775 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U776 ( .A1(n723), .A2(n722), .ZN(n731) );
  XOR2_X1 U777 ( .A(n724), .B(KEYINPUT126), .Z(n725) );
  XNOR2_X1 U778 ( .A(n726), .B(n725), .ZN(n727) );
  XOR2_X1 U779 ( .A(G101), .B(n727), .Z(n728) );
  NOR2_X1 U780 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n731), .B(n730), .ZN(G69) );
  XOR2_X1 U782 ( .A(n732), .B(KEYINPUT98), .Z(n733) );
  XNOR2_X1 U783 ( .A(n734), .B(n733), .ZN(n739) );
  INV_X1 U784 ( .A(n735), .ZN(n736) );
  XNOR2_X1 U785 ( .A(n739), .B(n736), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(n737), .ZN(n743) );
  XNOR2_X1 U787 ( .A(G227), .B(n739), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U789 ( .A1(G953), .A2(n741), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n743), .A2(n742), .ZN(G72) );
  XNOR2_X1 U791 ( .A(n744), .B(G122), .ZN(G24) );
  BUF_X1 U792 ( .A(n745), .Z(n746) );
  XOR2_X1 U793 ( .A(G137), .B(n746), .Z(n747) );
  XNOR2_X1 U794 ( .A(KEYINPUT127), .B(n747), .ZN(G39) );
endmodule

