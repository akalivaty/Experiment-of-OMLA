//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n205), .A2(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT17), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT92), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(G8gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT16), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G1gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n217), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(KEYINPUT17), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n214), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n217), .B(new_n220), .ZN(new_n225));
  INV_X1    g024(.A(new_n213), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT93), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n222), .A2(new_n213), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n227), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n229), .B(KEYINPUT13), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n230), .A2(new_n231), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n228), .A2(KEYINPUT93), .A3(KEYINPUT18), .A4(new_n229), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n224), .A2(new_n229), .A3(new_n227), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n241), .A2(KEYINPUT94), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243));
  INV_X1    g042(.A(G197gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT11), .B(G169gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT12), .Z(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(new_n241), .B2(KEYINPUT94), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n236), .A2(new_n241), .A3(new_n237), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n238), .A2(new_n250), .B1(new_n251), .B2(new_n248), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT95), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n248), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n236), .A2(new_n237), .A3(new_n242), .A4(new_n249), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n255), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G226gat), .ZN(new_n260));
  INV_X1    g059(.A(G233gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT24), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n266), .B(new_n267), .C1(G183gat), .C2(G190gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n274));
  NOR2_X1   g073(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n272), .B1(KEYINPUT64), .B2(KEYINPUT23), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n268), .A2(new_n271), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT25), .B1(new_n268), .B2(KEYINPUT66), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(G190gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n284), .A2(KEYINPUT28), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(KEYINPUT28), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n273), .A2(KEYINPUT26), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n273), .A2(KEYINPUT26), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(new_n271), .A3(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n285), .A2(new_n264), .A3(new_n286), .A4(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n263), .B1(new_n280), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(G211gat), .A2(G218gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT22), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(G211gat), .A2(G218gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(G211gat), .A2(G218gat), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT73), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301));
  OR2_X1    g100(.A1(G211gat), .A2(G218gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(new_n294), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n297), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n301), .A3(new_n294), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT73), .B1(new_n298), .B2(new_n299), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n305), .A2(new_n306), .A3(new_n296), .A4(new_n293), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT29), .B1(new_n280), .B2(new_n290), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n292), .B(new_n308), .C1(new_n262), .C2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n278), .A2(new_n279), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n278), .A2(new_n279), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n290), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n262), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n311), .B1(new_n317), .B2(new_n291), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G64gat), .B(G92gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT74), .ZN(new_n321));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n318), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(KEYINPUT30), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT30), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n319), .A2(new_n328), .A3(new_n323), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G78gat), .B(G106gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT31), .B(G50gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  INV_X1    g135(.A(G155gat), .ZN(new_n337));
  INV_X1    g136(.A(G162gat), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT78), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n336), .B1(new_n339), .B2(KEYINPUT2), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(G148gat), .ZN(new_n342));
  INV_X1    g141(.A(G148gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(G141gat), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT77), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(G141gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(G148gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n336), .ZN(new_n350));
  NOR2_X1   g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT78), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n340), .A2(new_n345), .A3(new_n349), .A4(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n342), .A2(new_n344), .ZN(new_n358));
  AND2_X1   g157(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n359));
  NOR2_X1   g158(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n357), .B(new_n336), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n304), .A2(new_n316), .A3(new_n307), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT79), .B(KEYINPUT3), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n363), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n353), .A2(new_n362), .A3(new_n365), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n368), .A2(new_n316), .B1(new_n307), .B2(new_n304), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT84), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n316), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n372), .A2(new_n370), .A3(new_n308), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n335), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G22gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n308), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n377));
  INV_X1    g176(.A(new_n335), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n364), .A2(new_n363), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n374), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n375), .B1(new_n374), .B2(new_n380), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n334), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT85), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n374), .A2(new_n375), .A3(new_n380), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n385), .B1(new_n382), .B2(KEYINPUT86), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n374), .A2(new_n387), .A3(new_n375), .A4(new_n380), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n388), .A3(new_n333), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n304), .A2(new_n316), .A3(new_n307), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n390), .A2(new_n365), .B1(new_n362), .B2(new_n353), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n376), .B2(KEYINPUT84), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n369), .A2(new_n370), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n378), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n380), .ZN(new_n395));
  OAI21_X1  g194(.A(G22gat), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n385), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n334), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n389), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT87), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n384), .A2(new_n389), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G113gat), .B(G120gat), .Z(new_n407));
  INV_X1    g206(.A(KEYINPUT1), .ZN(new_n408));
  XNOR2_X1  g207(.A(G127gat), .B(G134gat), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n407), .A2(KEYINPUT68), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G127gat), .B(G134gat), .Z(new_n411));
  XNOR2_X1  g210(.A(G113gat), .B(G120gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n408), .A2(KEYINPUT68), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n280), .A2(new_n415), .A3(new_n290), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n280), .B2(new_n290), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n406), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT32), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G15gat), .B(G43gat), .Z(new_n423));
  XNOR2_X1  g222(.A(G71gat), .B(G99gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n420), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT69), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT32), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n414), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n315), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n416), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n431), .B2(new_n406), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n425), .A2(KEYINPUT33), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n405), .B1(new_n430), .B2(new_n416), .ZN(new_n435));
  INV_X1    g234(.A(new_n433), .ZN(new_n436));
  NOR4_X1   g235(.A1(new_n435), .A2(KEYINPUT69), .A3(new_n428), .A4(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n426), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT34), .B1(new_n406), .B2(KEYINPUT71), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n431), .B2(new_n406), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n430), .A2(new_n405), .A3(new_n439), .A4(new_n416), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n438), .B(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n353), .A2(new_n362), .A3(new_n410), .A4(new_n414), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT4), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n415), .A2(new_n448), .A3(new_n362), .A4(new_n353), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n377), .A2(new_n429), .A3(new_n368), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT80), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n363), .A2(new_n429), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n446), .ZN(new_n457));
  INV_X1    g256(.A(new_n451), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(KEYINPUT81), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT81), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n459), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n461), .B1(new_n453), .B2(KEYINPUT80), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G1gat), .B(G29gat), .ZN(new_n467));
  INV_X1    g266(.A(G85gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT0), .B(G57gat), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n469), .B(new_n470), .Z(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT82), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n459), .B1(new_n453), .B2(new_n461), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n368), .A2(new_n429), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n478), .A2(new_n377), .B1(new_n447), .B2(new_n449), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(new_n451), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n476), .B1(new_n480), .B2(new_n461), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n471), .B1(new_n481), .B2(new_n460), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT82), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n471), .A3(new_n460), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n475), .A2(new_n483), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n485), .A2(new_n484), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT35), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND4_X1   g287(.A1(new_n330), .A2(new_n404), .A3(new_n445), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n443), .A2(KEYINPUT70), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n438), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n490), .B(new_n426), .C1(new_n434), .C2(new_n437), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n398), .B1(new_n397), .B2(new_n334), .ZN(new_n496));
  AOI211_X1 g295(.A(KEYINPUT85), .B(new_n333), .C1(new_n396), .C2(new_n385), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n402), .B1(new_n498), .B2(new_n389), .ZN(new_n499));
  INV_X1    g298(.A(new_n403), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT91), .ZN(new_n502));
  INV_X1    g301(.A(new_n330), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n484), .B1(new_n482), .B2(KEYINPUT82), .ZN(new_n505));
  AOI211_X1 g304(.A(new_n474), .B(new_n471), .C1(new_n481), .C2(new_n460), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n475), .A2(new_n483), .A3(KEYINPUT83), .A4(new_n484), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n485), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n503), .B1(new_n509), .B2(new_n487), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n404), .A2(new_n511), .A3(new_n495), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n502), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n489), .B1(new_n513), .B2(KEYINPUT35), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n495), .A2(KEYINPUT36), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n517));
  NAND2_X1  g316(.A1(new_n444), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n510), .B2(new_n404), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n519), .B(KEYINPUT88), .C1(new_n510), .C2(new_n404), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT37), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n319), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n310), .A2(new_n318), .A3(KEYINPUT37), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n325), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n324), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT90), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n532), .A3(new_n325), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n533), .A3(new_n525), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n530), .B1(new_n534), .B2(KEYINPUT38), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(new_n487), .A3(new_n486), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n450), .A2(new_n452), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n458), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(KEYINPUT89), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(KEYINPUT89), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT39), .ZN(new_n541));
  INV_X1    g340(.A(new_n457), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(new_n451), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n539), .A2(new_n540), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n472), .B(new_n544), .C1(new_n545), .C2(KEYINPUT39), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT40), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n548), .A2(new_n503), .A3(new_n485), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n536), .A2(new_n550), .A3(new_n404), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n522), .A2(new_n523), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n259), .B1(new_n515), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT102), .ZN(new_n554));
  NAND2_X1  g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555));
  INV_X1    g354(.A(G92gat), .ZN(new_n556));
  AOI22_X1  g355(.A1(KEYINPUT8), .A2(new_n555), .B1(new_n468), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT100), .ZN(new_n558));
  XOR2_X1   g357(.A(G99gat), .B(G106gat), .Z(new_n559));
  INV_X1    g358(.A(KEYINPUT101), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT7), .B1(new_n468), .B2(new_n556), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(G85gat), .A3(G92gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n559), .A2(new_n560), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n558), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n562), .B1(new_n558), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n554), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n558), .A2(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n561), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(KEYINPUT102), .A3(new_n567), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n213), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT41), .ZN(new_n575));
  INV_X1    g374(.A(G232gat), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n575), .A2(new_n576), .A3(new_n261), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT103), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n568), .A2(new_n554), .A3(new_n569), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT102), .B1(new_n572), .B2(new_n567), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n226), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT103), .ZN(new_n582));
  INV_X1    g381(.A(new_n577), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n579), .A2(new_n580), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(new_n214), .A3(new_n223), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G190gat), .B(G218gat), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n589), .A3(new_n587), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT104), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(new_n597), .A3(new_n592), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n585), .A2(KEYINPUT104), .A3(new_n587), .A4(new_n589), .ZN(new_n599));
  INV_X1    g398(.A(new_n595), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(new_n601), .A3(KEYINPUT105), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT105), .B1(new_n598), .B2(new_n601), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n596), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n606));
  INV_X1    g405(.A(G57gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G64gat), .ZN(new_n608));
  INV_X1    g407(.A(G64gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(G57gat), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT97), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G71gat), .B(G78gat), .Z(new_n614));
  OR2_X1    g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n611), .A2(KEYINPUT97), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n616), .B1(new_n613), .B2(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n618), .A2(KEYINPUT98), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(KEYINPUT98), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(KEYINPUT21), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n618), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n622), .A2(KEYINPUT21), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n225), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n623), .A2(new_n225), .ZN(new_n625));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT99), .ZN(new_n627));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR3_X1    g428(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n629), .B1(new_n624), .B2(new_n625), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n630), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n630), .B2(new_n634), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT106), .B1(new_n605), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n596), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n598), .A2(new_n601), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n640), .B1(new_n643), .B2(new_n602), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT106), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n637), .ZN(new_n646));
  INV_X1    g445(.A(G230gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n261), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n619), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(new_n586), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n622), .B1(new_n572), .B2(new_n567), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n618), .A2(new_n568), .A3(new_n569), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n648), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n648), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n655), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n655), .B2(new_n657), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n639), .A2(new_n646), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n553), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n509), .A2(new_n487), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n503), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT16), .B(G8gat), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT107), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n677), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n673), .A2(new_n672), .A3(new_n674), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n673), .A2(G8gat), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n676), .A2(new_n678), .A3(new_n679), .A4(new_n680), .ZN(G1325gat));
  AOI21_X1  g480(.A(G15gat), .B1(new_n667), .B2(new_n445), .ZN(new_n682));
  INV_X1    g481(.A(new_n519), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(G15gat), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n682), .B1(new_n667), .B2(new_n684), .ZN(G1326gat));
  INV_X1    g484(.A(new_n404), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n667), .A2(new_n375), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n553), .A2(new_n686), .A3(new_n666), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G22gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n690), .B(new_n692), .ZN(G1327gat));
  NOR3_X1   g492(.A1(new_n644), .A2(new_n637), .A3(new_n663), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n553), .A2(new_n203), .A3(new_n669), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n551), .B(new_n519), .C1(new_n510), .C2(new_n404), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n605), .B1(new_n514), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n644), .A2(new_n700), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n522), .A2(new_n523), .A3(new_n551), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n703), .B2(new_n514), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n255), .A2(new_n256), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n638), .A3(new_n664), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT109), .Z(new_n707));
  NAND3_X1  g506(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n668), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n696), .A2(new_n709), .ZN(G1328gat));
  NAND4_X1  g509(.A1(new_n553), .A2(new_n204), .A3(new_n503), .A4(new_n694), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n708), .B2(new_n330), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(G1329gat));
  NAND4_X1  g514(.A1(new_n701), .A2(new_n704), .A3(new_n683), .A4(new_n707), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G43gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n444), .A2(G43gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n553), .A2(new_n694), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1330gat));
  OAI21_X1  g521(.A(G50gat), .B1(new_n708), .B2(new_n404), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT111), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n404), .A2(G50gat), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT110), .Z(new_n726));
  NAND3_X1  g525(.A1(new_n553), .A2(new_n694), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n724), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n723), .B(new_n727), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  INV_X1    g531(.A(KEYINPUT35), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n511), .B1(new_n404), .B2(new_n495), .ZN(new_n734));
  AOI211_X1 g533(.A(KEYINPUT91), .B(new_n494), .C1(new_n401), .C2(new_n403), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n736), .B2(new_n510), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n697), .B1(new_n737), .B2(new_n489), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n705), .A2(new_n664), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n639), .A2(new_n646), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n639), .A2(new_n646), .A3(KEYINPUT112), .A4(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n738), .A2(new_n744), .A3(new_n669), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g545(.A1(new_n738), .A2(new_n744), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT113), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n738), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n330), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n756));
  INV_X1    g555(.A(new_n750), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n749), .B1(new_n738), .B2(new_n744), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n683), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G71gat), .ZN(new_n760));
  INV_X1    g559(.A(G71gat), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n738), .A2(new_n744), .A3(new_n761), .A4(new_n445), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n756), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n519), .B1(new_n748), .B2(new_n750), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n756), .B(new_n762), .C1(new_n764), .C2(new_n761), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n763), .A2(new_n766), .ZN(G1334gat));
  OAI21_X1  g566(.A(new_n686), .B1(new_n757), .B2(new_n758), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g568(.A1(new_n252), .A2(new_n638), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n664), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT114), .ZN(new_n772));
  AND4_X1   g571(.A1(new_n669), .A2(new_n701), .A3(new_n704), .A4(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n770), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n605), .B(new_n774), .C1(new_n514), .C2(new_n698), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT51), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n738), .A2(new_n777), .A3(new_n605), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n669), .A2(new_n468), .A3(new_n663), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n773), .A2(new_n468), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  AOI22_X1  g580(.A1(new_n776), .A2(new_n778), .B1(KEYINPUT115), .B2(new_n775), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n775), .A2(KEYINPUT115), .A3(new_n777), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n663), .A2(new_n503), .A3(new_n556), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n701), .A2(new_n704), .A3(new_n503), .A4(new_n772), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(G92gat), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT52), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n779), .B2(new_n784), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(G1337gat));
  NAND4_X1  g591(.A1(new_n701), .A2(new_n704), .A3(new_n683), .A4(new_n772), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G99gat), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n664), .A2(new_n444), .A3(G99gat), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n795), .A2(new_n796), .B1(new_n779), .B2(new_n797), .ZN(G1338gat));
  NOR3_X1   g597(.A1(new_n404), .A2(new_n664), .A3(G106gat), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT117), .Z(new_n800));
  NOR3_X1   g599(.A1(new_n782), .A2(new_n783), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n701), .A2(new_n704), .A3(new_n686), .A4(new_n772), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(G106gat), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT53), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n776), .A2(new_n778), .A3(new_n799), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT118), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n802), .A2(G106gat), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n806), .A4(new_n805), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n804), .A2(new_n808), .A3(new_n811), .ZN(G1339gat));
  NAND2_X1  g611(.A1(new_n650), .A2(new_n654), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n656), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n650), .A2(new_n648), .A3(new_n654), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n660), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n655), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT119), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n819), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n661), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n820), .A2(new_n826), .A3(new_n821), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n705), .A2(new_n823), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n232), .A2(new_n227), .A3(new_n234), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT120), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n228), .A2(new_n229), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n247), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(KEYINPUT121), .B(new_n247), .C1(new_n830), .C2(new_n831), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n663), .A3(new_n256), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n605), .B1(new_n828), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n825), .A3(new_n827), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n256), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n839), .A2(new_n644), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n638), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n639), .A2(new_n646), .A3(new_n252), .A4(new_n664), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n668), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n736), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n503), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n705), .ZN(new_n847));
  INV_X1    g646(.A(G113gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n686), .A2(new_n444), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n503), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n844), .A2(G113gat), .A3(new_n258), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n849), .A2(KEYINPUT122), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1340gat));
  INV_X1    g657(.A(G120gat), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n846), .A2(new_n859), .A3(new_n663), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n852), .ZN(new_n861));
  OAI21_X1  g660(.A(G120gat), .B1(new_n861), .B2(new_n664), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n861), .A2(new_n864), .A3(new_n638), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n637), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n864), .ZN(G1342gat));
  NAND2_X1  g666(.A1(new_n605), .A2(new_n330), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT123), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n845), .A2(G134gat), .A3(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n861), .B2(new_n644), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(G1343gat));
  INV_X1    g673(.A(new_n841), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n828), .A2(new_n837), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n644), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n637), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n843), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n686), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n683), .A2(new_n668), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n330), .ZN(new_n882));
  NOR4_X1   g681(.A1(new_n880), .A2(G141gat), .A3(new_n259), .A4(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n825), .A2(new_n822), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n254), .A2(new_n257), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n837), .B(KEYINPUT124), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n644), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n637), .B1(new_n889), .B2(new_n875), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT57), .B(new_n686), .C1(new_n890), .C2(new_n879), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n882), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n705), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n883), .B1(new_n893), .B2(G141gat), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n341), .B1(new_n892), .B2(new_n258), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n883), .A2(KEYINPUT58), .ZN(new_n897));
  OAI22_X1  g696(.A1(new_n894), .A2(new_n895), .B1(new_n896), .B2(new_n897), .ZN(G1344gat));
  NOR2_X1   g697(.A1(new_n880), .A2(new_n882), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n343), .A3(new_n663), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT59), .B(new_n343), .C1(new_n892), .C2(new_n663), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n665), .A2(new_n258), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n884), .B(new_n686), .C1(new_n890), .C2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n882), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n903), .A2(new_n905), .A3(new_n663), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n902), .B1(new_n907), .B2(G148gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n900), .B1(new_n901), .B2(new_n908), .ZN(G1345gat));
  AOI21_X1  g708(.A(G155gat), .B1(new_n899), .B2(new_n637), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n638), .A2(new_n337), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n892), .B2(new_n911), .ZN(G1346gat));
  AND2_X1   g711(.A1(new_n892), .A2(new_n605), .ZN(new_n913));
  INV_X1    g712(.A(new_n869), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n338), .A3(new_n881), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n913), .A2(new_n338), .B1(new_n880), .B2(new_n915), .ZN(G1347gat));
  AOI21_X1  g715(.A(new_n669), .B1(new_n842), .B2(new_n843), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n851), .A2(new_n330), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n259), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n668), .B1(new_n878), .B2(new_n879), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT125), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n503), .A3(new_n736), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n252), .A2(G169gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n920), .B1(new_n926), .B2(new_n927), .ZN(G1348gat));
  INV_X1    g727(.A(G176gat), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n919), .A2(new_n929), .A3(new_n664), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n330), .B1(new_n922), .B2(new_n924), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n736), .A3(new_n663), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n932), .B2(new_n929), .ZN(G1349gat));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n637), .A3(new_n918), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(G183gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n637), .A2(new_n282), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n926), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT60), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n936), .B(new_n940), .C1(new_n926), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n919), .B2(new_n644), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n605), .A2(new_n283), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n944), .A2(new_n945), .B1(new_n926), .B2(new_n946), .ZN(G1351gat));
  NOR3_X1   g746(.A1(new_n683), .A2(new_n669), .A3(new_n330), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n903), .A2(new_n905), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n259), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n683), .A2(new_n404), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n917), .A2(new_n923), .ZN(new_n952));
  AOI211_X1 g751(.A(KEYINPUT125), .B(new_n669), .C1(new_n842), .C2(new_n843), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n503), .B(new_n951), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n705), .A2(new_n244), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(G1352gat));
  NOR2_X1   g755(.A1(new_n664), .A2(G204gat), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n903), .A2(new_n905), .A3(new_n663), .A4(new_n948), .ZN(new_n961));
  AOI22_X1  g760(.A1(new_n959), .A2(new_n960), .B1(G204gat), .B2(new_n961), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n925), .A2(new_n503), .A3(new_n951), .A4(new_n957), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT127), .B1(new_n963), .B2(KEYINPUT62), .ZN(new_n964));
  OAI211_X1 g763(.A(KEYINPUT127), .B(KEYINPUT62), .C1(new_n954), .C2(new_n958), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n964), .B2(new_n966), .ZN(G1353gat));
  OR3_X1    g766(.A1(new_n954), .A2(G211gat), .A3(new_n638), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n903), .A2(new_n905), .A3(new_n637), .A4(new_n948), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  INV_X1    g772(.A(G218gat), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n949), .A2(new_n974), .A3(new_n644), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n931), .A2(new_n605), .A3(new_n951), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n974), .B2(new_n976), .ZN(G1355gat));
endmodule


