//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(KEYINPUT24), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(G169gat), .A3(G176gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n208), .A2(new_n210), .B1(KEYINPUT23), .B2(new_n202), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT24), .A3(new_n204), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n206), .A2(new_n211), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n206), .A2(new_n211), .A3(KEYINPUT25), .A4(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n202), .B(KEYINPUT26), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n208), .A2(new_n210), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n221), .A2(new_n222), .B1(G183gat), .B2(G190gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT27), .B(G183gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n213), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n213), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n224), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n223), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n220), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT70), .ZN(new_n232));
  NAND2_X1  g031(.A1(G226gat), .A2(G233gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n227), .A2(new_n229), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n223), .A2(new_n236), .B1(new_n218), .B2(new_n219), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT70), .B1(new_n237), .B2(new_n233), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n234), .B1(new_n231), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n235), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G211gat), .B(G218gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g042(.A(G197gat), .B(G204gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(G211gat), .A2(G218gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT22), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n246), .B1(new_n245), .B2(new_n247), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n243), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(KEYINPUT68), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(KEYINPUT68), .B(new_n242), .C1(new_n249), .C2(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT69), .B(KEYINPUT29), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n233), .B1(new_n237), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n231), .A2(new_n234), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n256), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(G64gat), .B(G92gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  NAND3_X1  g065(.A1(new_n257), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT30), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n257), .A2(new_n263), .ZN(new_n272));
  INV_X1    g071(.A(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n269), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(KEYINPUT82), .B(KEYINPUT0), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT83), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G57gat), .B(G85gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(KEYINPUT81), .ZN(new_n282));
  NAND2_X1  g081(.A1(G225gat), .A2(G233gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT76), .B(G162gat), .ZN(new_n289));
  INV_X1    g088(.A(G155gat), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT2), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G141gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT73), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G141gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .A4(G148gat), .ZN(new_n297));
  OR2_X1    g096(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(G141gat), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(G141gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n296), .B1(new_n302), .B2(G148gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n288), .B(new_n291), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G148gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G141gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n292), .A2(G148gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n306), .A2(new_n307), .B1(new_n308), .B2(KEYINPUT2), .ZN(new_n309));
  INV_X1    g108(.A(new_n286), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n284), .A2(KEYINPUT72), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n308), .A2(G155gat), .A3(G162gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n304), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G127gat), .B(G134gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G113gat), .A2(G120gat), .ZN(new_n318));
  INV_X1    g117(.A(G113gat), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT1), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G134gat), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n323), .A2(G127gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(G127gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(G113gat), .B2(G120gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n318), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n324), .A2(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n322), .A2(new_n329), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n301), .A2(new_n303), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n291), .A2(new_n288), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n315), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n283), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n282), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n283), .ZN(new_n339));
  INV_X1    g138(.A(new_n335), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n332), .B1(new_n304), .B2(new_n315), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n337), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(KEYINPUT81), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n332), .B1(new_n316), .B2(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n293), .A2(new_n295), .A3(G148gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT74), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n297), .A3(new_n300), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G162gat), .ZN(new_n350));
  INV_X1    g149(.A(G162gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT76), .ZN(new_n352));
  OAI21_X1  g151(.A(G155gat), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n287), .B1(new_n353), .B2(KEYINPUT2), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n314), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(new_n355), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n345), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n283), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n362));
  AOI211_X1 g161(.A(KEYINPUT79), .B(new_n362), .C1(new_n355), .C2(new_n332), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n364));
  INV_X1    g163(.A(new_n362), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n335), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n335), .A2(KEYINPUT4), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n363), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n338), .B(new_n344), .C1(new_n361), .C2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n335), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n335), .B2(new_n362), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n373), .A2(new_n360), .A3(new_n283), .A4(new_n337), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n281), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n331), .A2(new_n335), .A3(new_n283), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT39), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n360), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(new_n339), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT39), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n330), .B1(new_n355), .B2(new_n357), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT77), .B1(new_n316), .B2(KEYINPUT3), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n380), .B(new_n339), .C1(new_n384), .C2(new_n372), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n281), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n375), .B1(KEYINPUT40), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT40), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n389), .B1(new_n379), .B2(new_n386), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT87), .B(new_n389), .C1(new_n379), .C2(new_n386), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n275), .A2(new_n388), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n382), .A2(new_n383), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n256), .B1(new_n395), .B2(new_n258), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n253), .A2(new_n239), .A3(new_n254), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n355), .B1(new_n397), .B2(new_n357), .ZN(new_n398));
  OAI211_X1 g197(.A(G228gat), .B(G233gat), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G228gat), .A2(G233gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n357), .B1(new_n255), .B2(new_n259), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n316), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n259), .B1(new_n382), .B2(new_n383), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n400), .B(new_n402), .C1(new_n403), .C2(new_n256), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G50gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G22gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n258), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n398), .B1(new_n411), .B2(new_n255), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n404), .B(new_n410), .C1(new_n412), .C2(new_n400), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n409), .ZN(new_n415));
  INV_X1    g214(.A(new_n413), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n410), .B1(new_n399), .B2(new_n404), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n262), .B1(new_n241), .B2(new_n256), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n266), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n241), .A2(new_n255), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n260), .A2(new_n261), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n425), .B2(new_n256), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT38), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n420), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n273), .B1(new_n272), .B2(KEYINPUT37), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n421), .A2(new_n422), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT38), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n423), .A2(new_n420), .A3(new_n427), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n429), .A2(new_n432), .A3(new_n267), .A4(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n369), .A2(new_n374), .A3(new_n281), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT84), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n369), .A2(new_n374), .ZN(new_n437));
  INV_X1    g236(.A(new_n281), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n369), .A2(new_n441), .A3(new_n374), .A4(new_n281), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n436), .A2(new_n439), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n375), .A2(new_n444), .A3(KEYINPUT6), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT86), .B1(new_n439), .B2(new_n440), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n394), .B(new_n419), .C1(new_n434), .C2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT36), .ZN(new_n449));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n220), .A2(new_n332), .A3(new_n230), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n332), .B1(new_n220), .B2(new_n230), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT32), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(G15gat), .B(G43gat), .Z(new_n458));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n460), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n454), .B(KEYINPUT32), .C1(new_n456), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n452), .A2(new_n453), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT66), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n464), .A2(new_n450), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n461), .B2(new_n463), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n465), .A2(new_n466), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n461), .A2(new_n463), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n467), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n476), .B2(new_n469), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n449), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n473), .B1(new_n470), .B2(new_n471), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n472), .A3(new_n469), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT36), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT85), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n337), .A2(new_n283), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n384), .A2(new_n372), .A3(new_n485), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n336), .A2(new_n282), .A3(new_n337), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT81), .B1(new_n342), .B2(new_n343), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n366), .A2(new_n367), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n360), .B(new_n283), .C1(new_n490), .C2(new_n363), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n486), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n441), .B1(new_n492), .B2(new_n281), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n442), .A2(new_n440), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n484), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n436), .A2(KEYINPUT85), .A3(new_n440), .A4(new_n442), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n439), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n446), .A2(new_n445), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n275), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n448), .B(new_n483), .C1(new_n499), .C2(new_n419), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT35), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n414), .A2(new_n418), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n480), .B2(new_n479), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n275), .ZN(new_n505));
  AND4_X1   g304(.A1(new_n501), .A2(new_n503), .A3(new_n505), .A4(new_n447), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n500), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(G197gat), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT11), .B(G169gat), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT12), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  OR2_X1    g313(.A1(G43gat), .A2(G50gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(G43gat), .A2(G50gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT15), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT14), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT14), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n524), .A2(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n521), .A2(new_n523), .A3(KEYINPUT89), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n518), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n515), .A2(new_n529), .A3(new_n516), .ZN(new_n530));
  NAND2_X1  g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n532), .A2(new_n518), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n524), .A2(KEYINPUT90), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n521), .A2(new_n523), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n528), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(G1gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G1gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT16), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n539), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n545), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n547), .A2(new_n541), .A3(G8gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT92), .B1(new_n538), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n532), .A2(new_n536), .A3(new_n518), .A4(new_n534), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n551), .B(KEYINPUT17), .C1(new_n553), .C2(new_n528), .ZN(new_n554));
  INV_X1    g353(.A(new_n528), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n555), .A2(new_n552), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n550), .B1(new_n559), .B2(new_n549), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n546), .A2(new_n548), .ZN(new_n561));
  AOI211_X1 g360(.A(KEYINPUT92), .B(new_n561), .C1(new_n554), .C2(new_n558), .ZN(new_n562));
  OAI211_X1 g361(.A(KEYINPUT18), .B(new_n514), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n538), .B(new_n549), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(new_n514), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n559), .A2(new_n569), .A3(new_n549), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n561), .B1(new_n554), .B2(new_n558), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(new_n550), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT18), .B1(new_n572), .B2(new_n514), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n513), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n514), .B1(new_n560), .B2(new_n562), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT18), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n577), .A2(new_n512), .A3(new_n563), .A4(new_n567), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(KEYINPUT94), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n580), .B(new_n513), .C1(new_n568), .C2(new_n573), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n507), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT98), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(G85gat), .A3(G92gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n589), .A3(KEYINPUT7), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(KEYINPUT99), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n586), .A2(KEYINPUT7), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT100), .B(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n594), .A2(new_n595), .B1(KEYINPUT8), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n591), .A2(new_n599), .A3(new_n593), .A4(new_n597), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n554), .B2(new_n558), .ZN(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n602), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(new_n538), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n585), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n559), .A2(new_n607), .ZN(new_n612));
  INV_X1    g411(.A(new_n585), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n607), .A2(new_n538), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .A4(new_n606), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n616));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n609), .A2(new_n610), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n611), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n609), .A2(new_n615), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n624), .B2(new_n618), .ZN(new_n625));
  AOI211_X1 g424(.A(KEYINPUT101), .B(new_n619), .C1(new_n609), .C2(new_n615), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(G71gat), .A2(G78gat), .ZN(new_n630));
  XOR2_X1   g429(.A(G57gat), .B(G64gat), .Z(new_n631));
  AOI211_X1 g430(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(KEYINPUT9), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n629), .B1(KEYINPUT9), .B2(new_n630), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT95), .B(G57gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(G64gat), .ZN(new_n635));
  INV_X1    g434(.A(G64gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(G57gat), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n633), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(KEYINPUT21), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n561), .B1(KEYINPUT21), .B2(new_n639), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G127gat), .B(G155gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT20), .ZN(new_n646));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(KEYINPUT96), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n644), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n628), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(G230gat), .ZN(new_n655));
  INV_X1    g454(.A(G233gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n639), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n607), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n601), .A2(new_n639), .A3(new_n602), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n601), .A2(new_n639), .A3(new_n602), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT10), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n657), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n657), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n659), .B2(new_n661), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT103), .ZN(new_n670));
  XOR2_X1   g469(.A(G176gat), .B(G204gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n668), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n654), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n584), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n446), .A2(new_n445), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n436), .A2(new_n440), .A3(new_n442), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n375), .B1(new_n678), .B2(new_n484), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n679), .B2(new_n496), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  NAND4_X1  g481(.A1(new_n507), .A2(new_n275), .A3(new_n583), .A4(new_n674), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n683), .B2(new_n685), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT104), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n683), .A2(G8gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(G1325gat));
  INV_X1    g491(.A(new_n676), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n693), .B2(new_n483), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n479), .A2(new_n480), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(G15gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n694), .B1(new_n693), .B2(new_n697), .ZN(G1326gat));
  NAND2_X1  g497(.A1(new_n676), .A2(new_n502), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n497), .A2(new_n498), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n505), .A3(new_n503), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT35), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n419), .A2(new_n695), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n275), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n501), .A3(new_n447), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n502), .B1(new_n680), .B2(new_n275), .ZN(new_n709));
  INV_X1    g508(.A(new_n433), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n428), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n423), .B1(new_n422), .B2(new_n421), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n712), .A2(KEYINPUT38), .B1(new_n421), .B2(new_n266), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n498), .A2(new_n443), .A3(new_n711), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n387), .A2(KEYINPUT40), .ZN(new_n715));
  AND4_X1   g514(.A1(new_n439), .A2(new_n392), .A3(new_n393), .A4(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n502), .B1(new_n716), .B2(new_n275), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n482), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n705), .A2(new_n708), .B1(new_n709), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n702), .B1(new_n719), .B2(new_n628), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n507), .A2(KEYINPUT44), .A3(new_n627), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n673), .B(KEYINPUT107), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n724), .A2(new_n583), .A3(new_n652), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT108), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n703), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n628), .A2(new_n653), .A3(new_n673), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT106), .Z(new_n730));
  AND3_X1   g529(.A1(new_n507), .A2(new_n583), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n519), .A3(new_n680), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n733), .ZN(G1328gat));
  OAI21_X1  g533(.A(G36gat), .B1(new_n727), .B2(new_n505), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(new_n520), .A3(new_n275), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(G1329gat));
  NAND4_X1  g538(.A1(new_n720), .A2(new_n482), .A3(new_n721), .A4(new_n726), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G43gat), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n696), .A2(G43gat), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n507), .A2(new_n583), .A3(new_n730), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(KEYINPUT47), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n719), .A2(new_n582), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n745), .A2(KEYINPUT109), .A3(new_n730), .A4(new_n742), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(G43gat), .B2(new_n740), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n744), .B1(new_n750), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g550(.A1(new_n720), .A2(new_n502), .A3(new_n721), .A4(new_n726), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G50gat), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n419), .A2(G50gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n507), .A2(new_n583), .A3(new_n730), .A4(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(KEYINPUT48), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n745), .A2(new_n757), .A3(new_n730), .A4(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(KEYINPUT110), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(G50gat), .B2(new_n752), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n756), .B1(new_n761), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g561(.A1(new_n724), .A2(new_n583), .A3(new_n654), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT111), .Z(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n719), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n680), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(new_n634), .Z(G1332gat));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n505), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n768), .B1(new_n765), .B2(new_n769), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n771), .A2(new_n772), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n772), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n775), .A3(new_n770), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(G1333gat));
  INV_X1    g576(.A(G71gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n765), .B2(new_n482), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n764), .A2(new_n719), .A3(G71gat), .A4(new_n696), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n502), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n507), .A2(new_n627), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n583), .A2(new_n653), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n705), .A2(new_n708), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n628), .B1(new_n792), .B2(new_n500), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(KEYINPUT51), .A3(new_n789), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n791), .A2(new_n794), .A3(KEYINPUT113), .ZN(new_n798));
  INV_X1    g597(.A(new_n594), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n703), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n797), .A2(new_n673), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n789), .A2(new_n673), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n722), .A2(new_n680), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n799), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1336gat));
  NAND4_X1  g604(.A1(new_n720), .A2(new_n275), .A3(new_n721), .A4(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G92gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n724), .A2(G92gat), .A3(new_n505), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n793), .B2(new_n789), .ZN(new_n809));
  AND4_X1   g608(.A1(KEYINPUT51), .A2(new_n507), .A3(new_n627), .A4(new_n789), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n807), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(G1337gat));
  NOR2_X1   g615(.A1(new_n696), .A2(G99gat), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n797), .A2(new_n673), .A3(new_n798), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n722), .A2(new_n482), .A3(new_n802), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G99gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1338gat));
  NAND4_X1  g620(.A1(new_n720), .A2(new_n502), .A3(new_n721), .A4(new_n802), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G106gat), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n724), .A2(G106gat), .A3(new_n419), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n809), .B2(new_n810), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n824), .B(KEYINPUT114), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n795), .A2(new_n828), .B1(new_n822), .B2(G106gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n829), .B2(new_n826), .ZN(G1339gat));
  NAND2_X1  g629(.A1(new_n674), .A2(new_n582), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n572), .B2(new_n514), .ZN(new_n833));
  INV_X1    g632(.A(new_n560), .ZN(new_n834));
  INV_X1    g633(.A(new_n514), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n834), .A2(KEYINPUT116), .A3(new_n835), .A4(new_n570), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n833), .B(new_n836), .C1(new_n564), .C2(new_n566), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n511), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n627), .A2(new_n838), .A3(new_n578), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n639), .B1(new_n601), .B2(new_n602), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n663), .A2(new_n841), .A3(KEYINPUT10), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n661), .A2(new_n660), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n666), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n662), .A2(new_n664), .A3(new_n657), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n844), .A2(KEYINPUT115), .A3(KEYINPUT54), .A4(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n672), .B1(new_n665), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n662), .A2(new_n664), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n847), .B1(new_n850), .B2(new_n666), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT115), .B1(new_n851), .B2(new_n845), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n840), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n668), .A2(new_n672), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n844), .A2(KEYINPUT54), .A3(new_n845), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n857), .A2(KEYINPUT55), .A3(new_n846), .A4(new_n848), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n853), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n839), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n838), .A2(new_n578), .A3(new_n673), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n582), .B2(new_n859), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n862), .B2(new_n628), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n831), .B1(new_n863), .B2(new_n653), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n680), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n707), .ZN(new_n866));
  OAI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n582), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n582), .A2(G113gat), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT117), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n866), .B2(new_n869), .ZN(G1340gat));
  NOR3_X1   g669(.A1(new_n866), .A2(new_n320), .A3(new_n724), .ZN(new_n871));
  INV_X1    g670(.A(new_n866), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n673), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n320), .B2(new_n873), .ZN(G1341gat));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n653), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(G127gat), .ZN(G1342gat));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n866), .A2(new_n628), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n879), .B2(G134gat), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n878), .A2(KEYINPUT118), .A3(new_n323), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n878), .A2(KEYINPUT56), .A3(new_n323), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT56), .B1(new_n878), .B2(new_n323), .ZN(new_n883));
  OAI22_X1  g682(.A1(new_n880), .A2(new_n881), .B1(new_n882), .B2(new_n883), .ZN(G1343gat));
  NOR3_X1   g683(.A1(new_n703), .A2(new_n482), .A3(new_n275), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT119), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n864), .A2(new_n502), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n864), .A2(KEYINPUT57), .A3(new_n502), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n302), .B1(new_n891), .B2(new_n583), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n482), .A2(new_n419), .ZN(new_n893));
  AND4_X1   g692(.A1(new_n680), .A2(new_n864), .A3(new_n505), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n583), .A2(new_n292), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT120), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT58), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n885), .B(KEYINPUT119), .Z(new_n899));
  AND3_X1   g698(.A1(new_n864), .A2(KEYINPUT57), .A3(new_n502), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n864), .B2(new_n502), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n899), .B(new_n583), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT121), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n889), .A2(new_n890), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n583), .A4(new_n899), .ZN(new_n906));
  INV_X1    g705(.A(new_n302), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n897), .A2(KEYINPUT58), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n898), .B1(new_n908), .B2(new_n909), .ZN(G1344gat));
  AND2_X1   g709(.A1(new_n298), .A2(new_n299), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n911), .A3(new_n673), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n891), .A2(new_n673), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT59), .B(new_n911), .C1(new_n891), .C2(new_n673), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(G1345gat));
  AOI21_X1  g716(.A(new_n290), .B1(new_n891), .B2(new_n653), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n894), .A2(new_n290), .A3(new_n653), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n919), .ZN(G1346gat));
  NOR2_X1   g719(.A1(new_n628), .A2(new_n289), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n894), .A2(new_n627), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n891), .A2(new_n921), .B1(new_n922), .B2(new_n289), .ZN(G1347gat));
  AND2_X1   g722(.A1(new_n864), .A2(new_n703), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n706), .A2(new_n505), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(G169gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n929), .A3(new_n583), .ZN(new_n930));
  INV_X1    g729(.A(new_n926), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT123), .B(new_n929), .C1(new_n931), .C2(new_n583), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n583), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(G169gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n930), .B1(new_n932), .B2(new_n935), .ZN(G1348gat));
  AOI21_X1  g735(.A(G176gat), .B1(new_n928), .B2(new_n673), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n924), .A2(G176gat), .A3(new_n723), .A4(new_n925), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT124), .Z(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(G1349gat));
  NAND4_X1  g739(.A1(new_n864), .A2(new_n703), .A3(new_n653), .A4(new_n925), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n212), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(new_n226), .B2(new_n941), .ZN(new_n943));
  XNOR2_X1  g742(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n943), .A2(KEYINPUT126), .A3(new_n944), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n947), .B(new_n948), .C1(new_n949), .C2(new_n943), .ZN(G1350gat));
  NAND3_X1  g749(.A1(new_n928), .A2(new_n213), .A3(new_n627), .ZN(new_n951));
  AOI211_X1 g750(.A(KEYINPUT61), .B(new_n213), .C1(new_n931), .C2(new_n627), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n931), .A2(new_n627), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(G190gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n952), .B2(new_n955), .ZN(G1351gat));
  NAND2_X1  g755(.A1(new_n893), .A2(new_n275), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT127), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n924), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n583), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n680), .A2(new_n482), .A3(new_n505), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n904), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n583), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  INV_X1    g764(.A(G204gat), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n924), .A2(new_n958), .A3(new_n966), .A4(new_n673), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT62), .Z(new_n968));
  NAND3_X1  g767(.A1(new_n904), .A2(new_n723), .A3(new_n962), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n966), .B2(new_n970), .ZN(G1353gat));
  OR3_X1    g770(.A1(new_n959), .A2(G211gat), .A3(new_n652), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n904), .A2(new_n653), .A3(new_n962), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  INV_X1    g775(.A(G218gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n977), .A3(new_n627), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n627), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n978), .B1(new_n980), .B2(new_n977), .ZN(G1355gat));
endmodule


