

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749;

  XOR2_X1 U373 ( .A(n549), .B(n518), .Z(n614) );
  INV_X1 U374 ( .A(G953), .ZN(n736) );
  XNOR2_X1 U375 ( .A(n534), .B(KEYINPUT40), .ZN(n748) );
  AND2_X2 U376 ( .A1(n587), .A2(n397), .ZN(n432) );
  XNOR2_X2 U377 ( .A(n438), .B(n437), .ZN(n448) );
  XOR2_X2 U378 ( .A(G104), .B(G107), .Z(n438) );
  NAND2_X2 U379 ( .A1(n395), .A2(n391), .ZN(n403) );
  NOR2_X1 U380 ( .A1(n749), .A2(n748), .ZN(n535) );
  XNOR2_X1 U381 ( .A(n451), .B(G469), .ZN(n527) );
  XNOR2_X1 U382 ( .A(n526), .B(KEYINPUT42), .ZN(n749) );
  AND2_X1 U383 ( .A1(n533), .A2(n409), .ZN(n548) );
  NOR2_X1 U384 ( .A1(n527), .A2(n524), .ZN(n525) );
  BUF_X1 U385 ( .A(n537), .Z(n549) );
  OR2_X1 U386 ( .A1(n609), .A2(G902), .ZN(n495) );
  XNOR2_X1 U387 ( .A(n416), .B(n734), .ZN(n609) );
  XNOR2_X1 U388 ( .A(n733), .B(G146), .ZN(n508) );
  XNOR2_X1 U389 ( .A(n448), .B(n425), .ZN(n718) );
  XOR2_X1 U390 ( .A(G137), .B(G140), .Z(n484) );
  INV_X2 U391 ( .A(G143), .ZN(n440) );
  OR2_X2 U392 ( .A1(n666), .A2(G902), .ZN(n385) );
  XNOR2_X2 U393 ( .A(n431), .B(n358), .ZN(n537) );
  XNOR2_X1 U394 ( .A(n375), .B(KEYINPUT92), .ZN(n374) );
  NAND2_X1 U395 ( .A1(n373), .A2(n542), .ZN(n365) );
  NAND2_X1 U396 ( .A1(n578), .A2(n569), .ZN(n630) );
  XNOR2_X1 U397 ( .A(n483), .B(n484), .ZN(n734) );
  XNOR2_X1 U398 ( .A(n408), .B(KEYINPUT39), .ZN(n562) );
  INV_X1 U399 ( .A(n623), .ZN(n578) );
  INV_X1 U400 ( .A(KEYINPUT4), .ZN(n424) );
  INV_X1 U401 ( .A(KEYINPUT85), .ZN(n441) );
  AND2_X1 U402 ( .A1(n374), .A2(n594), .ZN(n597) );
  AND2_X1 U403 ( .A1(n388), .A2(n396), .ZN(n395) );
  NAND2_X1 U404 ( .A1(KEYINPUT65), .A2(n397), .ZN(n396) );
  NAND2_X1 U405 ( .A1(n394), .A2(n392), .ZN(n391) );
  INV_X1 U406 ( .A(n598), .ZN(n394) );
  NAND2_X1 U407 ( .A1(n393), .A2(n404), .ZN(n392) );
  XOR2_X1 U408 ( .A(KEYINPUT96), .B(KEYINPUT7), .Z(n469) );
  XNOR2_X1 U409 ( .A(n458), .B(n415), .ZN(n483) );
  INV_X1 U410 ( .A(KEYINPUT10), .ZN(n415) );
  XNOR2_X1 U411 ( .A(n467), .B(n355), .ZN(n733) );
  NAND2_X1 U412 ( .A1(G214), .A2(n511), .ZN(n613) );
  XNOR2_X1 U413 ( .A(n376), .B(n445), .ZN(n720) );
  XNOR2_X1 U414 ( .A(n436), .B(n435), .ZN(n376) );
  INV_X1 U415 ( .A(G119), .ZN(n435) );
  XNOR2_X1 U416 ( .A(n487), .B(n354), .ZN(n418) );
  XOR2_X1 U417 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n487) );
  XNOR2_X1 U418 ( .A(n486), .B(n485), .ZN(n488) );
  INV_X1 U419 ( .A(KEYINPUT23), .ZN(n485) );
  XNOR2_X1 U420 ( .A(G119), .B(KEYINPUT78), .ZN(n486) );
  XNOR2_X1 U421 ( .A(KEYINPUT76), .B(G110), .ZN(n437) );
  XOR2_X1 U422 ( .A(KEYINPUT68), .B(G101), .Z(n449) );
  XNOR2_X1 U423 ( .A(n446), .B(n407), .ZN(n659) );
  XNOR2_X1 U424 ( .A(n720), .B(n405), .ZN(n407) );
  XNOR2_X1 U425 ( .A(n718), .B(n421), .ZN(n446) );
  XNOR2_X1 U426 ( .A(n449), .B(n406), .ZN(n405) );
  XNOR2_X1 U427 ( .A(n584), .B(n583), .ZN(n649) );
  AND2_X1 U428 ( .A1(n386), .A2(n686), .ZN(n510) );
  XNOR2_X1 U429 ( .A(n590), .B(n410), .ZN(n409) );
  INV_X1 U430 ( .A(KEYINPUT104), .ZN(n410) );
  XNOR2_X1 U431 ( .A(n379), .B(n478), .ZN(n552) );
  OR2_X1 U432 ( .A1(n713), .A2(G902), .ZN(n379) );
  INV_X1 U433 ( .A(G472), .ZN(n384) );
  NAND2_X1 U434 ( .A1(n363), .A2(n362), .ZN(n591) );
  NAND2_X1 U435 ( .A1(n568), .A2(KEYINPUT0), .ZN(n362) );
  AND2_X1 U436 ( .A1(n364), .A2(n360), .ZN(n363) );
  BUF_X1 U437 ( .A(n631), .Z(n389) );
  NAND2_X1 U438 ( .A1(n404), .A2(KEYINPUT44), .ZN(n399) );
  XNOR2_X1 U439 ( .A(G146), .B(G125), .ZN(n458) );
  OR2_X1 U440 ( .A1(G237), .A2(G902), .ZN(n511) );
  XNOR2_X1 U441 ( .A(KEYINPUT3), .B(KEYINPUT70), .ZN(n436) );
  XNOR2_X1 U442 ( .A(G113), .B(G143), .ZN(n459) );
  XOR2_X1 U443 ( .A(G122), .B(G104), .Z(n460) );
  XOR2_X1 U444 ( .A(G140), .B(KEYINPUT94), .Z(n453) );
  INV_X1 U445 ( .A(n458), .ZN(n406) );
  XNOR2_X1 U446 ( .A(n422), .B(n444), .ZN(n421) );
  XNOR2_X1 U447 ( .A(n361), .B(n423), .ZN(n422) );
  XNOR2_X1 U448 ( .A(n441), .B(n424), .ZN(n423) );
  INV_X1 U449 ( .A(n745), .ZN(n411) );
  XNOR2_X1 U450 ( .A(n383), .B(n561), .ZN(n412) );
  AND2_X1 U451 ( .A1(n582), .A2(n521), .ZN(n509) );
  NAND2_X1 U452 ( .A1(n353), .A2(n351), .ZN(n364) );
  INV_X1 U453 ( .A(n352), .ZN(n367) );
  XNOR2_X1 U454 ( .A(n527), .B(KEYINPUT1), .ZN(n631) );
  XNOR2_X1 U455 ( .A(n592), .B(KEYINPUT6), .ZN(n582) );
  XNOR2_X1 U456 ( .A(n439), .B(G122), .ZN(n425) );
  XOR2_X1 U457 ( .A(KEYINPUT16), .B(KEYINPUT73), .Z(n439) );
  XNOR2_X1 U458 ( .A(n402), .B(KEYINPUT82), .ZN(n401) );
  INV_X1 U459 ( .A(G134), .ZN(n447) );
  XNOR2_X1 U460 ( .A(n470), .B(n380), .ZN(n472) );
  XNOR2_X1 U461 ( .A(n471), .B(n381), .ZN(n380) );
  INV_X1 U462 ( .A(KEYINPUT97), .ZN(n381) );
  NOR2_X1 U463 ( .A1(n617), .A2(n616), .ZN(n520) );
  XNOR2_X1 U464 ( .A(n427), .B(n426), .ZN(n587) );
  INV_X1 U465 ( .A(KEYINPUT35), .ZN(n426) );
  NAND2_X1 U466 ( .A1(n351), .A2(n365), .ZN(n568) );
  XNOR2_X1 U467 ( .A(n572), .B(KEYINPUT66), .ZN(n573) );
  NAND2_X1 U468 ( .A1(n529), .A2(n528), .ZN(n590) );
  XNOR2_X1 U469 ( .A(n377), .B(n720), .ZN(n507) );
  XNOR2_X1 U470 ( .A(n506), .B(n449), .ZN(n377) );
  XNOR2_X1 U471 ( .A(n417), .B(n490), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n418), .B(n488), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n705), .B(KEYINPUT120), .ZN(n706) );
  XNOR2_X1 U474 ( .A(n390), .B(n449), .ZN(n450) );
  XNOR2_X1 U475 ( .A(n484), .B(n357), .ZN(n390) );
  XNOR2_X1 U476 ( .A(n659), .B(n658), .ZN(n660) );
  INV_X1 U477 ( .A(n717), .ZN(n708) );
  AND2_X1 U478 ( .A1(n562), .A2(n686), .ZN(n534) );
  NAND2_X1 U479 ( .A1(n512), .A2(n356), .ZN(n387) );
  INV_X1 U480 ( .A(n587), .ZN(n746) );
  XNOR2_X1 U481 ( .A(n589), .B(KEYINPUT31), .ZN(n691) );
  AND2_X1 U482 ( .A1(n369), .A2(n371), .ZN(n351) );
  OR2_X1 U483 ( .A1(n567), .A2(n566), .ZN(n352) );
  AND2_X1 U484 ( .A1(n365), .A2(n366), .ZN(n353) );
  XOR2_X1 U485 ( .A(G128), .B(G110), .Z(n354) );
  XOR2_X1 U486 ( .A(KEYINPUT4), .B(G131), .Z(n355) );
  AND2_X1 U487 ( .A1(n537), .A2(n613), .ZN(n356) );
  AND2_X1 U488 ( .A1(G227), .A2(n736), .ZN(n357) );
  AND2_X1 U489 ( .A1(n511), .A2(G210), .ZN(n358) );
  AND2_X1 U490 ( .A1(n696), .A2(n599), .ZN(n359) );
  OR2_X1 U491 ( .A1(n352), .A2(n368), .ZN(n360) );
  INV_X1 U492 ( .A(KEYINPUT65), .ZN(n404) );
  INV_X1 U493 ( .A(KEYINPUT44), .ZN(n397) );
  XNOR2_X1 U494 ( .A(n361), .B(n447), .ZN(n467) );
  XNOR2_X2 U495 ( .A(n440), .B(G128), .ZN(n361) );
  NOR2_X1 U496 ( .A1(n367), .A2(KEYINPUT0), .ZN(n366) );
  INV_X1 U497 ( .A(KEYINPUT0), .ZN(n368) );
  NAND2_X1 U498 ( .A1(n537), .A2(n370), .ZN(n369) );
  NOR2_X1 U499 ( .A1(n372), .A2(n542), .ZN(n370) );
  NAND2_X1 U500 ( .A1(n372), .A2(n542), .ZN(n371) );
  INV_X1 U501 ( .A(n613), .ZN(n372) );
  INV_X1 U502 ( .A(n537), .ZN(n373) );
  NAND2_X1 U503 ( .A1(n691), .A2(n674), .ZN(n375) );
  XNOR2_X1 U504 ( .A(n510), .B(KEYINPUT101), .ZN(n538) );
  NAND2_X1 U505 ( .A1(n378), .A2(n575), .ZN(n695) );
  XNOR2_X1 U506 ( .A(n387), .B(n539), .ZN(n378) );
  XNOR2_X1 U507 ( .A(n530), .B(KEYINPUT30), .ZN(n531) );
  NOR2_X1 U508 ( .A1(n649), .A2(n591), .ZN(n585) );
  XNOR2_X2 U509 ( .A(n385), .B(n384), .ZN(n592) );
  NAND2_X1 U510 ( .A1(n623), .A2(n569), .ZN(n502) );
  XNOR2_X2 U511 ( .A(n495), .B(n494), .ZN(n623) );
  NOR2_X2 U512 ( .A1(n543), .A2(n568), .ZN(n685) );
  NOR2_X1 U513 ( .A1(n560), .A2(n414), .ZN(n413) );
  XNOR2_X2 U514 ( .A(n382), .B(KEYINPUT45), .ZN(n728) );
  NOR2_X2 U515 ( .A1(n403), .A2(n401), .ZN(n382) );
  NAND2_X1 U516 ( .A1(n413), .A2(n540), .ZN(n383) );
  INV_X1 U517 ( .A(n695), .ZN(n414) );
  OR2_X2 U518 ( .A1(n728), .A2(n419), .ZN(n420) );
  XNOR2_X1 U519 ( .A(n509), .B(KEYINPUT100), .ZN(n386) );
  NAND2_X1 U520 ( .A1(n703), .A2(G210), .ZN(n661) );
  XNOR2_X2 U521 ( .A(n608), .B(n607), .ZN(n703) );
  NAND2_X1 U522 ( .A1(n398), .A2(n598), .ZN(n388) );
  XNOR2_X1 U523 ( .A(n508), .B(n429), .ZN(n699) );
  NAND2_X1 U524 ( .A1(n432), .A2(n581), .ZN(n393) );
  NAND2_X1 U525 ( .A1(n400), .A2(n399), .ZN(n398) );
  NAND2_X1 U526 ( .A1(n432), .A2(KEYINPUT83), .ZN(n400) );
  NAND2_X1 U527 ( .A1(n434), .A2(n433), .ZN(n402) );
  NAND2_X1 U528 ( .A1(n548), .A2(n614), .ZN(n408) );
  AND2_X2 U529 ( .A1(n412), .A2(n411), .ZN(n605) );
  NAND2_X1 U530 ( .A1(n605), .A2(n359), .ZN(n419) );
  NAND2_X1 U531 ( .A1(n420), .A2(n601), .ZN(n606) );
  NOR2_X1 U532 ( .A1(n728), .A2(n735), .ZN(n644) );
  NAND2_X1 U533 ( .A1(n605), .A2(n696), .ZN(n735) );
  NAND2_X1 U534 ( .A1(n428), .A2(n586), .ZN(n427) );
  XNOR2_X1 U535 ( .A(n585), .B(KEYINPUT34), .ZN(n428) );
  XNOR2_X1 U536 ( .A(n450), .B(n448), .ZN(n429) );
  NOR2_X1 U537 ( .A1(n430), .A2(n582), .ZN(n595) );
  OR2_X1 U538 ( .A1(n430), .A2(n575), .ZN(n576) );
  XNOR2_X1 U539 ( .A(n574), .B(n573), .ZN(n430) );
  NAND2_X1 U540 ( .A1(n659), .A2(n479), .ZN(n431) );
  NAND2_X1 U541 ( .A1(n746), .A2(KEYINPUT44), .ZN(n433) );
  NOR2_X1 U542 ( .A1(n671), .A2(n597), .ZN(n434) );
  XNOR2_X1 U543 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U544 ( .A(n701), .B(n700), .ZN(n702) );
  INV_X1 U545 ( .A(KEYINPUT48), .ZN(n561) );
  XNOR2_X1 U546 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n583) );
  INV_X1 U547 ( .A(KEYINPUT64), .ZN(n607) );
  INV_X1 U548 ( .A(n527), .ZN(n528) );
  XNOR2_X1 U549 ( .A(n507), .B(n508), .ZN(n666) );
  XNOR2_X1 U550 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U551 ( .A(n713), .B(KEYINPUT122), .ZN(n714) );
  XNOR2_X1 U552 ( .A(n661), .B(n660), .ZN(n662) );
  INV_X1 U553 ( .A(n389), .ZN(n575) );
  XNOR2_X1 U554 ( .A(n610), .B(n609), .ZN(n612) );
  XNOR2_X1 U555 ( .A(n657), .B(n656), .ZN(G75) );
  XOR2_X2 U556 ( .A(G902), .B(KEYINPUT15), .Z(n599) );
  INV_X1 U557 ( .A(n599), .ZN(n479) );
  XOR2_X1 U558 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n443) );
  NAND2_X1 U559 ( .A1(G224), .A2(n736), .ZN(n442) );
  XNOR2_X1 U560 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U561 ( .A(G116), .B(G113), .ZN(n445) );
  NOR2_X1 U562 ( .A1(G902), .A2(n699), .ZN(n451) );
  XNOR2_X1 U563 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n465) );
  NOR2_X1 U564 ( .A1(G953), .A2(G237), .ZN(n503) );
  NAND2_X1 U565 ( .A1(G214), .A2(n503), .ZN(n452) );
  XNOR2_X1 U566 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U567 ( .A(KEYINPUT11), .B(KEYINPUT93), .Z(n455) );
  XNOR2_X1 U568 ( .A(G131), .B(KEYINPUT12), .ZN(n454) );
  XNOR2_X1 U569 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U570 ( .A(n457), .B(n456), .Z(n463) );
  XNOR2_X1 U571 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U572 ( .A(n483), .B(n461), .Z(n462) );
  XNOR2_X1 U573 ( .A(n463), .B(n462), .ZN(n704) );
  NOR2_X1 U574 ( .A1(G902), .A2(n704), .ZN(n464) );
  XNOR2_X1 U575 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U576 ( .A(G475), .B(n466), .ZN(n541) );
  XNOR2_X1 U577 ( .A(KEYINPUT98), .B(G478), .ZN(n478) );
  INV_X1 U578 ( .A(n467), .ZN(n473) );
  XNOR2_X1 U579 ( .A(G116), .B(KEYINPUT9), .ZN(n468) );
  XNOR2_X1 U580 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U581 ( .A(G107), .B(G122), .ZN(n471) );
  XNOR2_X1 U582 ( .A(n473), .B(n472), .ZN(n477) );
  NAND2_X1 U583 ( .A1(n736), .A2(G234), .ZN(n475) );
  XNOR2_X1 U584 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n474) );
  XNOR2_X1 U585 ( .A(n475), .B(n474), .ZN(n489) );
  NAND2_X1 U586 ( .A1(G217), .A2(n489), .ZN(n476) );
  XNOR2_X1 U587 ( .A(n477), .B(n476), .ZN(n713) );
  NOR2_X1 U588 ( .A1(n541), .A2(n552), .ZN(n686) );
  INV_X1 U589 ( .A(n686), .ZN(n689) );
  NAND2_X1 U590 ( .A1(n479), .A2(G234), .ZN(n480) );
  XNOR2_X1 U591 ( .A(n480), .B(KEYINPUT20), .ZN(n481) );
  XNOR2_X1 U592 ( .A(KEYINPUT90), .B(n481), .ZN(n491) );
  NAND2_X1 U593 ( .A1(n491), .A2(G221), .ZN(n482) );
  XOR2_X1 U594 ( .A(n482), .B(KEYINPUT21), .Z(n569) );
  NAND2_X1 U595 ( .A1(G221), .A2(n489), .ZN(n490) );
  XOR2_X1 U596 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n493) );
  NAND2_X1 U597 ( .A1(G217), .A2(n491), .ZN(n492) );
  XNOR2_X1 U598 ( .A(n493), .B(n492), .ZN(n494) );
  NAND2_X1 U599 ( .A1(G234), .A2(G237), .ZN(n496) );
  XNOR2_X1 U600 ( .A(n496), .B(KEYINPUT14), .ZN(n499) );
  NAND2_X1 U601 ( .A1(G902), .A2(n499), .ZN(n564) );
  NOR2_X1 U602 ( .A1(G900), .A2(n564), .ZN(n497) );
  NAND2_X1 U603 ( .A1(G953), .A2(n497), .ZN(n498) );
  XNOR2_X1 U604 ( .A(KEYINPUT99), .B(n498), .ZN(n500) );
  NAND2_X1 U605 ( .A1(G952), .A2(n499), .ZN(n643) );
  NOR2_X1 U606 ( .A1(G953), .A2(n643), .ZN(n567) );
  NOR2_X1 U607 ( .A1(n500), .A2(n567), .ZN(n501) );
  XOR2_X1 U608 ( .A(n501), .B(KEYINPUT79), .Z(n532) );
  NOR2_X1 U609 ( .A1(n502), .A2(n532), .ZN(n521) );
  XOR2_X1 U610 ( .A(G137), .B(KEYINPUT5), .Z(n505) );
  NAND2_X1 U611 ( .A1(n503), .A2(G210), .ZN(n504) );
  XNOR2_X1 U612 ( .A(n505), .B(n504), .ZN(n506) );
  INV_X1 U613 ( .A(n538), .ZN(n512) );
  NAND2_X1 U614 ( .A1(n512), .A2(n613), .ZN(n513) );
  NOR2_X1 U615 ( .A1(n575), .A2(n513), .ZN(n515) );
  XOR2_X1 U616 ( .A(KEYINPUT43), .B(KEYINPUT102), .Z(n514) );
  XNOR2_X1 U617 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U618 ( .A1(n373), .A2(n516), .ZN(n517) );
  XNOR2_X1 U619 ( .A(KEYINPUT103), .B(n517), .ZN(n745) );
  XOR2_X1 U620 ( .A(KEYINPUT38), .B(KEYINPUT75), .Z(n518) );
  NAND2_X1 U621 ( .A1(n614), .A2(n613), .ZN(n617) );
  INV_X1 U622 ( .A(n541), .ZN(n551) );
  NOR2_X1 U623 ( .A1(n552), .A2(n551), .ZN(n570) );
  INV_X1 U624 ( .A(n570), .ZN(n616) );
  XNOR2_X1 U625 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n519) );
  XNOR2_X1 U626 ( .A(n520), .B(n519), .ZN(n648) );
  XOR2_X1 U627 ( .A(KEYINPUT106), .B(KEYINPUT28), .Z(n523) );
  INV_X2 U628 ( .A(n592), .ZN(n628) );
  NAND2_X1 U629 ( .A1(n628), .A2(n521), .ZN(n522) );
  XOR2_X1 U630 ( .A(n523), .B(n522), .Z(n524) );
  XNOR2_X1 U631 ( .A(KEYINPUT107), .B(n525), .ZN(n543) );
  NOR2_X1 U632 ( .A1(n648), .A2(n543), .ZN(n526) );
  INV_X1 U633 ( .A(n630), .ZN(n529) );
  NAND2_X1 U634 ( .A1(n628), .A2(n613), .ZN(n530) );
  NOR2_X1 U635 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U636 ( .A(n535), .B(KEYINPUT46), .ZN(n540) );
  XNOR2_X1 U637 ( .A(KEYINPUT84), .B(KEYINPUT109), .ZN(n536) );
  XNOR2_X1 U638 ( .A(n536), .B(KEYINPUT36), .ZN(n539) );
  NAND2_X1 U639 ( .A1(n541), .A2(n552), .ZN(n692) );
  INV_X1 U640 ( .A(n692), .ZN(n681) );
  NOR2_X1 U641 ( .A1(n681), .A2(n686), .ZN(n618) );
  INV_X1 U642 ( .A(n618), .ZN(n594) );
  XNOR2_X1 U643 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n542) );
  NAND2_X1 U644 ( .A1(n594), .A2(n685), .ZN(n547) );
  INV_X1 U645 ( .A(n547), .ZN(n545) );
  INV_X1 U646 ( .A(KEYINPUT47), .ZN(n555) );
  NAND2_X1 U647 ( .A1(KEYINPUT74), .A2(n555), .ZN(n546) );
  INV_X1 U648 ( .A(n546), .ZN(n544) );
  NAND2_X1 U649 ( .A1(n545), .A2(n544), .ZN(n559) );
  NAND2_X1 U650 ( .A1(n547), .A2(n546), .ZN(n554) );
  NAND2_X1 U651 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U652 ( .A(KEYINPUT105), .B(n550), .ZN(n553) );
  AND2_X1 U653 ( .A1(n552), .A2(n551), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n553), .A2(n586), .ZN(n684) );
  NAND2_X1 U655 ( .A1(n554), .A2(n684), .ZN(n557) );
  NOR2_X1 U656 ( .A1(KEYINPUT74), .A2(n555), .ZN(n556) );
  NOR2_X1 U657 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U658 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U659 ( .A1(n562), .A2(n681), .ZN(n696) );
  NOR2_X1 U660 ( .A1(G898), .A2(n736), .ZN(n563) );
  XNOR2_X1 U661 ( .A(KEYINPUT87), .B(n563), .ZN(n722) );
  NOR2_X1 U662 ( .A1(n564), .A2(n722), .ZN(n565) );
  XNOR2_X1 U663 ( .A(n565), .B(KEYINPUT88), .ZN(n566) );
  INV_X1 U664 ( .A(n569), .ZN(n624) );
  NOR2_X1 U665 ( .A1(n591), .A2(n624), .ZN(n571) );
  NAND2_X1 U666 ( .A1(n571), .A2(n570), .ZN(n574) );
  XNOR2_X1 U667 ( .A(KEYINPUT22), .B(KEYINPUT72), .ZN(n572) );
  NOR2_X1 U668 ( .A1(n578), .A2(n576), .ZN(n577) );
  NAND2_X1 U669 ( .A1(n577), .A2(n592), .ZN(n679) );
  NOR2_X1 U670 ( .A1(n578), .A2(n389), .ZN(n579) );
  NAND2_X1 U671 ( .A1(n595), .A2(n579), .ZN(n580) );
  XNOR2_X2 U672 ( .A(n580), .B(KEYINPUT32), .ZN(n747) );
  NAND2_X1 U673 ( .A1(n679), .A2(n747), .ZN(n598) );
  INV_X1 U674 ( .A(KEYINPUT83), .ZN(n581) );
  NOR2_X2 U675 ( .A1(n631), .A2(n630), .ZN(n588) );
  NAND2_X1 U676 ( .A1(n588), .A2(n582), .ZN(n584) );
  NAND2_X1 U677 ( .A1(n628), .A2(n588), .ZN(n635) );
  NOR2_X1 U678 ( .A1(n591), .A2(n635), .ZN(n589) );
  NOR2_X1 U679 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U680 ( .A1(n593), .A2(n592), .ZN(n674) );
  NAND2_X1 U681 ( .A1(n389), .A2(n595), .ZN(n596) );
  NOR2_X1 U682 ( .A1(n623), .A2(n596), .ZN(n671) );
  NAND2_X1 U683 ( .A1(KEYINPUT2), .A2(n599), .ZN(n600) );
  XOR2_X1 U684 ( .A(n600), .B(KEYINPUT67), .Z(n601) );
  NAND2_X1 U685 ( .A1(KEYINPUT2), .A2(n696), .ZN(n602) );
  XNOR2_X1 U686 ( .A(KEYINPUT80), .B(n602), .ZN(n603) );
  NOR2_X1 U687 ( .A1(n728), .A2(n603), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n605), .A2(n604), .ZN(n647) );
  NAND2_X1 U689 ( .A1(n606), .A2(n647), .ZN(n608) );
  BUF_X2 U690 ( .A(n703), .Z(n712) );
  NAND2_X1 U691 ( .A1(G217), .A2(n712), .ZN(n610) );
  NOR2_X1 U692 ( .A1(G952), .A2(n736), .ZN(n611) );
  XNOR2_X1 U693 ( .A(KEYINPUT86), .B(n611), .ZN(n717) );
  NOR2_X1 U694 ( .A1(n612), .A2(n717), .ZN(G66) );
  NOR2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U699 ( .A1(n621), .A2(n649), .ZN(n622) );
  XOR2_X1 U700 ( .A(KEYINPUT117), .B(n622), .Z(n640) );
  XOR2_X1 U701 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n626) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n629), .B(KEYINPUT116), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n389), .A2(n630), .ZN(n632) );
  XNOR2_X1 U707 ( .A(KEYINPUT50), .B(n632), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U710 ( .A(KEYINPUT51), .B(n637), .ZN(n638) );
  NOR2_X1 U711 ( .A1(n648), .A2(n638), .ZN(n639) );
  NOR2_X1 U712 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n641), .B(KEYINPUT52), .ZN(n642) );
  NOR2_X1 U714 ( .A1(n643), .A2(n642), .ZN(n654) );
  NOR2_X1 U715 ( .A1(KEYINPUT2), .A2(n644), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(KEYINPUT81), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n652) );
  NOR2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U719 ( .A(KEYINPUT118), .B(n650), .Z(n651) );
  NAND2_X1 U720 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U722 ( .A1(n736), .A2(n655), .ZN(n657) );
  XNOR2_X1 U723 ( .A(KEYINPUT53), .B(KEYINPUT119), .ZN(n656) );
  XOR2_X1 U724 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n658) );
  NAND2_X1 U725 ( .A1(n662), .A2(n708), .ZN(n664) );
  INV_X1 U726 ( .A(KEYINPUT56), .ZN(n663) );
  XNOR2_X1 U727 ( .A(n664), .B(n663), .ZN(G51) );
  NAND2_X1 U728 ( .A1(n703), .A2(G472), .ZN(n668) );
  INV_X1 U729 ( .A(KEYINPUT62), .ZN(n665) );
  XNOR2_X1 U730 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U731 ( .A1(n669), .A2(n708), .ZN(n670) );
  XNOR2_X1 U732 ( .A(n670), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U733 ( .A(G101), .B(n671), .Z(G3) );
  NOR2_X1 U734 ( .A1(n689), .A2(n674), .ZN(n672) );
  XOR2_X1 U735 ( .A(KEYINPUT110), .B(n672), .Z(n673) );
  XNOR2_X1 U736 ( .A(G104), .B(n673), .ZN(G6) );
  NOR2_X1 U737 ( .A1(n674), .A2(n692), .ZN(n678) );
  XOR2_X1 U738 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n676) );
  XNOR2_X1 U739 ( .A(G107), .B(KEYINPUT111), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U741 ( .A(n678), .B(n677), .ZN(G9) );
  XNOR2_X1 U742 ( .A(G110), .B(KEYINPUT112), .ZN(n680) );
  XNOR2_X1 U743 ( .A(n680), .B(n679), .ZN(G12) );
  NAND2_X1 U744 ( .A1(n681), .A2(n685), .ZN(n683) );
  XOR2_X1 U745 ( .A(G128), .B(KEYINPUT29), .Z(n682) );
  XNOR2_X1 U746 ( .A(n683), .B(n682), .ZN(G30) );
  XNOR2_X1 U747 ( .A(G143), .B(n684), .ZN(G45) );
  NAND2_X1 U748 ( .A1(n686), .A2(n685), .ZN(n688) );
  XOR2_X1 U749 ( .A(G146), .B(KEYINPUT113), .Z(n687) );
  XNOR2_X1 U750 ( .A(n688), .B(n687), .ZN(G48) );
  NOR2_X1 U751 ( .A1(n689), .A2(n691), .ZN(n690) );
  XOR2_X1 U752 ( .A(G113), .B(n690), .Z(G15) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U754 ( .A(G116), .B(n693), .Z(G18) );
  XOR2_X1 U755 ( .A(G125), .B(KEYINPUT37), .Z(n694) );
  XNOR2_X1 U756 ( .A(n695), .B(n694), .ZN(G27) );
  XNOR2_X1 U757 ( .A(G134), .B(KEYINPUT114), .ZN(n697) );
  XNOR2_X1 U758 ( .A(n697), .B(n696), .ZN(G36) );
  NAND2_X1 U759 ( .A1(G469), .A2(n712), .ZN(n701) );
  XOR2_X1 U760 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n698) );
  XNOR2_X1 U761 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U762 ( .A1(n717), .A2(n702), .ZN(G54) );
  NAND2_X1 U763 ( .A1(n703), .A2(G475), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n704), .B(KEYINPUT59), .ZN(n705) );
  XNOR2_X1 U765 ( .A(n707), .B(n706), .ZN(n709) );
  NAND2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U767 ( .A(KEYINPUT60), .B(KEYINPUT121), .ZN(n710) );
  XNOR2_X1 U768 ( .A(n711), .B(n710), .ZN(G60) );
  NAND2_X1 U769 ( .A1(n712), .A2(G478), .ZN(n715) );
  NOR2_X1 U770 ( .A1(n717), .A2(n716), .ZN(G63) );
  XOR2_X1 U771 ( .A(n718), .B(KEYINPUT124), .Z(n719) );
  XNOR2_X1 U772 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U773 ( .A(G101), .B(n721), .ZN(n723) );
  NAND2_X1 U774 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U775 ( .A(n724), .B(KEYINPUT125), .ZN(n732) );
  XOR2_X1 U776 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n726) );
  NAND2_X1 U777 ( .A1(G224), .A2(G953), .ZN(n725) );
  XNOR2_X1 U778 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U779 ( .A1(n727), .A2(G898), .ZN(n730) );
  OR2_X1 U780 ( .A1(n728), .A2(G953), .ZN(n729) );
  NAND2_X1 U781 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U782 ( .A(n732), .B(n731), .ZN(G69) );
  XNOR2_X1 U783 ( .A(n734), .B(n733), .ZN(n738) );
  XNOR2_X1 U784 ( .A(n735), .B(n738), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n737), .A2(n736), .ZN(n743) );
  XNOR2_X1 U786 ( .A(G227), .B(n738), .ZN(n739) );
  XNOR2_X1 U787 ( .A(n739), .B(KEYINPUT126), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U789 ( .A1(n741), .A2(G953), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U791 ( .A(KEYINPUT127), .B(n744), .Z(G72) );
  XOR2_X1 U792 ( .A(G140), .B(n745), .Z(G42) );
  XOR2_X1 U793 ( .A(G122), .B(n746), .Z(G24) );
  XNOR2_X1 U794 ( .A(G119), .B(n747), .ZN(G21) );
  XOR2_X1 U795 ( .A(n748), .B(G131), .Z(G33) );
  XOR2_X1 U796 ( .A(G137), .B(n749), .Z(G39) );
endmodule

