//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G127gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(G134gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G127gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT69), .ZN(new_n208));
  XNOR2_X1  g007(.A(G113gat), .B(G120gat), .ZN(new_n209));
  OAI221_X1 g008(.A(new_n208), .B1(KEYINPUT69), .B2(new_n205), .C1(KEYINPUT1), .C2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n205), .A2(new_n207), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT70), .ZN(new_n213));
  INV_X1    g012(.A(G113gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(G120gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(G120gat), .ZN(new_n216));
  INV_X1    g015(.A(G120gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n212), .A2(new_n219), .A3(KEYINPUT71), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT71), .B1(new_n212), .B2(new_n219), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n210), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n227), .A2(new_n228), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n232), .B(new_n233), .C1(G183gat), .C2(G190gat), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT25), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n237), .A2(KEYINPUT64), .A3(new_n238), .A4(new_n231), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240));
  OAI22_X1  g039(.A1(new_n230), .A2(KEYINPUT65), .B1(new_n240), .B2(KEYINPUT24), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n238), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n239), .A2(new_n241), .B1(new_n233), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT25), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n233), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n237), .A2(new_n238), .B1(KEYINPUT64), .B2(new_n231), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n238), .A2(G183gat), .A3(G190gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n231), .A2(KEYINPUT64), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n244), .B(new_n246), .C1(new_n247), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n229), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n236), .B1(new_n245), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n246), .B1(new_n247), .B2(new_n250), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n227), .A2(new_n228), .ZN(new_n259));
  NAND2_X1  g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n261), .B1(new_n243), .B2(new_n244), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(KEYINPUT67), .A3(new_n236), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n255), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT27), .B(G183gat), .ZN(new_n266));
  INV_X1    g065(.A(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT28), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT26), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n225), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n271), .B2(new_n225), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n225), .A2(new_n271), .B1(new_n260), .B2(new_n270), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n230), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n224), .B1(new_n265), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n269), .A2(new_n275), .ZN(new_n278));
  AOI211_X1 g077(.A(new_n223), .B(new_n278), .C1(new_n255), .C2(new_n264), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n203), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT72), .B(G71gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G43gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  OR2_X1    g083(.A1(new_n284), .A2(KEYINPUT73), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(KEYINPUT73), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT33), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(KEYINPUT32), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT67), .B1(new_n263), .B2(new_n236), .ZN(new_n289));
  AOI211_X1 g088(.A(new_n254), .B(new_n235), .C1(new_n258), .C2(new_n262), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n276), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n223), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n265), .A2(new_n224), .A3(new_n276), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT32), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n294), .A2(new_n203), .B1(new_n295), .B2(KEYINPUT33), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n288), .B1(new_n296), .B2(new_n284), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(new_n202), .A3(new_n293), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT34), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n292), .A2(KEYINPUT34), .A3(new_n293), .A4(new_n202), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT33), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n280), .B1(KEYINPUT32), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n284), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n300), .A2(new_n301), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .A4(new_n288), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G211gat), .B(G218gat), .Z(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT76), .B(KEYINPUT22), .Z(new_n314));
  INV_X1    g113(.A(G211gat), .ZN(new_n315));
  INV_X1    g114(.A(G218gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n313), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n313), .A3(new_n318), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G226gat), .ZN(new_n324));
  INV_X1    g123(.A(G233gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(KEYINPUT29), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n265), .B2(new_n276), .ZN(new_n329));
  INV_X1    g128(.A(new_n326), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n235), .B1(new_n258), .B2(new_n262), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT77), .B1(new_n331), .B2(new_n278), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n276), .A2(new_n253), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n323), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n265), .A2(new_n326), .A3(new_n276), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(new_n334), .A3(new_n327), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n322), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(G92gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT78), .ZN(new_n343));
  INV_X1    g142(.A(G64gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n345), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n336), .A2(new_n339), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(KEYINPUT30), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n340), .A2(new_n350), .A3(new_n345), .ZN(new_n351));
  XOR2_X1   g150(.A(G141gat), .B(G148gat), .Z(new_n352));
  INV_X1    g151(.A(G155gat), .ZN(new_n353));
  INV_X1    g152(.A(G162gat), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT2), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G155gat), .B(G162gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n357), .A3(new_n355), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n359), .B2(new_n361), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n210), .B(new_n365), .C1(new_n221), .C2(new_n222), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n212), .A2(new_n219), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT71), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n220), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n365), .B1(new_n371), .B2(new_n210), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n364), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n361), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n223), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n376), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n378), .A2(new_n371), .A3(KEYINPUT4), .A4(new_n210), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n373), .A2(new_n374), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n374), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n223), .A2(KEYINPUT79), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n378), .B1(new_n382), .B2(new_n366), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n223), .A2(new_n376), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n380), .A2(new_n385), .A3(KEYINPUT5), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n366), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n387), .B2(new_n364), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT5), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT80), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT80), .B1(new_n377), .B2(new_n379), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n388), .B(new_n389), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(G85gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n386), .A2(new_n397), .A3(new_n392), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(KEYINPUT6), .A3(new_n398), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n349), .A2(new_n351), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G50gat), .ZN(new_n406));
  INV_X1    g205(.A(G78gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G106gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412));
  INV_X1    g211(.A(new_n321), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n412), .B1(new_n413), .B2(new_n319), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n378), .B1(new_n414), .B2(new_n360), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G22gat), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n323), .B1(KEYINPUT29), .B2(new_n362), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G228gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(new_n325), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n362), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n322), .B1(new_n423), .B2(new_n412), .ZN(new_n424));
  OAI21_X1  g223(.A(G22gat), .B1(new_n415), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n422), .B1(new_n419), .B2(new_n425), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n411), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n417), .B1(new_n416), .B2(new_n418), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n415), .A2(new_n424), .A3(G22gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n421), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n409), .B(KEYINPUT82), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n426), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n302), .B2(new_n297), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n311), .A2(new_n404), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT35), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n349), .A2(new_n351), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n402), .A2(new_n403), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n444), .A2(new_n446), .A3(KEYINPUT35), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n297), .A2(new_n302), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT75), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n297), .A2(KEYINPUT75), .A3(new_n302), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n450), .A2(new_n451), .B1(new_n303), .B2(new_n310), .ZN(new_n452));
  INV_X1    g251(.A(new_n435), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n404), .A2(new_n435), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT40), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT39), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n383), .A2(new_n381), .A3(new_n384), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n373), .B1(new_n390), .B2(new_n391), .ZN(new_n459));
  AOI211_X1 g258(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(new_n381), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n457), .A3(new_n381), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n397), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n456), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n349), .A2(new_n463), .A3(new_n351), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n458), .B1(new_n459), .B2(new_n381), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT39), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(new_n397), .A3(new_n461), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n399), .B1(new_n467), .B2(new_n456), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n336), .A2(KEYINPUT37), .A3(new_n339), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n471), .B1(new_n340), .B2(new_n472), .ZN(new_n473));
  AOI211_X1 g272(.A(KEYINPUT83), .B(KEYINPUT37), .C1(new_n336), .C2(new_n339), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n470), .B(new_n347), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n475), .A2(KEYINPUT38), .B1(new_n340), .B2(new_n345), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n291), .A2(new_n327), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n332), .A2(new_n334), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n326), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n322), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n337), .A2(new_n338), .A3(new_n322), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT83), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n340), .A2(new_n471), .A3(new_n472), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n345), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n329), .A2(new_n335), .A3(new_n323), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n322), .B1(new_n337), .B2(new_n338), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT38), .B1(new_n488), .B2(KEYINPUT37), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n445), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n469), .B1(new_n476), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n455), .B1(new_n491), .B2(new_n435), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n311), .A2(KEYINPUT36), .A3(new_n448), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n452), .B2(KEYINPUT36), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n442), .A2(new_n454), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G120gat), .B(G148gat), .ZN(new_n496));
  INV_X1    g295(.A(G176gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n498), .B(G204gat), .Z(new_n499));
  NAND2_X1  g298(.A1(G230gat), .A2(G233gat), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n500), .B(KEYINPUT101), .Z(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT100), .B(KEYINPUT10), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n504));
  INV_X1    g303(.A(G57gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(G64gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(G64gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n344), .A2(KEYINPUT93), .A3(G57gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G71gat), .A2(G78gat), .ZN(new_n510));
  INV_X1    g309(.A(G71gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n407), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT9), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n509), .A2(new_n514), .A3(KEYINPUT94), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT8), .ZN(new_n521));
  NAND2_X1  g320(.A1(G85gat), .A2(G92gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G85gat), .ZN(new_n525));
  INV_X1    g324(.A(G92gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n521), .A2(new_n524), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G99gat), .B(G106gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(KEYINPUT8), .A2(new_n520), .B1(new_n525), .B2(new_n526), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(new_n530), .A3(new_n524), .A4(new_n528), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n344), .A2(G57gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n505), .A2(G64gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n510), .A2(new_n513), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n344), .A2(G57gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n507), .A2(new_n541), .A3(KEYINPUT92), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n512), .A2(new_n510), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n519), .A2(new_n535), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n532), .A2(KEYINPUT98), .A3(new_n534), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT98), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n529), .A2(new_n548), .A3(new_n531), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n519), .A2(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n503), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n517), .A2(new_n518), .B1(new_n543), .B2(new_n544), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n549), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT10), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n501), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n501), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n546), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n499), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT94), .B1(new_n509), .B2(new_n514), .ZN(new_n559));
  INV_X1    g358(.A(new_n518), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n545), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n553), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n552), .A2(new_n535), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n502), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n554), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n556), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n557), .ZN(new_n567));
  INV_X1    g366(.A(new_n499), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n558), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G29gat), .ZN(new_n571));
  INV_X1    g370(.A(G36gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT14), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT14), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(G29gat), .B2(G36gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G29gat), .A2(G36gat), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(G43gat), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT88), .B1(new_n578), .B2(G50gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT88), .ZN(new_n580));
  INV_X1    g379(.A(G50gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(G43gat), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n579), .B(new_n582), .C1(G43gat), .C2(new_n581), .ZN(new_n583));
  XOR2_X1   g382(.A(KEYINPUT87), .B(KEYINPUT15), .Z(new_n584));
  NAND3_X1  g383(.A1(new_n577), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT15), .B1(new_n578), .B2(G50gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n581), .A2(G43gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n577), .A2(KEYINPUT86), .A3(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT86), .A4(new_n576), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n587), .B2(new_n586), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT91), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n593), .A2(KEYINPUT17), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(KEYINPUT17), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n590), .B(new_n588), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n597), .A2(new_n593), .A3(KEYINPUT17), .A4(new_n585), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n600));
  INV_X1    g399(.A(G15gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n417), .ZN(new_n602));
  NAND2_X1  g401(.A1(G15gat), .A2(G22gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT89), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n602), .A2(KEYINPUT89), .A3(new_n603), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(G1gat), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G1gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT16), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n606), .B2(new_n607), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n600), .B(G8gat), .C1(new_n609), .C2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n600), .A2(G8gat), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n600), .A2(G8gat), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .A4(new_n608), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n599), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n592), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n613), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n622), .B(KEYINPUT13), .Z(new_n626));
  INV_X1    g425(.A(new_n621), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n620), .B1(new_n613), .B2(new_n617), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n619), .A2(KEYINPUT18), .A3(new_n621), .A4(new_n622), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G169gat), .B(G197gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n625), .A2(new_n629), .A3(new_n630), .A4(new_n637), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n495), .A2(new_n570), .A3(new_n642), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n613), .A2(new_n617), .B1(KEYINPUT21), .B2(new_n552), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT96), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n552), .A2(KEYINPUT21), .ZN(new_n648));
  XOR2_X1   g447(.A(G127gat), .B(G155gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT95), .ZN(new_n652));
  XOR2_X1   g451(.A(G183gat), .B(G211gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n647), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n553), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n599), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G232gat), .A2(G233gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT97), .Z(new_n660));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n592), .B1(new_n549), .B2(new_n547), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n658), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(G190gat), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n664), .B1(new_n599), .B2(new_n657), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n267), .A3(new_n663), .ZN(new_n669));
  AOI21_X1  g468(.A(G218gat), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n267), .B1(new_n668), .B2(new_n663), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n553), .B1(new_n596), .B2(new_n598), .ZN(new_n672));
  NOR4_X1   g471(.A1(new_n672), .A2(G190gat), .A3(new_n662), .A4(new_n664), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n671), .A2(new_n673), .A3(new_n316), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT99), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n667), .A2(G218gat), .A3(new_n669), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n316), .B1(new_n671), .B2(new_n673), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n661), .ZN(new_n680));
  XNOR2_X1  g479(.A(G134gat), .B(G162gat), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n675), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n676), .A2(new_n677), .A3(new_n678), .A4(new_n682), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n656), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n643), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n445), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(new_n610), .ZN(G1324gat));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT103), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n643), .A2(new_n688), .A3(new_n444), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n696), .A2(new_n694), .A3(new_n693), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n696), .B(KEYINPUT102), .Z(new_n698));
  NOR2_X1   g497(.A1(new_n694), .A2(G8gat), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n695), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(G1325gat));
  NOR2_X1   g499(.A1(new_n689), .A2(new_n601), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n450), .A2(new_n451), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n311), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT36), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT104), .B1(new_n705), .B2(new_n493), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n493), .B(KEYINPUT104), .C1(new_n452), .C2(KEYINPUT36), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n643), .A2(new_n688), .A3(new_n452), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n701), .A2(new_n709), .B1(new_n601), .B2(new_n710), .ZN(G1326gat));
  NOR2_X1   g510(.A1(new_n689), .A2(new_n453), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT105), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n712), .B(new_n714), .ZN(G1327gat));
  INV_X1    g514(.A(new_n656), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n642), .A2(new_n570), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n495), .A2(new_n686), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n571), .A3(new_n446), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n492), .A2(new_n494), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n437), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT84), .B1(new_n437), .B2(KEYINPUT35), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n454), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n686), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT106), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n729), .B(KEYINPUT44), .C1(new_n495), .C2(new_n686), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n684), .A2(new_n685), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n491), .A2(new_n435), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n494), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n732), .A2(new_n455), .B1(new_n734), .B2(new_n707), .ZN(new_n735));
  INV_X1    g534(.A(new_n725), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n727), .B(new_n731), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n728), .A2(new_n730), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n718), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n738), .A2(new_n446), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n721), .B1(new_n571), .B2(new_n740), .ZN(G1328gat));
  NAND3_X1  g540(.A1(new_n738), .A2(new_n444), .A3(new_n739), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G36gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n719), .A2(new_n572), .A3(new_n444), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n744), .A2(new_n746), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n743), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT108), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n743), .A2(new_n752), .A3(new_n748), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1329gat));
  NAND3_X1  g553(.A1(new_n719), .A2(new_n578), .A3(new_n452), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT109), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n709), .A3(new_n739), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n756), .A2(new_n758), .A3(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1330gat));
  NAND4_X1  g562(.A1(new_n738), .A2(G50gat), .A3(new_n435), .A4(new_n739), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n719), .A2(new_n435), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(G50gat), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g566(.A(new_n570), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n492), .B1(new_n706), .B2(new_n708), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n725), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n687), .A2(new_n641), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n445), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT110), .B(G57gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1332gat));
  XNOR2_X1  g574(.A(new_n443), .B(KEYINPUT111), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  AND2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n778), .B2(new_n779), .ZN(G1333gat));
  OAI21_X1  g581(.A(new_n511), .B1(new_n772), .B2(new_n703), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n770), .A2(G71gat), .A3(new_n709), .A4(new_n771), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g585(.A1(new_n772), .A2(new_n453), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(new_n407), .ZN(G1335gat));
  AOI21_X1  g587(.A(new_n686), .B1(new_n769), .B2(new_n725), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n656), .A2(new_n641), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(KEYINPUT112), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n768), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n793), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(KEYINPUT112), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n789), .A2(new_n795), .A3(new_n790), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n525), .B1(new_n798), .B2(new_n445), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n656), .A2(new_n768), .A3(new_n641), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n738), .A2(G85gat), .A3(new_n446), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n799), .A2(new_n801), .ZN(G1336gat));
  NAND4_X1  g601(.A1(new_n794), .A2(new_n526), .A3(new_n797), .A4(new_n776), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n738), .A2(new_n776), .A3(new_n800), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n526), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n738), .A2(new_n444), .A3(new_n800), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n808), .A2(KEYINPUT113), .A3(new_n803), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT52), .B1(new_n808), .B2(KEYINPUT113), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(G1337gat));
  NAND3_X1  g610(.A1(new_n738), .A2(new_n709), .A3(new_n800), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G99gat), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n798), .A2(G99gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n703), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n738), .A2(new_n435), .A3(new_n800), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT114), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n738), .A2(new_n818), .A3(new_n435), .A4(new_n800), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(G106gat), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n453), .A2(G106gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n794), .A2(new_n797), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n816), .A2(G106gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n822), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1339gat));
  NOR3_X1   g628(.A1(new_n627), .A2(new_n628), .A3(new_n626), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n622), .B1(new_n619), .B2(new_n621), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n636), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n640), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT116), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n833), .A2(KEYINPUT116), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n551), .A2(new_n501), .A3(new_n554), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n566), .A2(new_n836), .A3(KEYINPUT54), .ZN(new_n837));
  XNOR2_X1  g636(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n555), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n839), .A3(new_n499), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n837), .A2(new_n839), .A3(KEYINPUT55), .A4(new_n499), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n842), .A2(new_n569), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n731), .A2(new_n834), .A3(new_n835), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n570), .A2(new_n640), .A3(new_n832), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n842), .A2(new_n569), .A3(new_n843), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n847), .B(new_n848), .C1(new_n642), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n686), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n656), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n687), .A2(new_n570), .A3(new_n641), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(new_n435), .A3(new_n703), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n776), .A2(new_n445), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n857), .B(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n214), .B1(new_n859), .B2(new_n641), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n854), .A2(new_n445), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n311), .A2(new_n436), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n777), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(G113gat), .A3(new_n642), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n860), .A2(new_n865), .ZN(G1340gat));
  AOI21_X1  g665(.A(new_n217), .B1(new_n859), .B2(new_n570), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n864), .A2(G120gat), .A3(new_n768), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  NAND3_X1  g668(.A1(new_n859), .A2(G127gat), .A3(new_n656), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n204), .B1(new_n864), .B2(new_n716), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  NOR2_X1   g671(.A1(new_n444), .A2(new_n686), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n863), .A2(new_n206), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT119), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(KEYINPUT121), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n731), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT120), .B1(new_n879), .B2(G134gat), .ZN(new_n881));
  OAI221_X1 g680(.A(new_n877), .B1(new_n875), .B2(new_n878), .C1(new_n880), .C2(new_n881), .ZN(G1343gat));
  NOR2_X1   g681(.A1(new_n709), .A2(new_n453), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(new_n861), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n777), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n885), .A2(G141gat), .A3(new_n642), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n854), .B2(new_n453), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n846), .A2(KEYINPUT123), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n844), .B2(new_n641), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n846), .A2(KEYINPUT123), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n892), .A2(new_n893), .B1(new_n685), .B2(new_n684), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n684), .A2(new_n844), .A3(new_n685), .A4(new_n835), .ZN(new_n895));
  INV_X1    g694(.A(new_n834), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n716), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n771), .A2(new_n768), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n453), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT57), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT122), .B(new_n887), .C1(new_n854), .C2(new_n453), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n890), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n709), .A2(new_n445), .A3(new_n776), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G141gat), .B1(new_n905), .B2(new_n642), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT58), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1344gat));
  OR3_X1    g710(.A1(new_n885), .A2(G148gat), .A3(new_n768), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n903), .A2(new_n570), .A3(new_n904), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(G148gat), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT124), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT57), .B(new_n435), .C1(new_n852), .C2(new_n853), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n570), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n904), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n914), .B1(new_n920), .B2(G148gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n912), .B1(new_n916), .B2(new_n921), .ZN(G1345gat));
  NOR3_X1   g721(.A1(new_n905), .A2(new_n353), .A3(new_n716), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n884), .A2(new_n656), .A3(new_n777), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n353), .B2(new_n924), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n905), .B2(new_n686), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n884), .A2(new_n354), .A3(new_n873), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n446), .A2(new_n443), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n855), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n642), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n854), .A2(new_n446), .A3(new_n777), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n862), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n933), .A2(G169gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n934), .B2(new_n642), .ZN(G1348gat));
  NOR3_X1   g734(.A1(new_n930), .A2(new_n497), .A3(new_n768), .ZN(new_n936));
  INV_X1    g735(.A(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n570), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n936), .B1(new_n497), .B2(new_n938), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n930), .B2(new_n716), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n656), .A2(new_n266), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n930), .B2(new_n686), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT61), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n937), .A2(new_n267), .A3(new_n731), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1351gat));
  NAND2_X1  g746(.A1(new_n883), .A2(new_n932), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(G197gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(new_n950), .A3(new_n641), .ZN(new_n951));
  INV_X1    g750(.A(new_n929), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n952), .B1(new_n734), .B2(new_n707), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n918), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(new_n641), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n955), .B2(new_n950), .ZN(G1352gat));
  OR3_X1    g755(.A1(new_n948), .A2(G204gat), .A3(new_n768), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n919), .A2(new_n953), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G204gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n959), .A2(new_n960), .A3(new_n962), .A4(new_n963), .ZN(G1353gat));
  NAND3_X1  g763(.A1(new_n918), .A2(new_n656), .A3(new_n953), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n918), .A2(new_n967), .A3(new_n656), .A4(new_n953), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n966), .A2(G211gat), .A3(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n966), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n949), .A2(new_n315), .A3(new_n656), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT127), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n973), .A2(new_n977), .A3(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n949), .B2(new_n731), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n686), .A2(new_n316), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n954), .B2(new_n981), .ZN(G1355gat));
endmodule


