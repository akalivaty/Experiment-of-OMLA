//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT41), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT88), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT83), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT84), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n214), .B2(KEYINPUT15), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n215), .B(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n210), .B(KEYINPUT85), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n221), .B(new_n222), .C1(new_n211), .C2(new_n212), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT17), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT90), .B(G85gat), .Z(new_n226));
  INV_X1    g025(.A(G92gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n226), .A2(new_n227), .B1(KEYINPUT8), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230));
  INV_X1    g029(.A(G85gat), .ZN(new_n231));
  OAI211_X1 g030(.A(KEYINPUT89), .B(new_n230), .C1(new_n231), .C2(new_n227), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT89), .B1(new_n231), .B2(new_n227), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT89), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(G85gat), .A3(G92gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT7), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n229), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G99gat), .B(G106gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT91), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n224), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n242), .B(new_n243), .C1(new_n203), .C2(new_n202), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G134gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(G190gat), .B(G218gat), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n245), .A2(new_n246), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n207), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n245), .A2(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(new_n246), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n206), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G15gat), .B(G22gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT16), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(G1gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(G1gat), .B2(new_n254), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G8gat), .ZN(new_n258));
  XOR2_X1   g057(.A(G57gat), .B(G64gat), .Z(new_n259));
  AND2_X1   g058(.A1(G71gat), .A2(G78gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(KEYINPUT9), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G71gat), .B(G78gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(KEYINPUT21), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(G183gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(G231gat), .A2(G233gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n265), .B(new_n266), .Z(new_n267));
  XOR2_X1   g066(.A(G127gat), .B(G155gat), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT20), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n267), .B(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n263), .A2(KEYINPUT21), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(G211gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n271), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n270), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n253), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(G85gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT0), .B(G57gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284));
  XNOR2_X1  g083(.A(G141gat), .B(G148gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n286), .B1(G155gat), .B2(G162gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G155gat), .B(G162gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n284), .B(new_n289), .C1(new_n285), .C2(new_n287), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G113gat), .B(G120gat), .ZN(new_n294));
  OAI21_X1  g093(.A(G127gat), .B1(new_n294), .B2(KEYINPUT1), .ZN(new_n295));
  INV_X1    g094(.A(G120gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G113gat), .ZN(new_n297));
  INV_X1    g096(.A(G113gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G120gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301));
  INV_X1    g100(.A(G127gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n295), .A2(new_n303), .A3(G134gat), .ZN(new_n304));
  INV_X1    g103(.A(G134gat), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n302), .B1(new_n300), .B2(new_n301), .ZN(new_n306));
  AOI211_X1 g105(.A(KEYINPUT1), .B(G127gat), .C1(new_n297), .C2(new_n299), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT73), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n293), .A2(new_n308), .A3(new_n311), .A4(new_n304), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n304), .ZN(new_n313));
  INV_X1    g112(.A(new_n293), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n310), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n283), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n310), .A2(new_n312), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT74), .ZN(new_n324));
  INV_X1    g123(.A(new_n309), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(new_n322), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n328), .A3(new_n322), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT3), .B1(new_n291), .B2(new_n292), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n313), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n317), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n320), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT75), .B1(new_n325), .B2(new_n322), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n321), .B2(new_n322), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n310), .A2(KEYINPUT75), .A3(KEYINPUT4), .A4(new_n312), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n318), .A2(KEYINPUT5), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n282), .B1(new_n337), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n328), .B1(new_n321), .B2(new_n322), .ZN(new_n346));
  AOI211_X1 g145(.A(KEYINPUT74), .B(KEYINPUT4), .C1(new_n310), .C2(new_n312), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n346), .A2(new_n347), .A3(new_n326), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n319), .B1(new_n348), .B2(new_n335), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n341), .A2(new_n343), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n281), .A3(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(KEYINPUT76), .B(KEYINPUT6), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n345), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G197gat), .B(G204gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(G211gat), .A2(G218gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT22), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  OR2_X1    g158(.A1(G211gat), .A2(G218gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT69), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n356), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n360), .B2(new_n356), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n359), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n356), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT69), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n367), .A2(new_n358), .A3(new_n355), .A4(new_n362), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G226gat), .ZN(new_n370));
  INV_X1    g169(.A(G233gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G190gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n375));
  AND2_X1   g174(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n374), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n380));
  AOI21_X1  g179(.A(G190gat), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n378), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR3_X1   g186(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G169gat), .ZN(new_n390));
  AND2_X1   g189(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT23), .B(new_n390), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(G183gat), .A3(G190gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT23), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(G169gat), .B2(G176gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT24), .ZN(new_n400));
  NOR2_X1   g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n397), .B(new_n399), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  OAI22_X1  g201(.A1(new_n383), .A2(new_n389), .B1(new_n395), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT65), .ZN(new_n405));
  INV_X1    g204(.A(G176gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n406), .A3(KEYINPUT23), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n407), .B2(new_n386), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n405), .A3(new_n386), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT25), .B1(new_n411), .B2(new_n402), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(KEYINPUT70), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT70), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n407), .A2(new_n405), .A3(new_n386), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(new_n408), .ZN(new_n417));
  INV_X1    g216(.A(new_n402), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n414), .B1(new_n419), .B2(new_n403), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n373), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n403), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n422), .A2(KEYINPUT29), .A3(new_n372), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n369), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n413), .A2(new_n420), .A3(new_n425), .A4(new_n373), .ZN(new_n426));
  INV_X1    g225(.A(new_n369), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n372), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT71), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT71), .B1(new_n424), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT37), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n424), .A2(new_n429), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n436), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT38), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n421), .A2(new_n423), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n438), .B1(new_n444), .B2(new_n427), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n428), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n369), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT38), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n440), .A2(new_n443), .B1(new_n439), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n282), .B(new_n352), .C1(new_n337), .C2(new_n344), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n354), .B(new_n449), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n369), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n454), .A2(KEYINPUT78), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n365), .A2(new_n368), .A3(new_n425), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT3), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n314), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n454), .A2(KEYINPUT78), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G228gat), .A2(G233gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT77), .Z(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n462), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(new_n465), .A3(new_n454), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT31), .B(G50gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G78gat), .B(G106gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(G22gat), .ZN(new_n471));
  INV_X1    g270(.A(new_n468), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n464), .A2(new_n472), .A3(new_n466), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n471), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n464), .B2(new_n466), .ZN(new_n476));
  INV_X1    g275(.A(new_n466), .ZN(new_n477));
  AOI211_X1 g276(.A(new_n468), .B(new_n477), .C1(new_n461), .C2(new_n463), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n435), .B1(new_n430), .B2(new_n431), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(KEYINPUT30), .A3(new_n441), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n441), .A2(KEYINPUT30), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n341), .A2(new_n318), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n281), .B1(new_n487), .B2(KEYINPUT39), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT39), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n316), .A2(new_n318), .ZN(new_n490));
  AOI211_X1 g289(.A(new_n489), .B(new_n490), .C1(new_n341), .C2(new_n318), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n486), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT79), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT79), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(new_n486), .C1(new_n488), .C2(new_n491), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n485), .A2(new_n493), .A3(new_n345), .A4(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n488), .ZN(new_n497));
  INV_X1    g296(.A(new_n491), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT40), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT80), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT80), .A4(KEYINPUT40), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n453), .B(new_n480), .C1(new_n496), .C2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G15gat), .B(G43gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(G71gat), .B(G99gat), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n505), .B(new_n506), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G227gat), .A2(G233gat), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n404), .A2(new_n412), .B1(new_n304), .B2(new_n308), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n313), .A2(new_n419), .A3(new_n403), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n404), .A2(new_n304), .A3(new_n308), .A4(new_n412), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n313), .B1(new_n419), .B2(new_n403), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n509), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT32), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT67), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n513), .A2(new_n521), .A3(KEYINPUT32), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n516), .A2(new_n509), .A3(new_n517), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT68), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n513), .B(KEYINPUT32), .C1(new_n514), .C2(new_n508), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n523), .B2(new_n530), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n531), .B2(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n354), .A2(new_n450), .B1(new_n482), .B2(new_n483), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n474), .A2(new_n479), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n504), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n354), .B1(new_n451), .B2(new_n452), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n530), .ZN(new_n544));
  INV_X1    g343(.A(new_n529), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT82), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT82), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n531), .B2(new_n532), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n540), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n543), .A2(new_n551), .A3(new_n484), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT35), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n540), .A2(new_n533), .ZN(new_n554));
  AOI221_X4 g353(.A(new_n553), .B1(new_n482), .B2(new_n483), .C1(new_n354), .C2(new_n450), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n552), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n542), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n258), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n225), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n224), .A2(new_n258), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(KEYINPUT18), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT86), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n224), .B2(new_n258), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(new_n561), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n560), .B(KEYINPUT13), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(KEYINPUT18), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  INV_X1    g370(.A(G197gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT11), .B(G169gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT12), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n563), .A2(new_n576), .A3(new_n569), .A4(new_n568), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n237), .A2(new_n238), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n263), .B1(new_n582), .B2(KEYINPUT92), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(new_n239), .Z(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT93), .Z(new_n587));
  INV_X1    g386(.A(KEYINPUT10), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n240), .A2(KEYINPUT10), .A3(new_n263), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n585), .B(KEYINPUT95), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595));
  INV_X1    g394(.A(G148gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT94), .B(G120gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n591), .A2(new_n585), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n581), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n277), .A2(new_n557), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT96), .Z(new_n607));
  NAND2_X1  g406(.A1(new_n354), .A2(new_n450), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT97), .B(G1gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(G1324gat));
  INV_X1    g411(.A(new_n607), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n484), .ZN(new_n614));
  NAND2_X1  g413(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n615));
  INV_X1    g414(.A(G8gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n255), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT42), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n616), .B2(new_n614), .ZN(G1325gat));
  NAND2_X1  g419(.A1(new_n550), .A2(new_n548), .ZN(new_n621));
  AOI21_X1  g420(.A(G15gat), .B1(new_n607), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n537), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n624), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n540), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G22gat), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT98), .B(KEYINPUT43), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1327gat));
  OAI21_X1  g428(.A(new_n623), .B1(new_n538), .B2(new_n480), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n496), .A2(new_n503), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n345), .A2(new_n351), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n349), .A2(new_n350), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT81), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n282), .A4(new_n352), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n632), .A2(new_n353), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n540), .B1(new_n637), .B2(new_n449), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n630), .B1(new_n631), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n621), .A2(new_n484), .A3(new_n480), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n553), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n538), .A2(KEYINPUT35), .A3(new_n554), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n253), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n605), .A2(new_n276), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n211), .A3(new_n609), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT99), .B(KEYINPUT45), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n557), .B2(new_n253), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n249), .A2(new_n252), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n621), .A2(new_n484), .A3(new_n480), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT35), .B1(new_n653), .B2(new_n543), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n538), .A2(KEYINPUT35), .A3(new_n554), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT100), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n657), .A3(new_n642), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n652), .B1(new_n659), .B2(new_n542), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n651), .B1(new_n660), .B2(new_n650), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT101), .B1(new_n661), .B2(new_n645), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n641), .A2(new_n657), .A3(new_n642), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n657), .B1(new_n641), .B2(new_n642), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n542), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n650), .A3(new_n253), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n644), .A2(KEYINPUT44), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n669));
  INV_X1    g468(.A(new_n645), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n662), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n609), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT102), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n649), .B1(new_n674), .B2(new_n211), .ZN(G1328gat));
  NAND3_X1  g474(.A1(new_n646), .A2(new_n212), .A3(new_n485), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT46), .Z(new_n677));
  AOI21_X1  g476(.A(new_n484), .B1(new_n662), .B2(new_n671), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n678), .B2(new_n212), .ZN(G1329gat));
  NAND2_X1  g478(.A1(new_n668), .A2(new_n670), .ZN(new_n680));
  OAI21_X1  g479(.A(G43gat), .B1(new_n680), .B2(new_n623), .ZN(new_n681));
  INV_X1    g480(.A(G43gat), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n646), .A2(new_n682), .A3(new_n621), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(KEYINPUT47), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n623), .B1(new_n662), .B2(new_n671), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT104), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n669), .B1(new_n668), .B2(new_n670), .ZN(new_n687));
  AOI211_X1 g486(.A(KEYINPUT101), .B(new_n645), .C1(new_n666), .C2(new_n667), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n537), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n690), .A3(G43gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n683), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n692), .B2(new_n694), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n684), .B1(new_n695), .B2(new_n696), .ZN(G1330gat));
  XOR2_X1   g496(.A(new_n646), .B(KEYINPUT106), .Z(new_n698));
  NOR2_X1   g497(.A1(new_n480), .A2(G50gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT107), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G50gat), .B1(new_n680), .B2(new_n480), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(KEYINPUT48), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT108), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n672), .A2(new_n540), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n705), .A2(G50gat), .B1(new_n700), .B2(new_n698), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(KEYINPUT48), .B2(new_n706), .ZN(G1331gat));
  AND3_X1   g506(.A1(new_n665), .A2(new_n277), .A3(new_n581), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n604), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n609), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g511(.A1(new_n709), .A2(new_n484), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  AND2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n713), .B2(new_n714), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n709), .B2(new_n623), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n621), .B(KEYINPUT109), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n719), .A2(G71gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n709), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g521(.A1(new_n710), .A2(new_n540), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g523(.A1(new_n275), .A2(new_n580), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n604), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT110), .Z(new_n727));
  AND2_X1   g526(.A1(new_n668), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(new_n608), .A3(new_n226), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n660), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n725), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n660), .A2(new_n725), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT51), .Z(new_n733));
  OAI211_X1 g532(.A(new_n604), .B(new_n731), .C1(new_n733), .C2(KEYINPUT111), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(new_n608), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n730), .B1(new_n735), .B2(new_n226), .ZN(G1336gat));
  AND4_X1   g535(.A1(new_n227), .A2(new_n733), .A3(new_n485), .A4(new_n604), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n227), .B1(new_n728), .B2(new_n485), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT52), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(KEYINPUT52), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n485), .A2(new_n227), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n734), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(G1337gat));
  XNOR2_X1  g542(.A(KEYINPUT112), .B(G99gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n729), .B2(new_n623), .ZN(new_n745));
  INV_X1    g544(.A(new_n621), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n746), .A2(new_n744), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n734), .B2(new_n747), .ZN(G1338gat));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749));
  OAI21_X1  g548(.A(G106gat), .B1(new_n729), .B2(new_n480), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n480), .A2(G106gat), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n749), .B(new_n750), .C1(new_n734), .C2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n733), .A2(new_n604), .A3(new_n751), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT113), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n733), .A2(new_n756), .A3(new_n604), .A4(new_n751), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n755), .A2(new_n750), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n758), .B2(new_n749), .ZN(G1339gat));
  NOR2_X1   g558(.A1(new_n593), .A2(KEYINPUT54), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n599), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n602), .B(KEYINPUT54), .C1(new_n592), .C2(new_n591), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(KEYINPUT55), .A3(new_n762), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(new_n603), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n762), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n580), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n566), .A2(new_n567), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n575), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n604), .A2(new_n579), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n652), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n764), .A2(new_n767), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n579), .A2(new_n773), .A3(new_n772), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n253), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n275), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n253), .A2(new_n276), .A3(new_n604), .A4(new_n580), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n609), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR4_X1   g581(.A1(new_n782), .A2(new_n485), .A3(new_n540), .A4(new_n533), .ZN(new_n783));
  AOI21_X1  g582(.A(G113gat), .B1(new_n783), .B2(new_n580), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n782), .A2(new_n640), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n581), .A2(new_n298), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(G1340gat));
  INV_X1    g586(.A(new_n785), .ZN(new_n788));
  INV_X1    g587(.A(new_n604), .ZN(new_n789));
  OAI21_X1  g588(.A(G120gat), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n783), .A2(new_n296), .A3(new_n604), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1341gat));
  OAI21_X1  g591(.A(G127gat), .B1(new_n788), .B2(new_n276), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n783), .A2(new_n302), .A3(new_n275), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(G1342gat));
  NAND3_X1  g594(.A1(new_n783), .A2(new_n305), .A3(new_n253), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT56), .Z(new_n797));
  OAI21_X1  g596(.A(G134gat), .B1(new_n788), .B2(new_n652), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1343gat));
  INV_X1    g598(.A(G141gat), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n774), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n765), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n764), .A2(new_n580), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n778), .A2(KEYINPUT115), .A3(new_n604), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n802), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n779), .B1(new_n807), .B2(new_n253), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n781), .B1(new_n808), .B2(new_n276), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT57), .B1(new_n809), .B2(new_n480), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n537), .A2(new_n608), .A3(new_n485), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n540), .C1(new_n780), .C2(new_n781), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n800), .B1(new_n814), .B2(new_n580), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n780), .A2(new_n781), .ZN(new_n816));
  INV_X1    g615(.A(new_n811), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n816), .A2(new_n480), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n800), .A3(new_n580), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT58), .B1(new_n820), .B2(KEYINPUT117), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(new_n822), .ZN(G1344gat));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n809), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n825), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n812), .B(new_n540), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT57), .B1(new_n816), .B2(new_n480), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n828), .A2(new_n604), .A3(new_n811), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n824), .B1(new_n830), .B2(G148gat), .ZN(new_n831));
  AOI211_X1 g630(.A(KEYINPUT59), .B(new_n596), .C1(new_n814), .C2(new_n604), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n537), .A2(new_n480), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(new_n604), .A3(new_n596), .A4(new_n484), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n831), .A2(new_n832), .B1(new_n782), .B2(new_n834), .ZN(G1345gat));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n275), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT119), .Z(new_n837));
  INV_X1    g636(.A(G155gat), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n276), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n837), .A2(new_n838), .B1(new_n814), .B2(new_n839), .ZN(G1346gat));
  INV_X1    g639(.A(G162gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n818), .A2(new_n841), .A3(new_n253), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n842), .B(KEYINPUT120), .Z(new_n843));
  AND2_X1   g642(.A1(new_n814), .A2(new_n253), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n841), .ZN(G1347gat));
  NAND2_X1  g644(.A1(new_n776), .A2(new_n779), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n276), .ZN(new_n847));
  INV_X1    g646(.A(new_n781), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n609), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT121), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n816), .B2(new_n609), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n533), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n540), .A2(new_n484), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n390), .A3(new_n580), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857));
  INV_X1    g656(.A(new_n719), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n849), .A2(new_n857), .A3(new_n858), .A4(new_n854), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n608), .B(new_n858), .C1(new_n780), .C2(new_n781), .ZN(new_n860));
  INV_X1    g659(.A(new_n854), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT122), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n863), .A2(new_n580), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n856), .B1(new_n390), .B2(new_n864), .ZN(G1348gat));
  NAND3_X1  g664(.A1(new_n853), .A2(new_n604), .A3(new_n854), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n406), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n391), .A2(new_n392), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n859), .A2(new_n862), .A3(new_n868), .A4(new_n604), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT123), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(KEYINPUT123), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n867), .A2(new_n870), .A3(KEYINPUT124), .A4(new_n871), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1349gat));
  AOI21_X1  g675(.A(new_n276), .B1(new_n379), .B2(new_n380), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n855), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n859), .A2(new_n862), .A3(new_n275), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n859), .A2(new_n862), .A3(KEYINPUT125), .A4(new_n275), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(G183gat), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT60), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n878), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1350gat));
  NAND4_X1  g687(.A1(new_n853), .A2(new_n374), .A3(new_n253), .A4(new_n854), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT126), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n859), .A2(new_n862), .A3(new_n253), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G190gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT61), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(KEYINPUT127), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(KEYINPUT127), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n891), .A2(new_n896), .A3(G190gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(KEYINPUT61), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n894), .A3(new_n898), .ZN(G1351gat));
  NAND2_X1  g698(.A1(new_n850), .A2(new_n852), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n485), .A3(new_n833), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n572), .A3(new_n580), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n828), .A2(new_n829), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n609), .A2(new_n484), .A3(new_n537), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n904), .A2(new_n580), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n572), .ZN(G1352gat));
  OR4_X1    g706(.A1(KEYINPUT62), .A2(new_n901), .A3(G204gat), .A4(new_n789), .ZN(new_n908));
  INV_X1    g707(.A(G204gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n902), .A2(new_n909), .A3(new_n604), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT62), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n904), .A2(new_n604), .A3(new_n905), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n908), .B(new_n911), .C1(new_n912), .C2(new_n909), .ZN(G1353gat));
  OR3_X1    g712(.A1(new_n901), .A2(G211gat), .A3(new_n276), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n828), .A2(new_n275), .A3(new_n829), .A4(new_n905), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n915), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT63), .B1(new_n915), .B2(G211gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1354gat));
  NAND3_X1  g717(.A1(new_n904), .A2(new_n253), .A3(new_n905), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G218gat), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n901), .A2(G218gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n652), .B2(new_n921), .ZN(G1355gat));
endmodule


