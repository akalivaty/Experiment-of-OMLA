//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n462), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n467), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G125), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n468), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(G136), .B2(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n470), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n469), .A2(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n487), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n492), .B1(new_n468), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(KEYINPUT66), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .A3(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(new_n506), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n499), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n501), .A2(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n513), .A2(G543), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT68), .B(G51), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n522), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n520), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n521), .A2(G90), .B1(new_n511), .B2(G52), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n501), .B2(new_n503), .ZN(new_n531));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(G651), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n529), .A2(KEYINPUT69), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT69), .B1(new_n529), .B2(new_n534), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n506), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n511), .A2(G43), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n514), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT70), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n511), .A2(G53), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n502), .A2(KEYINPUT5), .A3(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(G543), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(G91), .B2(new_n521), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n552), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND2_X1  g137(.A1(new_n521), .A2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n511), .A2(G49), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G288));
  AOI22_X1  g142(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n506), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n511), .A2(G48), .ZN(new_n570));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n514), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n521), .A2(G85), .B1(new_n511), .B2(G47), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT72), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(KEYINPUT71), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(KEYINPUT71), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(G651), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G66), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n556), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  INV_X1    g160(.A(G54), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n525), .B2(KEYINPUT73), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n511), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n521), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT10), .B1(new_n521), .B2(G92), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n585), .B(new_n590), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  MUX2_X1   g170(.A(new_n595), .B(G301), .S(G868), .Z(G321));
  XOR2_X1   g171(.A(G321), .B(KEYINPUT74), .Z(G284));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G299), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(G168), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(new_n598), .B2(G168), .ZN(G280));
  INV_X1    g176(.A(new_n595), .ZN(new_n602));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n468), .A2(new_n463), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n484), .A2(G135), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n469), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G123), .ZN(new_n618));
  OAI221_X1 g193(.A(new_n615), .B1(new_n616), .B2(new_n617), .C1(new_n481), .C2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G2096), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n613), .A2(new_n614), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT75), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT77), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2427), .B(G2430), .Z(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT78), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n630), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n638), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(G401));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(new_n612), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n645), .B2(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(new_n620), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT79), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT80), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT20), .Z(new_n662));
  OR2_X1    g237(.A1(new_n655), .A2(new_n657), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n660), .A3(new_n658), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n662), .B(new_n664), .C1(new_n660), .C2(new_n663), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT81), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT82), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G229));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G23), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n566), .B2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT86), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT33), .B(G1976), .Z(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(G6), .A2(G16), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n573), .B2(G16), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT32), .B(G1981), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n675), .A2(G22), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G166), .B2(new_n675), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(G1971), .Z(new_n688));
  AND4_X1   g263(.A1(new_n680), .A2(new_n684), .A3(new_n685), .A4(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G25), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT83), .Z(new_n694));
  OAI21_X1  g269(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n695));
  INV_X1    g270(.A(G107), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G2105), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT84), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n484), .A2(G131), .ZN(new_n700));
  INV_X1    g275(.A(G119), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n481), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n694), .B1(new_n703), .B2(G29), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  XOR2_X1   g280(.A(new_n704), .B(new_n705), .Z(new_n706));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(KEYINPUT87), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n691), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G24), .ZN(new_n710));
  XOR2_X1   g285(.A(G290), .B(KEYINPUT85), .Z(new_n711));
  AOI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n689), .A2(new_n690), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n709), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n707), .A2(KEYINPUT87), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G21), .ZN(new_n719));
  AOI21_X1  g294(.A(KEYINPUT92), .B1(new_n675), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(G168), .A2(G16), .ZN(new_n721));
  MUX2_X1   g296(.A(KEYINPUT92), .B(new_n720), .S(new_n721), .Z(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(G1966), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(new_n469), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT90), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(KEYINPUT90), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n484), .A2(G139), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n726), .A2(new_n727), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G33), .B(new_n731), .S(G29), .Z(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n722), .A2(G1966), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(G2072), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n723), .A2(new_n733), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G27), .A2(G29), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G164), .B2(G29), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT94), .B(G2078), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n692), .A2(G32), .ZN(new_n742));
  INV_X1    g317(.A(new_n481), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G129), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n484), .A2(G141), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n463), .A2(G105), .ZN(new_n746));
  AND3_X1   g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT91), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT26), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n742), .B1(new_n752), .B2(new_n692), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G34), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(KEYINPUT24), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(KEYINPUT24), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n692), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G160), .B2(new_n692), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G2084), .Z(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G11), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT30), .B(G28), .Z(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G29), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n619), .A2(new_n692), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(KEYINPUT93), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n761), .B(new_n766), .C1(KEYINPUT93), .C2(new_n765), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n755), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n675), .A2(G5), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G171), .B2(new_n675), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1961), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n736), .A2(new_n741), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT96), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n716), .A2(new_n717), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n692), .A2(G26), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT28), .Z(new_n776));
  AOI22_X1  g351(.A1(new_n743), .A2(G128), .B1(G140), .B2(new_n484), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(G116), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT88), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT89), .B(G2067), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n544), .A2(G16), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G16), .B2(G19), .ZN(new_n787));
  INV_X1    g362(.A(G1341), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G29), .A2(G35), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G162), .B2(G29), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT29), .B(G2090), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n787), .A2(new_n788), .ZN(new_n794));
  AND4_X1   g369(.A1(new_n785), .A2(new_n789), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n675), .A2(G20), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT23), .Z(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G299), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1956), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n675), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n602), .B2(new_n675), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n795), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n772), .B2(KEYINPUT96), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n718), .A2(new_n773), .A3(new_n774), .A4(new_n805), .ZN(G150));
  XOR2_X1   g381(.A(G150), .B(KEYINPUT97), .Z(G311));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n513), .B(G93), .C1(new_n554), .C2(new_n555), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n513), .A2(G55), .A3(G543), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n809), .A2(KEYINPUT98), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(G80), .A2(G543), .ZN(new_n816));
  INV_X1    g391(.A(G67), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n556), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G651), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n808), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n809), .A2(KEYINPUT98), .A3(new_n810), .ZN(new_n821));
  AOI21_X1  g396(.A(KEYINPUT98), .B1(new_n809), .B2(new_n810), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n819), .B(new_n808), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n820), .A2(new_n824), .B1(new_n540), .B2(new_n543), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT99), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n827), .A2(new_n544), .A3(new_n823), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n602), .A2(G559), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  AOI21_X1  g408(.A(G860), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n826), .A2(G860), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT100), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT101), .Z(G145));
  NAND2_X1  g415(.A1(new_n731), .A2(KEYINPUT102), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n751), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n703), .B(new_n610), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n782), .B(new_n497), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n743), .A2(G130), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n469), .A2(G118), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT103), .B1(new_n484), .B2(G142), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n484), .A2(KEYINPUT103), .A3(G142), .ZN(new_n850));
  OAI221_X1 g425(.A(new_n846), .B1(new_n847), .B2(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n845), .B(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n844), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n844), .A2(new_n852), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n477), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n484), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n619), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(G162), .Z(new_n860));
  AOI21_X1  g435(.A(G37), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n855), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g438(.A1(new_n826), .A2(new_n598), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n827), .A2(new_n544), .A3(new_n823), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n544), .B1(new_n827), .B2(new_n823), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n605), .ZN(new_n868));
  OR2_X1    g443(.A1(G299), .A2(new_n595), .ZN(new_n869));
  NAND2_X1  g444(.A1(G299), .A2(new_n595), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(KEYINPUT41), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  NOR2_X1   g447(.A1(G299), .A2(new_n595), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n591), .B(new_n592), .ZN(new_n874));
  AOI22_X1  g449(.A1(G651), .A2(new_n584), .B1(new_n587), .B2(new_n589), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n874), .A2(new_n875), .B1(new_n552), .B2(new_n559), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n872), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n868), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT105), .Z(new_n881));
  NOR2_X1   g456(.A1(new_n873), .A2(new_n876), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n868), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT104), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n887));
  INV_X1    g462(.A(new_n569), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n889));
  INV_X1    g464(.A(new_n572), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT106), .B1(new_n569), .B2(new_n572), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n891), .A2(G166), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(G166), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(G290), .A2(G288), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n576), .A2(new_n566), .A3(new_n580), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n887), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(KEYINPUT108), .A3(new_n895), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(new_n901), .B2(new_n895), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n899), .B(KEYINPUT107), .C1(new_n893), .C2(new_n894), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n886), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n864), .B1(new_n910), .B2(new_n598), .ZN(G295));
  OAI21_X1  g486(.A(new_n864), .B1(new_n910), .B2(new_n598), .ZN(G331));
  OAI21_X1  g487(.A(KEYINPUT110), .B1(new_n535), .B2(new_n536), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT69), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n504), .A2(G64), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n506), .B1(new_n915), .B2(new_n532), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n504), .A2(G90), .A3(new_n513), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n511), .A2(G52), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n914), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n529), .A2(KEYINPUT69), .A3(new_n534), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n913), .A2(G168), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(G168), .B1(new_n913), .B2(new_n923), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n828), .B(new_n825), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n913), .A2(G168), .A3(new_n923), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT110), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n921), .B1(new_n920), .B2(new_n922), .ZN(new_n929));
  OAI21_X1  g504(.A(G286), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n927), .B(new_n930), .C1(new_n865), .C2(new_n866), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n878), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n927), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT111), .B1(new_n867), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n924), .A2(new_n925), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n829), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n883), .B1(new_n867), .B2(new_n933), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT112), .B1(new_n940), .B2(new_n908), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n900), .A2(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n926), .A2(new_n882), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n934), .B2(new_n937), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n942), .B(new_n943), .C1(new_n945), .C2(new_n932), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n939), .A2(new_n931), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n936), .B1(new_n935), .B2(new_n829), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n926), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n948), .B1(new_n951), .B2(new_n879), .ZN(new_n952));
  AOI21_X1  g527(.A(G37), .B1(new_n952), .B2(new_n908), .ZN(new_n953));
  XOR2_X1   g528(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n878), .B1(new_n938), .B2(new_n926), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n942), .B1(new_n956), .B2(new_n948), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(new_n958), .B2(new_n954), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n952), .A2(new_n908), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n957), .A3(new_n964), .A4(new_n954), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT44), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n947), .A2(new_n953), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(KEYINPUT113), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n947), .A2(new_n953), .A3(new_n970), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n962), .B(new_n966), .C1(new_n969), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(KEYINPUT113), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(KEYINPUT43), .A3(new_n971), .ZN(new_n974));
  INV_X1    g549(.A(new_n966), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT114), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n961), .B1(new_n972), .B2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n497), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n980), .B2(new_n979), .ZN(new_n982));
  INV_X1    g557(.A(G40), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT116), .B1(new_n858), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  NAND3_X1  g560(.A1(G160), .A2(new_n985), .A3(G40), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n989), .A2(G1986), .A3(G290), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT48), .ZN(new_n991));
  INV_X1    g566(.A(G1996), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n751), .B(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G2067), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n782), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n703), .B(new_n705), .Z(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n991), .B1(new_n989), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n990), .A2(KEYINPUT48), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n988), .A2(new_n992), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n1002), .B(KEYINPUT46), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n995), .A2(new_n752), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n988), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT126), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  INV_X1    g583(.A(new_n703), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n705), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT125), .Z(new_n1011));
  OAI22_X1  g586(.A1(new_n1011), .A2(new_n996), .B1(G2067), .B2(new_n782), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1001), .B(new_n1008), .C1(new_n988), .C2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n858), .A2(KEYINPUT116), .A3(new_n983), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n985), .B1(G160), .B2(G40), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n979), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n497), .A2(new_n1023), .A3(new_n978), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1022), .A2(new_n984), .A3(new_n986), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1956), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(G299), .B(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1021), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1016), .A2(new_n1032), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1025), .A2(KEYINPUT121), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n802), .ZN(new_n1035));
  INV_X1    g610(.A(new_n979), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1016), .A2(new_n994), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n595), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1030), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1031), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(KEYINPUT60), .A3(new_n1037), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n595), .A2(KEYINPUT122), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n595), .A2(KEYINPUT122), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1035), .A2(KEYINPUT60), .A3(new_n1037), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1043), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1039), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n1031), .A3(KEYINPUT61), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1031), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n1039), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(G1996), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT58), .B(G1341), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n1016), .B2(new_n1036), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n544), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(KEYINPUT59), .B(new_n544), .C1(new_n1057), .C2(new_n1059), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1052), .A2(new_n1055), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1040), .B1(new_n1050), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1016), .A2(new_n1036), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n566), .A2(G1976), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(G8), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT52), .ZN(new_n1069));
  INV_X1    g644(.A(G1976), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT52), .B1(G288), .B2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1066), .A2(G8), .A3(new_n1067), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT49), .ZN(new_n1073));
  INV_X1    g648(.A(G1981), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n573), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n573), .A2(new_n1074), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1077), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(KEYINPUT49), .A3(new_n1075), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(new_n1080), .A3(new_n1066), .A4(G8), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1069), .A2(new_n1072), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G8), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT117), .B(G1971), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n1056), .A2(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1025), .A2(G2090), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G166), .A2(new_n1083), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(KEYINPUT55), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(G2090), .B1(new_n1025), .B2(KEYINPUT119), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(KEYINPUT119), .B2(new_n1025), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1083), .B1(new_n1092), .B2(new_n1085), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1082), .B(new_n1090), .C1(new_n1089), .C2(new_n1093), .ZN(new_n1094));
  AND4_X1   g669(.A1(new_n984), .A2(new_n1019), .A3(new_n986), .A4(new_n1017), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(G1966), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1025), .A2(G2084), .ZN(new_n1097));
  OAI21_X1  g672(.A(G286), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI221_X1 g673(.A(G168), .B1(new_n1025), .B2(G2084), .C1(new_n1095), .C2(G1966), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(G8), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT51), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1102), .A3(G8), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1094), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1056), .B2(G2078), .ZN(new_n1107));
  INV_X1    g682(.A(G1961), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1033), .A2(new_n1034), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G2078), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1095), .A2(KEYINPUT53), .A3(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1107), .A2(new_n1109), .A3(G301), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n858), .A2(new_n983), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1106), .A2(G2078), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n982), .A2(new_n1114), .A3(new_n1017), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1107), .A2(new_n1109), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1112), .A2(new_n1113), .B1(new_n1117), .B2(G171), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1105), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1117), .A2(G171), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1123), .A2(new_n1124), .A3(KEYINPUT54), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1065), .B(new_n1104), .C1(new_n1120), .C2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1082), .A2(new_n1089), .A3(new_n1087), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1066), .A2(G8), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n566), .A2(new_n1070), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT118), .Z(new_n1130));
  AOI21_X1  g705(.A(new_n1076), .B1(new_n1081), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1127), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  OAI211_X1 g708(.A(G8), .B(G168), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1094), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1136), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(new_n1090), .A3(new_n1082), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1132), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1126), .A2(KEYINPUT124), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT124), .B1(new_n1126), .B2(new_n1139), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1142), .A2(KEYINPUT62), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(KEYINPUT62), .ZN(new_n1144));
  NOR4_X1   g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n1122), .A4(new_n1094), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1140), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(G290), .B(new_n713), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n989), .B1(new_n998), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1013), .B1(new_n1146), .B2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g724(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1151));
  XNOR2_X1  g725(.A(new_n1151), .B(KEYINPUT127), .ZN(new_n1152));
  NOR2_X1   g726(.A1(G229), .A2(new_n1152), .ZN(new_n1153));
  AND3_X1   g727(.A1(new_n1153), .A2(new_n862), .A3(new_n959), .ZN(G308));
  NAND3_X1  g728(.A1(new_n1153), .A2(new_n862), .A3(new_n959), .ZN(G225));
endmodule


