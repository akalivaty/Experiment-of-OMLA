//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT72), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT78), .B(G469), .Z(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT73), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT73), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n195), .A2(G104), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n193), .A2(KEYINPUT73), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n199), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT74), .B1(new_n205), .B2(KEYINPUT3), .ZN(new_n206));
  AOI21_X1  g020(.A(G107), .B1(new_n194), .B2(new_n196), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT74), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n207), .A2(new_n208), .A3(new_n198), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n202), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT75), .A3(G101), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT75), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n208), .B1(new_n207), .B2(new_n198), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT73), .B(G104), .ZN(new_n214));
  OAI211_X1 g028(.A(KEYINPUT74), .B(KEYINPUT3), .C1(new_n214), .C2(G107), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n201), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(new_n216), .B2(new_n217), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n211), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n225), .A3(G143), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n222), .A2(G143), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(KEYINPUT65), .A3(new_n228), .A4(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT0), .B(G128), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n223), .A2(new_n225), .ZN(new_n236));
  INV_X1    g050(.A(G143), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(G146), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n235), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n216), .A2(new_n217), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(new_n219), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n221), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT11), .A3(G134), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G137), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n252));
  INV_X1    g066(.A(G131), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n249), .B2(G137), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n251), .A2(new_n252), .A3(new_n253), .A4(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n248), .A3(new_n253), .A4(new_n250), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n255), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n256), .A2(new_n258), .B1(new_n259), .B2(G131), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n217), .B(new_n202), .C1(new_n206), .C2(new_n209), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n193), .A2(G107), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n217), .B1(new_n205), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n226), .A2(new_n228), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n226), .A2(new_n228), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n240), .B2(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n261), .A2(new_n264), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT10), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n263), .B1(new_n216), .B2(new_n217), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n265), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n239), .B1(new_n236), .B2(new_n237), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n267), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(KEYINPUT10), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n246), .A2(new_n260), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G110), .B(G140), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G227), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n280), .B(new_n282), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n271), .B1(new_n276), .B2(new_n273), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n259), .A2(G131), .ZN(new_n287));
  INV_X1    g101(.A(new_n258), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT12), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT12), .B1(new_n286), .B2(new_n290), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n285), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n246), .A2(new_n278), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n290), .ZN(new_n300));
  AOI211_X1 g114(.A(KEYINPUT76), .B(new_n260), .C1(new_n246), .C2(new_n278), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n279), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n283), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n297), .B1(new_n303), .B2(KEYINPUT79), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT79), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n305), .A3(new_n283), .ZN(new_n306));
  AOI211_X1 g120(.A(G902), .B(new_n192), .C1(new_n304), .C2(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n279), .A2(new_n284), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n300), .B2(new_n301), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n279), .B1(new_n293), .B2(new_n295), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n283), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(G469), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n309), .B2(new_n311), .ZN(new_n317));
  INV_X1    g131(.A(G469), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT77), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n191), .B1(new_n307), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G214), .B1(G237), .B2(G902), .ZN(new_n322));
  NAND2_X1  g136(.A1(G234), .A2(G237), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(G952), .A3(new_n281), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT96), .Z(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT21), .B(G898), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(G902), .A3(G953), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n326), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G116), .B(G119), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n333), .A2(KEYINPUT67), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT2), .B(G113), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n334), .B(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n244), .B2(new_n219), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n221), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n340));
  INV_X1    g154(.A(G116), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n341), .A2(KEYINPUT5), .A3(G119), .ZN(new_n342));
  INV_X1    g156(.A(G113), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n340), .A2(new_n344), .B1(new_n336), .B2(new_n332), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n273), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G110), .B(G122), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n261), .A2(new_n264), .ZN(new_n351));
  INV_X1    g165(.A(new_n345), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n338), .B2(new_n221), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n348), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(KEYINPUT6), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G125), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n357), .B(new_n267), .C1(new_n274), .C2(new_n275), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n243), .B2(G125), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT80), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n241), .B1(new_n232), .B2(new_n233), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(new_n357), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n281), .A2(G224), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n366), .B(KEYINPUT81), .Z(new_n367));
  AND3_X1   g181(.A1(new_n362), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(new_n362), .B2(new_n365), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT6), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n347), .A2(new_n371), .A3(new_n349), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n356), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n351), .A2(new_n352), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n346), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n348), .B(KEYINPUT8), .Z(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT7), .B1(new_n366), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(new_n380), .B2(new_n366), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n365), .B(new_n382), .C1(new_n360), .C2(new_n363), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n377), .B1(new_n374), .B2(new_n346), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n366), .A2(KEYINPUT7), .ZN(new_n386));
  OAI22_X1  g200(.A1(new_n385), .A2(new_n376), .B1(new_n360), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(G902), .B1(new_n388), .B2(new_n355), .ZN(new_n389));
  OAI21_X1  g203(.A(G210), .B1(G237), .B2(G902), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n373), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n390), .B1(new_n373), .B2(new_n389), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n322), .B(new_n331), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT15), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G478), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n188), .A2(new_n397), .A3(G953), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(KEYINPUT94), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(KEYINPUT89), .A2(G122), .ZN(new_n401));
  NOR2_X1   g215(.A1(KEYINPUT89), .A2(G122), .ZN(new_n402));
  OAI21_X1  g216(.A(G116), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT90), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT90), .B(G116), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n341), .A2(G122), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n199), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G128), .B(G143), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(G134), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(KEYINPUT92), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n408), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n405), .A2(new_n406), .B1(KEYINPUT14), .B2(new_n408), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(KEYINPUT92), .ZN(new_n422));
  OAI21_X1  g236(.A(G107), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n421), .A2(KEYINPUT92), .B1(new_n418), .B2(new_n417), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n407), .A2(new_n415), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT92), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(KEYINPUT93), .A3(G107), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n414), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n411), .A2(KEYINPUT13), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n237), .A2(G128), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n433), .B(G134), .C1(KEYINPUT13), .C2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n435), .A2(KEYINPUT91), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n411), .A2(new_n249), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(KEYINPUT91), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n199), .B1(new_n407), .B2(new_n408), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n410), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n400), .B1(new_n432), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT93), .B1(new_n430), .B2(G107), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n424), .B(new_n199), .C1(new_n426), .C2(new_n429), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n413), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n442), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n399), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n448), .A3(new_n313), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT95), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n443), .A2(new_n448), .A3(KEYINPUT95), .A4(new_n313), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n396), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n449), .A2(new_n450), .B1(new_n395), .B2(G478), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  NOR2_X1   g269(.A1(G475), .A2(G902), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT88), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G125), .B(G140), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n223), .A3(new_n225), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n459), .A2(new_n222), .ZN(new_n461));
  NOR2_X1   g275(.A1(G237), .A2(G953), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G214), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n237), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(G143), .A3(G214), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(KEYINPUT18), .A2(G131), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n460), .A2(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT84), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n466), .A2(KEYINPUT84), .A3(new_n467), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n466), .A2(G131), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT17), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n464), .A2(new_n253), .A3(new_n465), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n459), .A2(KEYINPUT16), .ZN(new_n478));
  INV_X1    g292(.A(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G125), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(KEYINPUT16), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n222), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n478), .B(G146), .C1(KEYINPUT16), .C2(new_n480), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n466), .A2(KEYINPUT17), .A3(G131), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n477), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G113), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n193), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n473), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n473), .A2(new_n485), .A3(KEYINPUT87), .A4(new_n487), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n474), .A2(new_n476), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g308(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n459), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n459), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n498), .A2(new_n236), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(new_n483), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n493), .A2(KEYINPUT85), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n473), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n487), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n455), .B(new_n458), .C1(new_n492), .C2(new_n504), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n490), .A2(new_n491), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT20), .B1(new_n506), .B2(new_n457), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n487), .B1(new_n473), .B2(new_n485), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n490), .B2(new_n491), .ZN(new_n510));
  OAI21_X1  g324(.A(G475), .B1(new_n510), .B2(G902), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n453), .A2(new_n454), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n394), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n187), .B1(new_n321), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n316), .A2(new_n319), .ZN(new_n516));
  INV_X1    g330(.A(new_n279), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n299), .A2(new_n290), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT76), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n299), .A2(new_n298), .A3(new_n290), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT79), .B1(new_n521), .B2(new_n284), .ZN(new_n522));
  INV_X1    g336(.A(new_n297), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n306), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n192), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n313), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n190), .B1(new_n516), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n453), .A2(new_n454), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n393), .A2(new_n528), .A3(new_n512), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(KEYINPUT97), .A3(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n265), .A2(G119), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n531), .A2(KEYINPUT23), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n265), .A2(G119), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(KEYINPUT70), .A2(KEYINPUT23), .ZN(new_n536));
  OAI22_X1  g350(.A1(new_n532), .A2(new_n535), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n531), .A2(new_n533), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT24), .B(G110), .Z(new_n539));
  OAI22_X1  g353(.A1(new_n537), .A2(G110), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n483), .A3(new_n460), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n537), .A2(G110), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n482), .A2(new_n483), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT22), .B(G137), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n546), .B(new_n547), .Z(new_n548));
  XNOR2_X1  g362(.A(new_n545), .B(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n550));
  AOI21_X1  g364(.A(G902), .B1(new_n550), .B2(KEYINPUT71), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G234), .ZN(new_n555));
  OAI21_X1  g369(.A(G217), .B1(new_n555), .B2(G902), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n552), .B2(new_n553), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n549), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n313), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n462), .A2(G210), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT27), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT26), .B(G101), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n364), .A2(new_n290), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n256), .A2(new_n258), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n247), .A2(G134), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n250), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G131), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n276), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n566), .A2(new_n337), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n337), .B1(new_n566), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT28), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n256), .A2(new_n258), .B1(G131), .B2(new_n569), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n364), .A2(new_n290), .B1(new_n575), .B2(new_n276), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT28), .B1(new_n576), .B2(new_n337), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n565), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n337), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT30), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n566), .A2(new_n581), .A3(new_n571), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n566), .B2(new_n571), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n576), .A2(new_n337), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n565), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT31), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n571), .B1(new_n243), .B2(new_n260), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT30), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n576), .A2(new_n581), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n572), .B1(new_n592), .B2(new_n580), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(KEYINPUT31), .A3(new_n565), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n579), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(G472), .A2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT68), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n579), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT31), .B1(new_n593), .B2(new_n565), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n337), .B1(new_n590), .B2(new_n591), .ZN(new_n601));
  INV_X1    g415(.A(new_n565), .ZN(new_n602));
  NOR4_X1   g416(.A1(new_n601), .A2(new_n587), .A3(new_n572), .A4(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n599), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT68), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n596), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT32), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n598), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n588), .A2(new_n594), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n597), .B1(new_n609), .B2(new_n599), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT29), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n601), .A2(new_n572), .A3(new_n565), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n602), .B1(new_n574), .B2(new_n578), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT69), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n578), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n602), .A2(new_n611), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n589), .A2(new_n580), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n585), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n577), .B1(new_n619), .B2(KEYINPUT28), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n616), .B(new_n617), .C1(new_n620), .C2(new_n615), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n614), .A2(new_n313), .A3(new_n621), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n610), .A2(KEYINPUT32), .B1(new_n622), .B2(G472), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n561), .B1(new_n608), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n515), .A2(new_n530), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  OAI21_X1  g440(.A(G472), .B1(new_n595), .B2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n598), .A2(new_n627), .A3(new_n606), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n561), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n527), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n512), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n443), .A2(new_n448), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n443), .A2(new_n448), .A3(new_n632), .A4(KEYINPUT33), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(G478), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n449), .A2(new_n638), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n639), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n635), .B2(new_n636), .ZN(new_n645));
  INV_X1    g459(.A(new_n642), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT99), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n631), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n648), .A2(new_n394), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n630), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NAND2_X1  g466(.A1(new_n528), .A2(new_n631), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n393), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n527), .A2(new_n654), .A3(new_n629), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  INV_X1    g471(.A(new_n548), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n545), .B(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n313), .A3(new_n556), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n558), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n628), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n515), .A2(new_n530), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT100), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NAND2_X1  g482(.A1(new_n608), .A2(new_n623), .ZN(new_n669));
  INV_X1    g483(.A(new_n322), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n373), .A2(new_n389), .ZN(new_n671));
  INV_X1    g485(.A(new_n390), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n373), .A2(new_n389), .A3(new_n390), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n669), .A2(new_n675), .A3(new_n662), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n325), .B(KEYINPUT101), .Z(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(G900), .B2(new_n328), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n631), .B(new_n678), .C1(new_n453), .C2(new_n454), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n676), .A2(new_n527), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XNOR2_X1  g496(.A(new_n678), .B(KEYINPUT39), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n527), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n619), .A2(new_n602), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT103), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n586), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n313), .ZN(new_n689));
  AOI22_X1  g503(.A1(G472), .A2(new_n689), .B1(new_n610), .B2(KEYINPUT32), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n690), .A2(new_n691), .A3(new_n608), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n691), .B1(new_n690), .B2(new_n608), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n673), .A2(new_n674), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n512), .B1(new_n453), .B2(new_n454), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n662), .A2(new_n670), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n694), .A2(new_n697), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n685), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n237), .ZN(G45));
  INV_X1    g518(.A(new_n678), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n631), .B(new_n705), .C1(new_n643), .C2(new_n647), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n676), .A2(new_n527), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  AOI21_X1  g522(.A(new_n318), .B1(new_n524), .B2(new_n313), .ZN(new_n709));
  INV_X1    g523(.A(new_n189), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n307), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n649), .A2(new_n711), .A3(new_n624), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NAND3_X1  g528(.A1(new_n711), .A2(new_n624), .A3(new_n654), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  AND2_X1   g530(.A1(new_n513), .A2(new_n331), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n711), .A2(new_n676), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  OAI21_X1  g533(.A(new_n322), .B1(new_n391), .B2(new_n392), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n698), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n600), .A2(new_n603), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n574), .A2(new_n578), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT69), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n565), .B1(new_n724), .B2(new_n616), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n596), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n627), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n727), .A2(new_n561), .A3(new_n330), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n711), .A2(new_n721), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NOR2_X1   g544(.A1(new_n727), .A2(new_n663), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n711), .A2(new_n675), .A3(new_n706), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  OAI21_X1  g547(.A(new_n607), .B1(new_n595), .B2(new_n597), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n561), .B1(new_n623), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT106), .Z(new_n736));
  NAND4_X1  g550(.A1(new_n673), .A2(new_n189), .A3(new_n322), .A4(new_n674), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n314), .A2(G469), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n737), .B1(new_n526), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n643), .A2(new_n647), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n512), .A3(new_n678), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n736), .A2(new_n739), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n526), .A2(new_n738), .ZN(new_n745));
  INV_X1    g559(.A(new_n737), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n624), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n742), .B1(new_n747), .B2(new_n741), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(KEYINPUT105), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n706), .A2(new_n624), .A3(new_n739), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n751), .B2(new_n742), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n744), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  INV_X1    g568(.A(new_n747), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n679), .B(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NAND2_X1  g572(.A1(new_n740), .A2(new_n631), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n628), .A3(new_n662), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n312), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT45), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(G469), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n526), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n189), .A3(new_n683), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n391), .A2(new_n392), .A3(new_n670), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT108), .Z(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n764), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n763), .B2(new_n762), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  NAND4_X1  g594(.A1(new_n775), .A2(new_n608), .A3(new_n623), .A4(new_n561), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n773), .A2(new_n189), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n773), .A2(KEYINPUT47), .A3(new_n189), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n741), .B(new_n781), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n479), .ZN(G42));
  INV_X1    g601(.A(new_n677), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n761), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n711), .A2(new_n775), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n736), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT48), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT48), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n789), .A2(new_n793), .A3(new_n736), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n694), .A2(new_n561), .A3(new_n325), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n790), .ZN(new_n797));
  INV_X1    g611(.A(new_n648), .ZN(new_n798));
  OAI211_X1 g612(.A(G952), .B(new_n281), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n727), .A2(new_n561), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n761), .A2(new_n788), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n711), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n801), .A2(new_n720), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n795), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT115), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n795), .A2(new_n807), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n307), .A2(new_n709), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(new_n191), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n784), .A2(new_n785), .A3(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n812), .A2(new_n776), .ZN(new_n813));
  NOR2_X1   g627(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n697), .A2(new_n322), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n711), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(KEYINPUT114), .B2(KEYINPUT50), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n800), .B(new_n789), .C1(new_n813), .C2(new_n817), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n797), .A2(new_n512), .A3(new_n740), .ZN(new_n819));
  OAI211_X1 g633(.A(KEYINPUT114), .B(KEYINPUT50), .C1(new_n801), .C2(new_n816), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n789), .A2(new_n731), .A3(new_n790), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n818), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n818), .B2(new_n822), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n809), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n676), .B(new_n527), .C1(new_n706), .C2(new_n680), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n678), .A2(new_n189), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n720), .A2(new_n698), .A3(new_n662), .A4(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n831), .B(new_n745), .C1(new_n692), .C2(new_n693), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n732), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n732), .A2(new_n829), .A3(new_n832), .A4(KEYINPUT113), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n665), .B2(new_n655), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n648), .A2(KEYINPUT110), .A3(new_n394), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT110), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n798), .B2(new_n393), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n630), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n625), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n712), .A2(new_n715), .A3(new_n718), .A4(new_n729), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n748), .A2(KEYINPUT105), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n751), .A2(new_n750), .A3(new_n742), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n853), .B2(new_n744), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n665), .A2(new_n842), .A3(new_n655), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n512), .A2(new_n740), .A3(new_n678), .A4(new_n731), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n755), .A2(new_n756), .B1(new_n856), .B2(new_n739), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n663), .B1(new_n608), .B2(new_n623), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n453), .A2(new_n512), .A3(new_n454), .A4(new_n705), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n859), .A2(new_n775), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n527), .A2(new_n858), .A3(KEYINPUT112), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n669), .A2(new_n859), .A3(new_n775), .A4(new_n662), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n321), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n857), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n849), .A2(new_n854), .A3(new_n855), .A4(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n841), .A2(new_n867), .A3(KEYINPUT53), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n665), .A2(new_n655), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT111), .ZN(new_n871));
  INV_X1    g685(.A(new_n848), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n872), .A3(new_n855), .ZN(new_n873));
  INV_X1    g687(.A(new_n850), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n753), .A2(new_n866), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n836), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(new_n835), .B2(new_n836), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n869), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n868), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n836), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n839), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n869), .B1(new_n883), .B2(new_n867), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n857), .A2(KEYINPUT53), .A3(new_n865), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n753), .A3(new_n874), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n873), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n840), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n878), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT54), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n881), .A2(KEYINPUT54), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n809), .B(KEYINPUT116), .C1(new_n824), .C2(new_n825), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n828), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  NOR4_X1   g708(.A1(new_n759), .A2(new_n561), .A3(new_n190), .A4(new_n670), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT109), .Z(new_n896));
  XNOR2_X1  g710(.A(new_n810), .B(KEYINPUT49), .ZN(new_n897));
  OR4_X1    g711(.A1(new_n694), .A2(new_n896), .A3(new_n697), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(G75));
  OR2_X1    g713(.A1(new_n281), .A2(G952), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT118), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n887), .A2(new_n889), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n313), .B1(new_n884), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(G210), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n356), .A2(new_n372), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n370), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n902), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n904), .A2(KEYINPUT117), .A3(G210), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n911), .A2(new_n916), .ZN(G51));
  AOI21_X1  g731(.A(KEYINPUT53), .B1(new_n876), .B2(new_n879), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n849), .A2(new_n854), .A3(new_n855), .A4(new_n885), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n841), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n921), .A2(new_n313), .A3(new_n768), .ZN(new_n922));
  INV_X1    g736(.A(new_n524), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n841), .B2(new_n919), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n918), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT54), .B1(new_n918), .B2(new_n920), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n890), .A2(new_n884), .A3(KEYINPUT119), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n769), .B(KEYINPUT57), .Z(new_n931));
  AOI21_X1  g745(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n922), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n931), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT119), .B1(new_n890), .B2(new_n884), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n925), .B1(new_n884), .B2(new_n903), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n935), .B1(new_n938), .B2(new_n929), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT120), .B1(new_n939), .B2(new_n923), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n902), .B1(new_n934), .B2(new_n940), .ZN(G54));
  NAND2_X1  g755(.A1(KEYINPUT58), .A2(G475), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n904), .A2(new_n506), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n506), .B1(new_n904), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n901), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G60));
  XNOR2_X1  g762(.A(new_n637), .B(KEYINPUT122), .ZN(new_n949));
  NAND2_X1  g763(.A1(G478), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT59), .Z(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n902), .B1(new_n930), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n949), .B1(new_n891), .B2(new_n951), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(G63));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n959));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n921), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n959), .B1(new_n962), .B2(new_n660), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(KEYINPUT61), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n902), .B1(new_n962), .B2(new_n660), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n559), .B1(new_n921), .B2(new_n961), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n966), .B(new_n965), .C1(new_n963), .C2(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G66));
  INV_X1    g784(.A(new_n327), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n281), .B1(new_n971), .B2(G224), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n849), .A2(new_n855), .A3(new_n874), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(new_n281), .ZN(new_n974));
  INV_X1    g788(.A(G898), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n908), .B1(new_n975), .B2(G953), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n974), .B(new_n976), .ZN(G69));
  NAND2_X1  g791(.A1(G900), .A2(G953), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n732), .A2(new_n829), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n736), .A2(new_n721), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n757), .B1(new_n774), .B2(new_n980), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n786), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n779), .A2(new_n753), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n978), .B1(new_n983), .B2(G953), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n498), .B(KEYINPUT126), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT125), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n592), .B(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n703), .A2(new_n979), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n624), .A2(new_n775), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n991), .B(new_n684), .C1(new_n798), .C2(new_n653), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n786), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n989), .A2(new_n779), .A3(new_n990), .A4(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n987), .A2(G953), .ZN(new_n995));
  AOI22_X1  g809(.A1(new_n984), .A2(new_n987), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n994), .B2(new_n973), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n593), .A2(new_n602), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1000), .B1(new_n983), .B2(new_n973), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n612), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1003), .A2(new_n901), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n612), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n1000), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1008), .A2(new_n1002), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1006), .B1(new_n881), .B2(new_n1009), .ZN(G57));
endmodule


