

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  XOR2_X2 U323 ( .A(n344), .B(n343), .Z(n562) );
  XNOR2_X1 U324 ( .A(n334), .B(n333), .ZN(n338) );
  XNOR2_X1 U325 ( .A(n332), .B(KEYINPUT67), .ZN(n333) );
  NOR2_X1 U326 ( .A1(n571), .A2(n464), .ZN(n551) );
  XNOR2_X1 U327 ( .A(n327), .B(n326), .ZN(n523) );
  XOR2_X1 U328 ( .A(n368), .B(n330), .Z(n291) );
  XOR2_X1 U329 ( .A(n373), .B(n372), .Z(n292) );
  XOR2_X1 U330 ( .A(n368), .B(KEYINPUT75), .Z(n293) );
  XOR2_X1 U331 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n294) );
  INV_X1 U332 ( .A(KEYINPUT99), .ZN(n316) );
  NOR2_X1 U333 ( .A1(n523), .A2(n531), .ZN(n405) );
  XNOR2_X1 U334 ( .A(n402), .B(KEYINPUT114), .ZN(n403) );
  XNOR2_X1 U335 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U336 ( .A(n374), .B(n292), .ZN(n375) );
  XNOR2_X1 U337 ( .A(n404), .B(n403), .ZN(n531) );
  XNOR2_X1 U338 ( .A(n319), .B(n318), .ZN(n322) );
  XNOR2_X1 U339 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U340 ( .A(KEYINPUT65), .B(KEYINPUT41), .ZN(n394) );
  XNOR2_X1 U341 ( .A(n474), .B(KEYINPUT106), .ZN(n475) );
  XNOR2_X1 U342 ( .A(n477), .B(n394), .ZN(n454) );
  XNOR2_X1 U343 ( .A(n476), .B(n475), .ZN(n519) );
  XNOR2_X1 U344 ( .A(n484), .B(KEYINPUT58), .ZN(n485) );
  INV_X1 U345 ( .A(G43GAT), .ZN(n480) );
  XNOR2_X1 U346 ( .A(n486), .B(n485), .ZN(n488) );
  XNOR2_X1 U347 ( .A(n480), .B(KEYINPUT40), .ZN(n481) );
  XNOR2_X1 U348 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  XNOR2_X1 U349 ( .A(n482), .B(n481), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U351 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U353 ( .A(KEYINPUT19), .B(n297), .Z(n325) );
  XOR2_X1 U354 ( .A(G190GAT), .B(G134GAT), .Z(n330) );
  XOR2_X1 U355 ( .A(n330), .B(G99GAT), .Z(n300) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(G15GAT), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n298), .B(G113GAT), .ZN(n381) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(n381), .ZN(n299) );
  XNOR2_X1 U359 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n325), .B(n301), .ZN(n310) );
  XOR2_X1 U361 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n303) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U364 ( .A(n304), .B(KEYINPUT20), .Z(n308) );
  XNOR2_X1 U365 ( .A(G71GAT), .B(G176GAT), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n305), .B(G120GAT), .ZN(n371) );
  XNOR2_X1 U367 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n306), .B(KEYINPUT84), .ZN(n409) );
  XNOR2_X1 U369 ( .A(n371), .B(n409), .ZN(n307) );
  XNOR2_X1 U370 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n310), .B(n309), .ZN(n532) );
  XOR2_X1 U372 ( .A(KEYINPUT100), .B(G176GAT), .Z(n312) );
  XNOR2_X1 U373 ( .A(G169GAT), .B(G8GAT), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n312), .B(n311), .ZN(n324) );
  XOR2_X1 U375 ( .A(G204GAT), .B(G64GAT), .Z(n367) );
  XOR2_X1 U376 ( .A(G92GAT), .B(G218GAT), .Z(n314) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(G190GAT), .ZN(n313) );
  XNOR2_X1 U378 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U379 ( .A(n367), .B(n315), .Z(n319) );
  NAND2_X1 U380 ( .A1(G226GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n320), .B(G211GAT), .ZN(n444) );
  XNOR2_X1 U383 ( .A(n444), .B(KEYINPUT79), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n327) );
  INV_X1 U386 ( .A(n325), .ZN(n326) );
  XOR2_X1 U387 ( .A(G92GAT), .B(G85GAT), .Z(n329) );
  XNOR2_X1 U388 ( .A(G99GAT), .B(G106GAT), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n368) );
  NAND2_X1 U390 ( .A1(G232GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n291), .B(n331), .ZN(n334) );
  XOR2_X1 U392 ( .A(G218GAT), .B(G162GAT), .Z(n445) );
  XOR2_X1 U393 ( .A(n445), .B(KEYINPUT10), .Z(n332) );
  XOR2_X1 U394 ( .A(KEYINPUT68), .B(KEYINPUT11), .Z(n336) );
  XNOR2_X1 U395 ( .A(KEYINPUT77), .B(KEYINPUT9), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n344) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n339), .B(G29GAT), .ZN(n340) );
  XOR2_X1 U400 ( .A(n340), .B(KEYINPUT8), .Z(n342) );
  XNOR2_X1 U401 ( .A(G43GAT), .B(G50GAT), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n392) );
  INV_X1 U403 ( .A(n392), .ZN(n343) );
  XNOR2_X1 U404 ( .A(KEYINPUT78), .B(n562), .ZN(n483) );
  XNOR2_X1 U405 ( .A(KEYINPUT36), .B(n483), .ZN(n458) );
  XOR2_X1 U406 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n346) );
  XNOR2_X1 U407 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n352) );
  XOR2_X1 U409 ( .A(KEYINPUT13), .B(KEYINPUT73), .Z(n348) );
  XNOR2_X1 U410 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n370) );
  XOR2_X1 U412 ( .A(n370), .B(G78GAT), .Z(n350) );
  XOR2_X1 U413 ( .A(G8GAT), .B(G1GAT), .Z(n388) );
  XNOR2_X1 U414 ( .A(n388), .B(G211GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n365) );
  XOR2_X1 U417 ( .A(G155GAT), .B(G71GAT), .Z(n354) );
  XNOR2_X1 U418 ( .A(G22GAT), .B(G183GAT), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U420 ( .A(G64GAT), .B(KEYINPUT79), .Z(n356) );
  XNOR2_X1 U421 ( .A(G15GAT), .B(G127GAT), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U423 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U424 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n360) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U427 ( .A(KEYINPUT14), .B(n361), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n559) );
  NOR2_X1 U430 ( .A1(n458), .A2(n559), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n366), .B(KEYINPUT45), .ZN(n379) );
  XOR2_X1 U432 ( .A(G148GAT), .B(G78GAT), .Z(n442) );
  XNOR2_X1 U433 ( .A(n442), .B(n367), .ZN(n378) );
  NAND2_X1 U434 ( .A1(G230GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n293), .B(n369), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n374) );
  XOR2_X1 U437 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n373) );
  XNOR2_X1 U438 ( .A(KEYINPUT32), .B(KEYINPUT76), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n477) );
  NAND2_X1 U440 ( .A1(n379), .A2(n477), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n380), .B(KEYINPUT113), .ZN(n393) );
  XOR2_X1 U442 ( .A(n381), .B(KEYINPUT70), .Z(n383) );
  NAND2_X1 U443 ( .A1(G229GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U445 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n385) );
  XNOR2_X1 U446 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U448 ( .A(n387), .B(n386), .Z(n390) );
  XOR2_X1 U449 ( .A(G141GAT), .B(G22GAT), .Z(n439) );
  XNOR2_X1 U450 ( .A(n439), .B(n388), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U452 ( .A(n392), .B(n391), .Z(n552) );
  INV_X1 U453 ( .A(n552), .ZN(n573) );
  XOR2_X1 U454 ( .A(KEYINPUT72), .B(n573), .Z(n530) );
  NAND2_X1 U455 ( .A1(n393), .A2(n530), .ZN(n401) );
  INV_X1 U456 ( .A(n562), .ZN(n398) );
  NOR2_X1 U457 ( .A1(n552), .A2(n454), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n395), .B(n294), .ZN(n396) );
  NAND2_X1 U459 ( .A1(n396), .A2(n559), .ZN(n397) );
  NOR2_X1 U460 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U461 ( .A(KEYINPUT47), .B(n399), .ZN(n400) );
  NAND2_X1 U462 ( .A1(n401), .A2(n400), .ZN(n404) );
  XOR2_X1 U463 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n402) );
  XNOR2_X1 U464 ( .A(KEYINPUT54), .B(n405), .ZN(n431) );
  XOR2_X1 U465 ( .A(G85GAT), .B(G162GAT), .Z(n407) );
  XNOR2_X1 U466 ( .A(G29GAT), .B(G134GAT), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n430) );
  XOR2_X1 U469 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n411) );
  XNOR2_X1 U470 ( .A(G1GAT), .B(G57GAT), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U472 ( .A(G148GAT), .B(G120GAT), .Z(n413) );
  XNOR2_X1 U473 ( .A(G141GAT), .B(G113GAT), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n428) );
  XOR2_X1 U476 ( .A(KEYINPUT96), .B(KEYINPUT4), .Z(n417) );
  XNOR2_X1 U477 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U479 ( .A(KEYINPUT95), .B(n418), .Z(n420) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U482 ( .A(n421), .B(KEYINPUT97), .Z(n426) );
  XOR2_X1 U483 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n423) );
  XNOR2_X1 U484 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U486 ( .A(KEYINPUT3), .B(n424), .Z(n451) );
  XNOR2_X1 U487 ( .A(n451), .B(KEYINPUT94), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n549) );
  NAND2_X1 U491 ( .A1(n431), .A2(n549), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n432), .B(KEYINPUT66), .ZN(n572) );
  XOR2_X1 U493 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n434) );
  NAND2_X1 U494 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(KEYINPUT23), .B(n435), .ZN(n449) );
  XOR2_X1 U497 ( .A(G204GAT), .B(KEYINPUT22), .Z(n437) );
  XNOR2_X1 U498 ( .A(KEYINPUT93), .B(KEYINPUT91), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U500 ( .A(n438), .B(G106GAT), .Z(n441) );
  XNOR2_X1 U501 ( .A(G50GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U503 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(n466) );
  NOR2_X1 U508 ( .A1(n572), .A2(n466), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n452), .B(KEYINPUT55), .ZN(n453) );
  NOR2_X2 U510 ( .A1(n532), .A2(n453), .ZN(n568) );
  INV_X1 U511 ( .A(n454), .ZN(n537) );
  NAND2_X1 U512 ( .A1(n568), .A2(n537), .ZN(n457) );
  XOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(G176GAT), .ZN(n456) );
  BUF_X1 U515 ( .A(n458), .Z(n586) );
  XNOR2_X1 U516 ( .A(KEYINPUT88), .B(n532), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT27), .B(n523), .Z(n463) );
  XNOR2_X1 U518 ( .A(KEYINPUT28), .B(KEYINPUT69), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n459), .B(n466), .ZN(n527) );
  NAND2_X1 U520 ( .A1(n463), .A2(n527), .ZN(n460) );
  NOR2_X1 U521 ( .A1(n549), .A2(n460), .ZN(n534) );
  NAND2_X1 U522 ( .A1(n461), .A2(n534), .ZN(n472) );
  NAND2_X1 U523 ( .A1(n466), .A2(n532), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(KEYINPUT26), .ZN(n571) );
  INV_X1 U525 ( .A(n463), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n551), .B(KEYINPUT101), .ZN(n469) );
  NOR2_X1 U527 ( .A1(n532), .A2(n523), .ZN(n465) );
  NOR2_X1 U528 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U529 ( .A(KEYINPUT25), .B(n467), .ZN(n468) );
  NAND2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n549), .A2(n470), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n491) );
  NAND2_X1 U533 ( .A1(n559), .A2(n491), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n586), .A2(n473), .ZN(n476) );
  XNOR2_X1 U535 ( .A(KEYINPUT107), .B(KEYINPUT37), .ZN(n474) );
  INV_X1 U536 ( .A(n477), .ZN(n578) );
  NOR2_X1 U537 ( .A1(n530), .A2(n578), .ZN(n492) );
  NAND2_X1 U538 ( .A1(n519), .A2(n492), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(KEYINPUT108), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT38), .B(n479), .ZN(n507) );
  NOR2_X1 U541 ( .A1(n532), .A2(n507), .ZN(n482) );
  INV_X1 U542 ( .A(n483), .ZN(n543) );
  NAND2_X1 U543 ( .A1(n568), .A2(n543), .ZN(n486) );
  XOR2_X1 U544 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n484) );
  XOR2_X1 U545 ( .A(G190GAT), .B(KEYINPUT123), .Z(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(G1351GAT) );
  XNOR2_X1 U547 ( .A(KEYINPUT103), .B(KEYINPUT34), .ZN(n495) );
  INV_X1 U548 ( .A(n559), .ZN(n581) );
  NAND2_X1 U549 ( .A1(n483), .A2(n581), .ZN(n489) );
  XOR2_X1 U550 ( .A(KEYINPUT16), .B(n489), .Z(n490) );
  AND2_X1 U551 ( .A1(n491), .A2(n490), .ZN(n509) );
  NAND2_X1 U552 ( .A1(n492), .A2(n509), .ZN(n493) );
  XNOR2_X1 U553 ( .A(KEYINPUT102), .B(n493), .ZN(n501) );
  NOR2_X1 U554 ( .A1(n549), .A2(n501), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  NOR2_X1 U557 ( .A1(n501), .A2(n523), .ZN(n497) );
  XOR2_X1 U558 ( .A(G8GAT), .B(n497), .Z(G1325GAT) );
  XNOR2_X1 U559 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n532), .A2(n501), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G15GAT), .B(n500), .ZN(G1326GAT) );
  NOR2_X1 U563 ( .A1(n501), .A2(n527), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1327GAT) );
  NOR2_X1 U566 ( .A1(n549), .A2(n507), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n523), .A2(n507), .ZN(n506) );
  XOR2_X1 U570 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  NOR2_X1 U571 ( .A1(n527), .A2(n507), .ZN(n508) );
  XOR2_X1 U572 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  NOR2_X1 U573 ( .A1(n454), .A2(n573), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n509), .A2(n520), .ZN(n515) );
  NOR2_X1 U575 ( .A1(n549), .A2(n515), .ZN(n510) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n510), .Z(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n523), .A2(n515), .ZN(n512) );
  XOR2_X1 U579 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U580 ( .A1(n532), .A2(n515), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n527), .A2(n515), .ZN(n517) );
  XNOR2_X1 U584 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U588 ( .A1(n549), .A2(n526), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U591 ( .A1(n523), .A2(n526), .ZN(n524) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n532), .A2(n526), .ZN(n525) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  INV_X1 U598 ( .A(n530), .ZN(n565) );
  BUF_X1 U599 ( .A(n531), .Z(n548) );
  NOR2_X1 U600 ( .A1(n548), .A2(n532), .ZN(n533) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(KEYINPUT115), .B(n535), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n565), .A2(n544), .ZN(n536) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U606 ( .A1(n544), .A2(n537), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n541) );
  NAND2_X1 U609 ( .A1(n544), .A2(n581), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U613 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n552), .A2(n561), .ZN(n553) );
  XOR2_X1 U619 ( .A(KEYINPUT118), .B(n553), .Z(n554) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  NOR2_X1 U621 ( .A1(n561), .A2(n454), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n561), .ZN(n560) );
  XOR2_X1 U627 ( .A(G155GAT), .B(n560), .Z(G1346GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT120), .B(n563), .Z(n564) );
  XNOR2_X1 U630 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  XOR2_X1 U631 ( .A(G169GAT), .B(KEYINPUT121), .Z(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1348GAT) );
  NAND2_X1 U634 ( .A1(n581), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT122), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G183GAT), .B(n570), .ZN(G1350GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U638 ( .A1(n573), .A2(n584), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT127), .Z(n583) );
  NAND2_X1 U647 ( .A1(n584), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  INV_X1 U649 ( .A(n584), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

