

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U321 ( .A(n407), .B(KEYINPUT94), .ZN(n408) );
  XNOR2_X1 U322 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U323 ( .A(n390), .B(n389), .ZN(n394) );
  NOR2_X1 U324 ( .A1(n538), .A2(n466), .ZN(n583) );
  XOR2_X1 U325 ( .A(n406), .B(n405), .Z(n521) );
  AND2_X1 U326 ( .A1(G228GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U327 ( .A(G162GAT), .B(G50GAT), .Z(n433) );
  XNOR2_X1 U328 ( .A(n433), .B(n432), .ZN(n434) );
  INV_X1 U329 ( .A(KEYINPUT73), .ZN(n439) );
  XNOR2_X1 U330 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U331 ( .A(n388), .B(n289), .ZN(n389) );
  INV_X1 U332 ( .A(KEYINPUT96), .ZN(n421) );
  NOR2_X1 U333 ( .A1(n494), .A2(n465), .ZN(n552) );
  XNOR2_X1 U334 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U335 ( .A(n422), .B(n421), .ZN(n472) );
  XNOR2_X1 U336 ( .A(n409), .B(n408), .ZN(n538) );
  INV_X1 U337 ( .A(G218GAT), .ZN(n467) );
  XOR2_X1 U338 ( .A(KEYINPUT38), .B(n447), .Z(n490) );
  XNOR2_X1 U339 ( .A(n467), .B(KEYINPUT62), .ZN(n468) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n448) );
  XNOR2_X1 U341 ( .A(n469), .B(n468), .ZN(G1355GAT) );
  XNOR2_X1 U342 ( .A(n449), .B(n448), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n291) );
  XNOR2_X1 U344 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n290) );
  XNOR2_X1 U345 ( .A(n291), .B(n290), .ZN(n306) );
  XOR2_X1 U346 ( .A(G64GAT), .B(G204GAT), .Z(n369) );
  XOR2_X1 U347 ( .A(KEYINPUT33), .B(n369), .Z(n294) );
  XNOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT66), .ZN(n292) );
  XNOR2_X1 U349 ( .A(n292), .B(KEYINPUT13), .ZN(n327) );
  XNOR2_X1 U350 ( .A(n327), .B(G176GAT), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n299) );
  XNOR2_X1 U352 ( .A(G85GAT), .B(KEYINPUT70), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n295), .B(G92GAT), .ZN(n438) );
  XOR2_X1 U354 ( .A(n438), .B(KEYINPUT31), .Z(n297) );
  NAND2_X1 U355 ( .A1(G230GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U356 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U357 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U358 ( .A(KEYINPUT69), .B(G78GAT), .Z(n301) );
  XNOR2_X1 U359 ( .A(G148GAT), .B(G106GAT), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n388) );
  XNOR2_X1 U361 ( .A(G120GAT), .B(G99GAT), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n302), .B(G71GAT), .ZN(n396) );
  XNOR2_X1 U363 ( .A(n388), .B(n396), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U365 ( .A(n306), .B(n305), .Z(n579) );
  XOR2_X1 U366 ( .A(KEYINPUT64), .B(KEYINPUT29), .Z(n312) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n307), .B(KEYINPUT8), .ZN(n430) );
  XOR2_X1 U369 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n309) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(G169GAT), .ZN(n308) );
  XNOR2_X1 U371 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n430), .B(n310), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n317) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(G15GAT), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n313), .B(G8GAT), .ZN(n323) );
  XOR2_X1 U376 ( .A(n323), .B(G50GAT), .Z(n315) );
  NAND2_X1 U377 ( .A1(G229GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U378 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U379 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U380 ( .A(G197GAT), .B(G22GAT), .Z(n319) );
  XNOR2_X1 U381 ( .A(G141GAT), .B(G43GAT), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U383 ( .A(G36GAT), .B(n320), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n573) );
  NOR2_X1 U385 ( .A1(n579), .A2(n573), .ZN(n473) );
  XOR2_X1 U386 ( .A(G155GAT), .B(G22GAT), .Z(n383) );
  XOR2_X1 U387 ( .A(n323), .B(n383), .Z(n325) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U390 ( .A(n326), .B(KEYINPUT77), .Z(n329) );
  XNOR2_X1 U391 ( .A(n327), .B(KEYINPUT15), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U393 ( .A(G183GAT), .B(G71GAT), .Z(n331) );
  XNOR2_X1 U394 ( .A(G78GAT), .B(G211GAT), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U396 ( .A(n333), .B(n332), .Z(n341) );
  XOR2_X1 U397 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n335) );
  XNOR2_X1 U398 ( .A(KEYINPUT78), .B(KEYINPUT76), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U400 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n337) );
  XNOR2_X1 U401 ( .A(G127GAT), .B(G64GAT), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n582) );
  XOR2_X1 U405 ( .A(G113GAT), .B(G127GAT), .Z(n343) );
  XNOR2_X1 U406 ( .A(KEYINPUT81), .B(KEYINPUT0), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n397) );
  XOR2_X1 U408 ( .A(G29GAT), .B(n397), .Z(n345) );
  NAND2_X1 U409 ( .A1(G225GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U411 ( .A(G85GAT), .B(n346), .ZN(n363) );
  XOR2_X1 U412 ( .A(G1GAT), .B(KEYINPUT91), .Z(n348) );
  XNOR2_X1 U413 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n347) );
  XNOR2_X1 U414 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U415 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n350) );
  XNOR2_X1 U416 ( .A(G120GAT), .B(G57GAT), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U419 ( .A(G155GAT), .B(G148GAT), .Z(n354) );
  XNOR2_X1 U420 ( .A(G162GAT), .B(G134GAT), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U423 ( .A(n357), .B(KEYINPUT6), .Z(n361) );
  XOR2_X1 U424 ( .A(G141GAT), .B(KEYINPUT2), .Z(n359) );
  XNOR2_X1 U425 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n359), .B(n358), .ZN(n392) );
  XNOR2_X1 U427 ( .A(n392), .B(KEYINPUT1), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n494) );
  XOR2_X1 U430 ( .A(KEYINPUT86), .B(G197GAT), .Z(n365) );
  XNOR2_X1 U431 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U433 ( .A(G211GAT), .B(n366), .Z(n391) );
  XOR2_X1 U434 ( .A(G8GAT), .B(KEYINPUT93), .Z(n368) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U436 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U437 ( .A(n370), .B(n369), .Z(n372) );
  XOR2_X1 U438 ( .A(KEYINPUT75), .B(G36GAT), .Z(n431) );
  XNOR2_X1 U439 ( .A(G92GAT), .B(n431), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U441 ( .A(n391), .B(n373), .ZN(n380) );
  XOR2_X1 U442 ( .A(G169GAT), .B(G176GAT), .Z(n375) );
  XNOR2_X1 U443 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U445 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n377) );
  XNOR2_X1 U446 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n376) );
  XNOR2_X1 U447 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n395) );
  XOR2_X1 U449 ( .A(n380), .B(n395), .Z(n510) );
  XNOR2_X1 U450 ( .A(n510), .B(KEYINPUT27), .ZN(n417) );
  XOR2_X1 U451 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n382) );
  XNOR2_X1 U452 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n382), .B(n381), .ZN(n387) );
  XOR2_X1 U454 ( .A(KEYINPUT22), .B(G204GAT), .Z(n385) );
  XNOR2_X1 U455 ( .A(n433), .B(n383), .ZN(n384) );
  XNOR2_X1 U456 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U457 ( .A(n387), .B(n386), .Z(n390) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n553) );
  INV_X1 U460 ( .A(n395), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n404) );
  XOR2_X1 U462 ( .A(G134GAT), .B(G43GAT), .Z(n428) );
  XOR2_X1 U463 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n399) );
  XNOR2_X1 U464 ( .A(G15GAT), .B(KEYINPUT84), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U466 ( .A(n428), .B(n400), .Z(n402) );
  NAND2_X1 U467 ( .A1(G227GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U469 ( .A(n404), .B(n403), .ZN(n405) );
  INV_X1 U470 ( .A(n521), .ZN(n555) );
  NOR2_X1 U471 ( .A1(n553), .A2(n555), .ZN(n409) );
  INV_X1 U472 ( .A(KEYINPUT26), .ZN(n407) );
  NOR2_X1 U473 ( .A1(n417), .A2(n538), .ZN(n413) );
  INV_X1 U474 ( .A(n510), .ZN(n497) );
  NAND2_X1 U475 ( .A1(n497), .A2(n555), .ZN(n410) );
  NAND2_X1 U476 ( .A1(n553), .A2(n410), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n411), .B(KEYINPUT25), .ZN(n412) );
  NOR2_X1 U478 ( .A1(n413), .A2(n412), .ZN(n414) );
  NOR2_X1 U479 ( .A1(n494), .A2(n414), .ZN(n415) );
  XNOR2_X1 U480 ( .A(n415), .B(KEYINPUT95), .ZN(n420) );
  XOR2_X1 U481 ( .A(n553), .B(KEYINPUT28), .Z(n502) );
  XNOR2_X1 U482 ( .A(KEYINPUT85), .B(n521), .ZN(n416) );
  NOR2_X1 U483 ( .A1(n502), .A2(n416), .ZN(n418) );
  INV_X1 U484 ( .A(n494), .ZN(n508) );
  NOR2_X1 U485 ( .A1(n508), .A2(n417), .ZN(n520) );
  NAND2_X1 U486 ( .A1(n418), .A2(n520), .ZN(n419) );
  NAND2_X1 U487 ( .A1(n420), .A2(n419), .ZN(n422) );
  NOR2_X1 U488 ( .A1(n582), .A2(n472), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n423), .B(KEYINPUT101), .ZN(n445) );
  XOR2_X1 U490 ( .A(KEYINPUT74), .B(KEYINPUT72), .Z(n425) );
  XNOR2_X1 U491 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n444) );
  XOR2_X1 U493 ( .A(G106GAT), .B(G99GAT), .Z(n427) );
  XNOR2_X1 U494 ( .A(G218GAT), .B(G190GAT), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U496 ( .A(n429), .B(n428), .Z(n437) );
  XOR2_X1 U497 ( .A(n431), .B(n430), .Z(n435) );
  NAND2_X1 U498 ( .A1(G232GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n438), .B(KEYINPUT11), .ZN(n440) );
  XOR2_X1 U501 ( .A(n444), .B(n443), .Z(n569) );
  XNOR2_X1 U502 ( .A(KEYINPUT36), .B(n569), .ZN(n450) );
  NOR2_X1 U503 ( .A1(n445), .A2(n450), .ZN(n446) );
  XOR2_X1 U504 ( .A(KEYINPUT37), .B(n446), .Z(n507) );
  NAND2_X1 U505 ( .A1(n473), .A2(n507), .ZN(n447) );
  NAND2_X1 U506 ( .A1(n490), .A2(n555), .ZN(n449) );
  XOR2_X1 U507 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n464) );
  INV_X1 U508 ( .A(n582), .ZN(n565) );
  NOR2_X1 U509 ( .A1(n450), .A2(n565), .ZN(n452) );
  XNOR2_X1 U510 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n579), .A2(n453), .ZN(n454) );
  NAND2_X1 U513 ( .A1(n454), .A2(n573), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n579), .B(KEYINPUT41), .ZN(n559) );
  NOR2_X1 U515 ( .A1(n573), .A2(n559), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n455), .B(KEYINPUT46), .ZN(n456) );
  NOR2_X1 U517 ( .A1(n582), .A2(n456), .ZN(n457) );
  NAND2_X1 U518 ( .A1(n457), .A2(n569), .ZN(n459) );
  XOR2_X1 U519 ( .A(KEYINPUT47), .B(KEYINPUT110), .Z(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U522 ( .A(KEYINPUT48), .B(n462), .ZN(n519) );
  NAND2_X1 U523 ( .A1(n519), .A2(n497), .ZN(n463) );
  XOR2_X1 U524 ( .A(n464), .B(n463), .Z(n465) );
  INV_X1 U525 ( .A(n552), .ZN(n466) );
  INV_X1 U526 ( .A(n583), .ZN(n572) );
  NOR2_X1 U527 ( .A1(n450), .A2(n572), .ZN(n469) );
  INV_X1 U528 ( .A(n569), .ZN(n548) );
  NOR2_X1 U529 ( .A1(n548), .A2(n565), .ZN(n470) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  NOR2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n492) );
  NAND2_X1 U532 ( .A1(n473), .A2(n492), .ZN(n482) );
  NOR2_X1 U533 ( .A1(n508), .A2(n482), .ZN(n474) );
  XOR2_X1 U534 ( .A(G1GAT), .B(n474), .Z(n475) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(n475), .ZN(G1324GAT) );
  NOR2_X1 U536 ( .A1(n510), .A2(n482), .ZN(n477) );
  XNOR2_X1 U537 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(G1325GAT) );
  NOR2_X1 U539 ( .A1(n482), .A2(n521), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n479) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  INV_X1 U544 ( .A(n502), .ZN(n523) );
  NOR2_X1 U545 ( .A1(n523), .A2(n482), .ZN(n483) );
  XOR2_X1 U546 ( .A(G22GAT), .B(n483), .Z(G1327GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n485) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U550 ( .A(KEYINPUT100), .B(n486), .Z(n488) );
  NAND2_X1 U551 ( .A1(n494), .A2(n490), .ZN(n487) );
  XNOR2_X1 U552 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n490), .A2(n497), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n489), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n490), .A2(n502), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n491), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U557 ( .A(n573), .ZN(n539) );
  NOR2_X1 U558 ( .A1(n539), .A2(n559), .ZN(n506) );
  NAND2_X1 U559 ( .A1(n506), .A2(n492), .ZN(n493) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(n493), .Z(n501) );
  NAND2_X1 U561 ( .A1(n501), .A2(n494), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n495), .B(KEYINPUT42), .ZN(n496) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(n496), .ZN(G1332GAT) );
  XOR2_X1 U564 ( .A(G64GAT), .B(KEYINPUT105), .Z(n499) );
  NAND2_X1 U565 ( .A1(n501), .A2(n497), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n499), .B(n498), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n501), .A2(n555), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n500), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n504) );
  NAND2_X1 U570 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(n505), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n507), .A2(n506), .ZN(n515) );
  NOR2_X1 U574 ( .A1(n508), .A2(n515), .ZN(n509) );
  XOR2_X1 U575 ( .A(G85GAT), .B(n509), .Z(G1336GAT) );
  NOR2_X1 U576 ( .A1(n510), .A2(n515), .ZN(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G92GAT), .B(n513), .ZN(G1337GAT) );
  NOR2_X1 U580 ( .A1(n521), .A2(n515), .ZN(n514) );
  XOR2_X1 U581 ( .A(G99GAT), .B(n514), .Z(G1338GAT) );
  NOR2_X1 U582 ( .A1(n523), .A2(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n518), .ZN(G1339GAT) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n537) );
  NOR2_X1 U588 ( .A1(n521), .A2(n537), .ZN(n522) );
  XNOR2_X1 U589 ( .A(KEYINPUT112), .B(n522), .ZN(n524) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT113), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n533), .A2(n539), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n529) );
  INV_X1 U595 ( .A(n559), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n533), .A2(n543), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U598 ( .A(G120GAT), .B(n530), .Z(G1341GAT) );
  NAND2_X1 U599 ( .A1(n533), .A2(n582), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n531), .B(KEYINPUT50), .ZN(n532) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n535) );
  NAND2_X1 U603 ( .A1(n533), .A2(n548), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n536), .ZN(G1343GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n541) );
  NOR2_X1 U607 ( .A1(n538), .A2(n537), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n549), .A2(n539), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  NAND2_X1 U612 ( .A1(n549), .A2(n543), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n549), .A2(n582), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n547), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U617 ( .A(G162GAT), .B(KEYINPUT119), .Z(n551) );
  NAND2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT55), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n568) );
  NOR2_X1 U623 ( .A1(n573), .A2(n568), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n568), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(KEYINPUT122), .B(n562), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n568), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT124), .B(n566), .Z(n567) );
  XNOR2_X1 U634 ( .A(G183GAT), .B(n567), .ZN(G1350GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT58), .B(n570), .Z(n571) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(n571), .ZN(G1351GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(KEYINPUT59), .B(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U645 ( .A1(n583), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
endmodule

