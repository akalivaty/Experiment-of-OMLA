//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT67), .B(G128), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n193), .B1(G143), .B2(new_n187), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n193), .A3(G128), .ZN(new_n197));
  XOR2_X1   g011(.A(G134), .B(G137), .Z(new_n198));
  AOI22_X1  g012(.A1(new_n195), .A2(new_n197), .B1(G131), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  OAI22_X1  g016(.A1(KEYINPUT65), .A2(new_n201), .B1(new_n202), .B2(G134), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI22_X1  g019(.A1(new_n204), .A2(KEYINPUT11), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT65), .A4(G134), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n203), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n200), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n207), .ZN(new_n211));
  AOI22_X1  g025(.A1(new_n204), .A2(KEYINPUT11), .B1(new_n205), .B2(G137), .ZN(new_n212));
  AND4_X1   g026(.A1(new_n200), .A2(new_n211), .A3(new_n209), .A4(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n199), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G116), .B(G119), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(KEYINPUT2), .B(G113), .Z(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n215), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(KEYINPUT68), .A3(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND4_X1   g038(.A1(KEYINPUT65), .A2(new_n201), .A3(new_n202), .A4(G134), .ZN(new_n225));
  AOI22_X1  g039(.A1(KEYINPUT65), .A2(new_n201), .B1(new_n202), .B2(G134), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n209), .B(new_n212), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n211), .A2(new_n200), .A3(new_n209), .A4(new_n212), .ZN(new_n229));
  INV_X1    g043(.A(new_n208), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n228), .A2(new_n229), .B1(G131), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(KEYINPUT0), .B(G128), .Z(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT64), .A3(new_n191), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  OAI211_X1 g048(.A(KEYINPUT0), .B(G128), .C1(new_n196), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n214), .B(new_n224), .C1(new_n231), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT28), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n240));
  NOR2_X1   g054(.A1(G237), .A2(G953), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G210), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n240), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G101), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n239), .A2(KEYINPUT29), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n237), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n230), .A2(G131), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n210), .B2(new_n213), .ZN(new_n251));
  INV_X1    g065(.A(new_n236), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n253), .A2(KEYINPUT69), .A3(new_n214), .A4(new_n224), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT72), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n222), .A2(new_n223), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n228), .A2(new_n229), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n236), .B1(new_n258), .B2(new_n250), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n198), .A2(G131), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT67), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n265), .A2(new_n266), .B1(new_n188), .B2(new_n190), .ZN(new_n267));
  AND4_X1   g081(.A1(new_n193), .A2(new_n188), .A3(new_n190), .A4(G128), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n260), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n229), .B2(new_n228), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n257), .B1(new_n259), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n249), .A2(new_n254), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n256), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n247), .B1(new_n274), .B2(KEYINPUT28), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT73), .B1(new_n275), .B2(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n271), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n272), .B1(new_n249), .B2(new_n254), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT28), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n247), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n238), .B1(new_n249), .B2(new_n254), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n239), .A2(new_n271), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(new_n245), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT30), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n253), .B2(new_n214), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n259), .A2(KEYINPUT30), .A3(new_n270), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n257), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n294), .A2(new_n246), .A3(new_n255), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n285), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n276), .A2(new_n284), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G472), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n249), .A2(new_n254), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n293), .A3(new_n246), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT31), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n245), .B1(new_n286), .B2(new_n287), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n299), .A2(new_n293), .A3(new_n303), .A4(new_n246), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT32), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT71), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(KEYINPUT71), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n298), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n305), .A2(new_n306), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT32), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT71), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n306), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n310), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n298), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n314), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G217), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(G234), .B2(new_n283), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n330));
  OR3_X1    g144(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G146), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n327), .A2(new_n329), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n187), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n261), .A2(G119), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n192), .B2(G119), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT24), .B(G110), .Z(new_n338));
  OR2_X1    g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT23), .B1(new_n261), .B2(G119), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(new_n336), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI22_X1  g157(.A1(new_n339), .A2(KEYINPUT77), .B1(G110), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n339), .A2(KEYINPUT77), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n335), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n330), .A2(new_n331), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n187), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n330), .A2(new_n331), .A3(new_n350), .A4(G146), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n343), .A2(G110), .B1(new_n337), .B2(new_n338), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n352), .B2(new_n353), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n346), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G953), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(G221), .A3(G234), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT78), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT22), .B(G137), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n346), .B(new_n362), .C1(new_n355), .C2(new_n356), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT25), .B1(new_n366), .B2(new_n283), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  AOI211_X1 g182(.A(new_n368), .B(G902), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n325), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(KEYINPUT79), .B(new_n325), .C1(new_n367), .C2(new_n369), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n325), .A2(G902), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT80), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT81), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n372), .A2(new_n379), .A3(new_n373), .A4(new_n376), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT3), .B1(new_n383), .B2(G107), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G104), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G101), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n382), .B1(new_n390), .B2(KEYINPUT4), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n389), .A2(KEYINPUT83), .A3(new_n392), .A4(G101), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT82), .B(G101), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n390), .B(KEYINPUT4), .C1(new_n395), .C2(new_n389), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n386), .A2(G104), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n388), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n389), .B2(new_n395), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n215), .A2(KEYINPUT5), .ZN(new_n403));
  INV_X1    g217(.A(G116), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n404), .A2(KEYINPUT5), .A3(G119), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(G113), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n220), .ZN(new_n407));
  OAI22_X1  g221(.A1(new_n397), .A2(new_n224), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(G110), .B(G122), .Z(new_n409));
  OR2_X1    g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n409), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT90), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n410), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n267), .A2(new_n268), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n328), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n236), .A2(G125), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G224), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(G953), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n408), .B(new_n409), .C1(new_n412), .C2(new_n413), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n415), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT7), .B1(new_n420), .B2(G953), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n419), .B(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n407), .A2(new_n402), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n427), .A2(KEYINPUT92), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n407), .A2(new_n402), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(KEYINPUT92), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT91), .B(KEYINPUT8), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n409), .B(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n426), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(G902), .B1(new_n434), .B2(new_n410), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n424), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G210), .B1(G237), .B2(G902), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n424), .A2(new_n435), .A3(new_n437), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(KEYINPUT93), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n440), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT93), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n446), .B(KEYINPUT89), .Z(new_n447));
  NOR2_X1   g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n416), .A2(new_n402), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n451));
  INV_X1    g265(.A(new_n395), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n400), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n191), .B1(new_n194), .B2(new_n261), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n197), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n251), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT12), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n449), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n459), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n457), .A2(new_n251), .A3(KEYINPUT85), .A4(KEYINPUT12), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G140), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n358), .A2(G227), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n394), .A2(new_n252), .A3(new_n396), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT10), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n195), .B2(new_n197), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n456), .A2(new_n471), .B1(new_n453), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n473), .A3(new_n231), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n470), .A2(new_n473), .A3(KEYINPUT84), .A4(new_n231), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT87), .A4(new_n462), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n465), .A2(new_n469), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n470), .A2(new_n473), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n251), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT88), .A3(new_n468), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n476), .A2(new_n477), .B1(new_n251), .B2(new_n481), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n486), .B2(new_n469), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n480), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n283), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n478), .A2(new_n463), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n478), .B2(new_n463), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n468), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n478), .A2(new_n469), .A3(new_n482), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(G469), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(G469), .A2(G902), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT9), .B(G234), .ZN(new_n499));
  OAI21_X1  g313(.A(G221), .B1(new_n499), .B2(G902), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n261), .A2(G143), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT95), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n192), .A2(G143), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n503), .A2(new_n504), .ZN(new_n508));
  OAI21_X1  g322(.A(G134), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n503), .A2(new_n205), .A3(new_n506), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT96), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n404), .A2(G122), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n404), .A2(G122), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n386), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n514), .ZN(new_n516));
  OAI21_X1  g330(.A(G107), .B1(new_n516), .B2(new_n512), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n510), .A2(new_n511), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n509), .B(new_n518), .C1(new_n511), .C2(new_n510), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n520));
  INV_X1    g334(.A(new_n515), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n205), .B1(new_n503), .B2(new_n506), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n523), .B2(new_n510), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n514), .A2(KEYINPUT14), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT97), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n512), .B1(new_n516), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n386), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n520), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n510), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n515), .B1(new_n532), .B2(new_n522), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n533), .A2(KEYINPUT98), .A3(new_n529), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n519), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n499), .A2(new_n324), .A3(G953), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n519), .B(new_n536), .C1(new_n534), .C2(new_n531), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n283), .ZN(new_n541));
  INV_X1    g355(.A(G478), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(G902), .B1(new_n538), .B2(new_n539), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(KEYINPUT15), .B2(new_n542), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n241), .A2(G214), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(G143), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT18), .A2(G131), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n333), .B2(new_n187), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n333), .A2(new_n187), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n333), .A2(new_n552), .A3(new_n187), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n549), .A2(new_n209), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT17), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n549), .B(new_n209), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(KEYINPUT17), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n558), .B1(new_n562), .B2(new_n352), .ZN(new_n563));
  XNOR2_X1  g377(.A(G113), .B(G122), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(new_n383), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n558), .B(new_n565), .C1(new_n562), .C2(new_n352), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n283), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G475), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n333), .B(KEYINPUT19), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n187), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n561), .A2(new_n332), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n551), .A2(new_n557), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n568), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT20), .ZN(new_n578));
  NOR2_X1   g392(.A1(G475), .A2(G902), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n577), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n571), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(G234), .A2(G237), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(G952), .A3(new_n358), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(G902), .A3(G953), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT21), .B(G898), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n547), .A2(new_n583), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n448), .A2(new_n501), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n323), .A2(new_n381), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n395), .ZN(G3));
  NAND2_X1  g408(.A1(new_n305), .A2(new_n283), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n315), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n501), .A2(new_n598), .A3(new_n378), .A4(new_n380), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n447), .B1(new_n439), .B2(new_n440), .ZN(new_n600));
  INV_X1    g414(.A(new_n590), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n540), .A2(KEYINPUT33), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n538), .A2(new_n604), .A3(new_n539), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(G478), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n542), .A2(new_n283), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n545), .B2(new_n542), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n583), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  OR3_X1    g423(.A1(new_n602), .A2(KEYINPUT99), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT99), .B1(new_n602), .B2(new_n609), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n599), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT34), .B(G104), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  INV_X1    g428(.A(new_n547), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n581), .A2(KEYINPUT100), .ZN(new_n616));
  INV_X1    g430(.A(new_n582), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n580), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n616), .B(new_n571), .C1(new_n618), .C2(KEYINPUT100), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(new_n601), .A3(new_n600), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n599), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT35), .B(G107), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NOR2_X1   g438(.A1(new_n362), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n357), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n375), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n372), .A2(new_n373), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n591), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n501), .A3(new_n448), .A4(new_n598), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  NAND2_X1  g446(.A1(new_n501), .A2(new_n628), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n585), .B(KEYINPUT101), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n637), .B2(new_n588), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n620), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n600), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI221_X4 g456(.A(new_n313), .B1(new_n297), .B2(G472), .C1(new_n320), .C2(new_n310), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT74), .B1(new_n321), .B2(new_n298), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n634), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  XOR2_X1   g460(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n638), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n501), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT40), .Z(new_n650));
  AOI21_X1  g464(.A(new_n245), .B1(new_n299), .B2(new_n293), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n652), .B(new_n283), .C1(new_n246), .C2(new_n274), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n320), .A2(new_n310), .B1(G472), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n547), .A2(new_n583), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n445), .B(KEYINPUT38), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n657), .A2(new_n447), .A3(new_n628), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n650), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  NOR2_X1   g474(.A1(new_n609), .A2(new_n638), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n641), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n634), .B(new_n663), .C1(new_n643), .C2(new_n644), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n323), .A2(KEYINPUT103), .A3(new_n634), .A4(new_n663), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  NAND2_X1  g483(.A1(new_n488), .A2(new_n283), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G469), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n500), .A3(new_n490), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n610), .B2(new_n611), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n323), .A2(new_n381), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT41), .B(G113), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G15));
  NOR2_X1   g490(.A1(new_n621), .A2(new_n672), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n323), .A2(new_n381), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  NOR2_X1   g493(.A1(new_n672), .A2(new_n641), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(new_n629), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n323), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G119), .ZN(G21));
  NOR4_X1   g497(.A1(new_n672), .A2(new_n641), .A3(new_n590), .A4(new_n655), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n377), .A2(KEYINPUT105), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n372), .A2(new_n686), .A3(new_n373), .A4(new_n376), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n306), .B(KEYINPUT104), .Z(new_n690));
  AOI21_X1  g504(.A(new_n246), .B1(new_n279), .B2(new_n239), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n301), .A2(new_n304), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n596), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n688), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n689), .B1(new_n688), .B2(new_n694), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n684), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  AND2_X1   g512(.A1(new_n694), .A2(new_n628), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n661), .A3(new_n680), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G125), .ZN(G27));
  NAND3_X1  g515(.A1(new_n298), .A2(new_n317), .A3(new_n319), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n688), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n498), .A2(KEYINPUT107), .A3(new_n500), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n498), .B2(new_n500), .ZN(new_n707));
  INV_X1    g521(.A(new_n447), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n445), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n710), .A2(new_n661), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n705), .A2(KEYINPUT42), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n710), .B(new_n381), .C1(new_n643), .C2(new_n644), .ZN(new_n714));
  OAI211_X1 g528(.A(KEYINPUT108), .B(new_n713), .C1(new_n714), .C2(new_n662), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n323), .A2(new_n381), .A3(new_n661), .A4(new_n710), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT108), .B1(new_n717), .B2(new_n713), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n712), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  OR2_X1    g534(.A1(new_n714), .A2(new_n640), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  AOI22_X1  g536(.A1(new_n617), .A2(new_n580), .B1(new_n570), .B2(G475), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n606), .A3(new_n608), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT43), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT43), .B1(new_n724), .B2(new_n725), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n597), .A3(new_n628), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n500), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n494), .A2(new_n495), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n489), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n734), .B2(new_n733), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT46), .B1(new_n736), .B2(new_n497), .ZN(new_n737));
  INV_X1    g551(.A(new_n490), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n497), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n732), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n709), .B1(new_n729), .B2(new_n730), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n731), .A2(new_n741), .A3(new_n742), .A4(new_n648), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G137), .ZN(G39));
  NOR4_X1   g558(.A1(new_n323), .A2(new_n381), .A3(new_n662), .A4(new_n709), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n741), .A2(KEYINPUT47), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n747), .B(new_n732), .C1(new_n739), .C2(new_n740), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G140), .ZN(G42));
  NOR3_X1   g564(.A1(new_n726), .A2(new_n727), .A3(new_n635), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT113), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n709), .A2(new_n672), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n705), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT48), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n381), .A2(new_n753), .A3(new_n654), .A4(new_n586), .ZN(new_n757));
  OAI211_X1 g571(.A(G952), .B(new_n358), .C1(new_n757), .C2(new_n609), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n695), .A2(new_n696), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n759), .A2(new_n752), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n758), .B1(new_n760), .B2(new_n680), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n709), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n746), .A2(new_n748), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT114), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n671), .A2(new_n490), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n500), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT115), .Z(new_n769));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n764), .A2(KEYINPUT114), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n763), .B(new_n760), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n447), .A2(new_n657), .A3(new_n500), .A4(new_n766), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n759), .A2(new_n752), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT50), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n754), .A2(new_n699), .ZN(new_n776));
  INV_X1    g590(.A(new_n757), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n583), .B1(new_n606), .B2(new_n608), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n772), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n762), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n763), .B(new_n760), .C1(new_n764), .C2(new_n768), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT116), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n781), .A2(new_n788), .A3(KEYINPUT51), .A4(new_n785), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT117), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n645), .A2(new_n700), .ZN(new_n793));
  INV_X1    g607(.A(new_n501), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n628), .A2(new_n638), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(KEYINPUT112), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n794), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n600), .B(new_n656), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n633), .B1(new_n314), .B2(new_n322), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT103), .B1(new_n801), .B2(new_n663), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n664), .A2(new_n665), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n793), .B(new_n800), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n609), .B1(new_n615), .B2(new_n583), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n448), .A2(new_n601), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n630), .B1(new_n599), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n323), .B2(new_n681), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n323), .B(new_n381), .C1(new_n673), .C2(new_n592), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n678), .A4(new_n697), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n711), .A2(new_n699), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n615), .A2(new_n639), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n709), .A2(new_n619), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n801), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n812), .B(new_n816), .C1(new_n640), .C2(new_n714), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n668), .A2(new_n819), .A3(new_n793), .A4(new_n800), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n805), .A2(new_n719), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n645), .A2(new_n700), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT52), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n822), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n823), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT54), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n825), .A2(KEYINPUT53), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n823), .B(new_n830), .C1(new_n821), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n784), .A2(new_n833), .A3(new_n790), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n792), .A2(new_n829), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(G952), .B2(G953), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n767), .A2(KEYINPUT49), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n724), .A2(new_n447), .A3(new_n732), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n688), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT111), .Z(new_n840));
  OR2_X1    g654(.A1(new_n767), .A2(KEYINPUT49), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n654), .A3(new_n657), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(new_n842), .ZN(G75));
  NOR2_X1   g657(.A1(new_n358), .A2(G952), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n823), .B1(new_n821), .B2(new_n831), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(G902), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT56), .B1(new_n847), .B2(G210), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n415), .A2(new_n423), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n422), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT55), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n845), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n848), .B2(new_n851), .ZN(G51));
  AOI21_X1  g667(.A(new_n824), .B1(new_n666), .B2(new_n667), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n819), .B1(new_n854), .B2(new_n800), .ZN(new_n855));
  INV_X1    g669(.A(new_n820), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n705), .A2(KEYINPUT42), .A3(new_n711), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n717), .A2(new_n713), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT108), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n858), .B1(new_n861), .B2(new_n715), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n810), .A2(new_n678), .ZN(new_n863));
  INV_X1    g677(.A(new_n808), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n682), .A2(new_n697), .A3(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n711), .A2(new_n699), .B1(new_n801), .B2(new_n815), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n863), .A2(new_n721), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n857), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n821), .A2(new_n831), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT54), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(KEYINPUT118), .A3(new_n832), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n846), .A2(new_n873), .A3(KEYINPUT54), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n497), .B(KEYINPUT57), .Z(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n872), .A2(KEYINPUT119), .A3(new_n874), .A4(new_n875), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n488), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n736), .B(KEYINPUT120), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n847), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n844), .B1(new_n880), .B2(new_n882), .ZN(G54));
  AND2_X1   g697(.A1(KEYINPUT58), .A2(G475), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n847), .A2(new_n577), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n846), .A2(G902), .A3(new_n884), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n576), .A3(new_n568), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n845), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT121), .ZN(G60));
  XNOR2_X1  g703(.A(new_n607), .B(KEYINPUT59), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n829), .B2(new_n832), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n603), .A2(new_n605), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n603), .B2(new_n605), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n872), .A2(new_n874), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n893), .A2(new_n894), .A3(new_n845), .A4(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n845), .B1(new_n891), .B2(new_n892), .ZN(new_n898));
  INV_X1    g712(.A(new_n896), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT122), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(G63));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT60), .Z(new_n903));
  NAND2_X1  g717(.A1(new_n846), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT123), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n846), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n365), .A3(new_n364), .A4(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n846), .A2(new_n906), .A3(new_n903), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n846), .B2(new_n903), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n626), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n911), .A3(new_n845), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n908), .A2(new_n911), .A3(KEYINPUT61), .A4(new_n845), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(G66));
  OAI21_X1  g730(.A(G953), .B1(new_n589), .B2(new_n420), .ZN(new_n917));
  INV_X1    g731(.A(new_n811), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n849), .B1(G898), .B2(new_n358), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  NOR2_X1   g735(.A1(new_n291), .A2(new_n292), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n572), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AND4_X1   g738(.A1(new_n501), .A2(new_n763), .A3(new_n648), .A4(new_n806), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n323), .A2(new_n381), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n743), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n743), .A2(KEYINPUT124), .A3(new_n926), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n929), .A2(new_n930), .B1(new_n764), .B2(new_n745), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n854), .A2(new_n659), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n854), .A2(new_n934), .A3(new_n659), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n924), .B1(new_n936), .B2(new_n358), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n923), .B1(G900), .B2(G953), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n641), .A2(new_n655), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n705), .A2(new_n648), .A3(new_n942), .A4(new_n741), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n749), .A2(new_n721), .A3(new_n743), .A4(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n854), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n862), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n941), .B1(new_n946), .B2(new_n358), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n938), .A2(new_n939), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT125), .B1(new_n937), .B2(new_n947), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n358), .B1(G227), .B2(G900), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n949), .A2(new_n951), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n959), .B2(new_n952), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n957), .A2(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(new_n946), .A2(new_n918), .ZN(new_n962));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n295), .B(KEYINPUT127), .Z(new_n966));
  AOI21_X1  g780(.A(new_n844), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n295), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n828), .A2(new_n968), .A3(new_n652), .A4(new_n964), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n936), .B2(new_n811), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n651), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n967), .A2(new_n969), .A3(new_n971), .ZN(G57));
endmodule


