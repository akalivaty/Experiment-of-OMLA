//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  INV_X1    g009(.A(G22gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G15gat), .ZN(new_n212));
  INV_X1    g011(.A(G15gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G22gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT100), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT100), .B1(new_n212), .B2(new_n214), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n210), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(new_n214), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT100), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n209), .A3(new_n215), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT101), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G8gat), .ZN(new_n225));
  INV_X1    g024(.A(G8gat), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n218), .A2(new_n222), .A3(new_n223), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G29gat), .A2(G36gat), .ZN(new_n229));
  OR2_X1    g028(.A1(KEYINPUT95), .A2(KEYINPUT14), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT95), .A2(KEYINPUT14), .ZN(new_n231));
  INV_X1    g030(.A(G29gat), .ZN(new_n232));
  INV_X1    g031(.A(G36gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n230), .A2(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n229), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G50gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G43gat), .ZN(new_n239));
  INV_X1    g038(.A(G43gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(G50gat), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT94), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT15), .ZN(new_n243));
  XNOR2_X1  g042(.A(G43gat), .B(G50gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT94), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n237), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT102), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(KEYINPUT96), .A2(G43gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(KEYINPUT96), .A2(G43gat), .ZN(new_n252));
  AOI21_X1  g051(.A(G50gat), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT97), .B1(new_n238), .B2(G43gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT97), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n240), .A3(G50gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n243), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT98), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT98), .B(new_n243), .C1(new_n253), .C2(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n242), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT99), .B1(new_n234), .B2(new_n236), .ZN(new_n264));
  AND2_X1   g063(.A1(KEYINPUT95), .A2(KEYINPUT14), .ZN(new_n265));
  NOR2_X1   g064(.A1(KEYINPUT95), .A2(KEYINPUT14), .ZN(new_n266));
  OAI22_X1  g065(.A1(new_n265), .A2(new_n266), .B1(G29gat), .B2(G36gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT99), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(new_n268), .A3(new_n235), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n263), .A2(new_n264), .A3(new_n229), .A4(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n247), .B(new_n250), .C1(new_n262), .C2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n248), .A2(new_n249), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n267), .A2(new_n268), .A3(new_n235), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n268), .B1(new_n267), .B2(new_n235), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n246), .A2(new_n242), .B1(G29gat), .B2(G36gat), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n260), .A4(new_n261), .ZN(new_n278));
  INV_X1    g077(.A(new_n272), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n278), .A2(new_n247), .A3(new_n250), .A4(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n228), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G229gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n278), .A2(new_n247), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n228), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n281), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n278), .A2(new_n225), .A3(new_n247), .A4(new_n227), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n282), .B(KEYINPUT13), .Z(new_n290));
  AOI21_X1  g089(.A(KEYINPUT103), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT103), .ZN(new_n292));
  INV_X1    g091(.A(new_n290), .ZN(new_n293));
  AOI211_X1 g092(.A(new_n292), .B(new_n293), .C1(new_n285), .C2(new_n288), .ZN(new_n294));
  OAI22_X1  g093(.A1(new_n287), .A2(KEYINPUT18), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n280), .ZN(new_n296));
  INV_X1    g095(.A(new_n228), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(new_n282), .A3(new_n285), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT18), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n208), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n300), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n287), .A2(KEYINPUT18), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n290), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n292), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n289), .A2(KEYINPUT103), .A3(new_n290), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n303), .A2(new_n304), .A3(new_n308), .A4(new_n207), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(KEYINPUT24), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT67), .ZN(new_n327));
  AOI211_X1 g126(.A(new_n312), .B(new_n318), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n329));
  INV_X1    g128(.A(new_n318), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(KEYINPUT65), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n320), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n322), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n318), .A2(new_n332), .B1(new_n333), .B2(new_n326), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n329), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n328), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(KEYINPUT66), .B(new_n329), .C1(new_n331), .C2(new_n334), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT27), .B(G183gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(G190gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT69), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n344), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n346), .ZN(new_n350));
  INV_X1    g149(.A(new_n315), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n351), .A2(new_n313), .A3(KEYINPUT26), .ZN(new_n352));
  AOI211_X1 g151(.A(new_n323), .B(new_n352), .C1(KEYINPUT26), .C2(new_n313), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n349), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(KEYINPUT75), .A3(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n357), .B(KEYINPUT74), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n354), .B1(new_n337), .B2(new_n338), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(KEYINPUT29), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n362), .B2(new_n357), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT22), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT72), .B(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G197gat), .B(G204gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n375), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n366), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n356), .A2(new_n360), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n377), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n362), .A2(KEYINPUT29), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n358), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(KEYINPUT76), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n385), .A3(new_n378), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(G8gat), .B(G36gat), .Z(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n387), .A2(KEYINPUT30), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n384), .A2(new_n386), .A3(new_n392), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(G127gat), .B(G134gat), .Z(new_n398));
  INV_X1    g197(.A(KEYINPUT70), .ZN(new_n399));
  INV_X1    g198(.A(G127gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(G134gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402));
  OAI221_X1 g201(.A(new_n398), .B1(new_n399), .B2(new_n401), .C1(KEYINPUT1), .C2(new_n402), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n402), .A2(KEYINPUT1), .B1(new_n399), .B2(new_n401), .ZN(new_n404));
  INV_X1    g203(.A(new_n398), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n409));
  XOR2_X1   g208(.A(G141gat), .B(G148gat), .Z(new_n410));
  NAND2_X1  g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT2), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G155gat), .B(G162gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(new_n414), .A3(new_n412), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n408), .B1(new_n409), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n417), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n416), .A2(KEYINPUT79), .A3(new_n417), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n420), .B1(new_n425), .B2(KEYINPUT3), .ZN(new_n426));
  AOI211_X1 g225(.A(KEYINPUT80), .B(new_n409), .C1(new_n423), .C2(new_n424), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n419), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT81), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n408), .A2(new_n418), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n407), .A2(new_n421), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n433), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n428), .A2(new_n431), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n435), .B1(new_n425), .B2(new_n407), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT5), .B1(new_n442), .B2(new_n431), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(G1gat), .B(G29gat), .Z(new_n445));
  XNOR2_X1  g244(.A(G57gat), .B(G85gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n438), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n435), .A2(KEYINPUT4), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n431), .A2(KEYINPUT5), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n424), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT79), .B1(new_n416), .B2(new_n417), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT3), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT80), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n425), .A2(new_n420), .A3(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n454), .B1(new_n460), .B2(new_n419), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n450), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT85), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n441), .B2(new_n443), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT6), .A4(new_n450), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n466), .A2(new_n450), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT6), .B1(new_n466), .B2(new_n450), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n387), .A2(new_n393), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n397), .A2(KEYINPUT86), .A3(new_n473), .A4(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n473), .A3(new_n395), .A4(new_n394), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n376), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n482), .B(new_n483), .C1(KEYINPUT87), .C2(new_n381), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n409), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n483), .B1(new_n376), .B2(new_n481), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n481), .B2(new_n378), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT88), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n421), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n483), .B1(new_n421), .B2(KEYINPUT3), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n378), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G228gat), .ZN(new_n493));
  INV_X1    g292(.A(G233gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n409), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n425), .ZN(new_n499));
  AOI211_X1 g298(.A(new_n493), .B(new_n494), .C1(new_n499), .C2(new_n492), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(G22gat), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n485), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n378), .A2(new_n481), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n504), .A2(KEYINPUT88), .A3(new_n483), .A4(new_n482), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n409), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n495), .B1(new_n506), .B2(new_n421), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n211), .B1(new_n507), .B2(new_n500), .ZN(new_n508));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT31), .B(G50gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n502), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n502), .B2(new_n508), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n477), .A2(new_n480), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n356), .A2(new_n407), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n362), .A2(new_n408), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G227gat), .A2(G233gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT71), .ZN(new_n524));
  OAI22_X1  g323(.A1(new_n521), .A2(new_n523), .B1(new_n524), .B2(KEYINPUT34), .ZN(new_n525));
  XOR2_X1   g324(.A(G15gat), .B(G43gat), .Z(new_n526));
  XNOR2_X1  g325(.A(G71gat), .B(G99gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n522), .B1(new_n519), .B2(new_n520), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(KEYINPUT33), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT34), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT71), .ZN(new_n535));
  AOI221_X4 g334(.A(new_n531), .B1(KEYINPUT33), .B2(new_n528), .C1(new_n521), .C2(new_n523), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n535), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n356), .A2(new_n407), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n362), .A2(new_n408), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n523), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT32), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT33), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n544), .A3(new_n528), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n532), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n525), .B1(new_n537), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n535), .B1(new_n533), .B2(new_n536), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(new_n546), .A3(new_n538), .ZN(new_n550));
  INV_X1    g349(.A(new_n525), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n548), .A2(KEYINPUT36), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT36), .B1(new_n548), .B2(new_n552), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n518), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT90), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n518), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT40), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n431), .B1(new_n428), .B2(new_n440), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n449), .B1(new_n562), .B2(KEYINPUT39), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n442), .A2(new_n431), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT39), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n560), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n463), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n563), .A2(new_n560), .A3(new_n566), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT30), .B1(new_n387), .B2(new_n393), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n396), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n517), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n387), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT38), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n366), .A2(new_n381), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n380), .B(new_n378), .C1(new_n382), .C2(new_n358), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(KEYINPUT37), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n576), .A2(new_n577), .A3(new_n392), .A4(new_n580), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n465), .A2(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n581), .A2(KEYINPUT91), .A3(new_n582), .A4(new_n474), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT91), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n474), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT37), .B1(new_n384), .B2(new_n386), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n577), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n586), .A2(new_n587), .A3(new_n393), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n584), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n576), .A2(new_n392), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n387), .A2(new_n575), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT38), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n574), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n557), .A2(new_n559), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT35), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n517), .B1(new_n548), .B2(new_n552), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(KEYINPUT92), .B2(new_n478), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n478), .A2(KEYINPUT92), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n477), .A2(new_n480), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(KEYINPUT35), .A3(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n311), .B1(new_n596), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT8), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  INV_X1    g408(.A(G92gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n608), .A2(KEYINPUT106), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT106), .B1(new_n608), .B2(new_n611), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT107), .ZN(new_n615));
  XOR2_X1   g414(.A(G99gat), .B(G106gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT7), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n614), .A2(new_n615), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n612), .B2(new_n613), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n616), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n617), .B(new_n619), .C1(new_n612), .C2(new_n613), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(KEYINPUT107), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n296), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT108), .Z(new_n627));
  NAND2_X1  g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT41), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n620), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n284), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n625), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT109), .ZN(new_n634));
  XOR2_X1   g433(.A(G134gat), .B(G162gat), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n628), .A2(new_n629), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n625), .A2(new_n632), .ZN(new_n639));
  INV_X1    g438(.A(new_n627), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n633), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n638), .A2(new_n642), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G57gat), .B(G64gat), .Z(new_n646));
  INV_X1    g445(.A(KEYINPUT9), .ZN(new_n647));
  INV_X1    g446(.A(G71gat), .ZN(new_n648));
  INV_X1    g447(.A(G78gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G71gat), .B(G78gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(KEYINPUT21), .ZN(new_n654));
  XNOR2_X1  g453(.A(G127gat), .B(G155gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n228), .B1(KEYINPUT21), .B2(new_n653), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT105), .ZN(new_n660));
  NAND2_X1  g459(.A1(G231gat), .A2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT104), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G183gat), .B(G211gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n658), .B(new_n665), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n645), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n651), .B(new_n652), .Z(new_n670));
  NAND3_X1  g469(.A1(new_n624), .A2(new_n620), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n624), .A2(new_n670), .A3(KEYINPUT110), .A4(new_n620), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n653), .A2(new_n623), .A3(new_n622), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n631), .A2(KEYINPUT10), .A3(new_n653), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n669), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n668), .B1(new_n675), .B2(new_n677), .ZN(new_n681));
  XNOR2_X1  g480(.A(G120gat), .B(G148gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(G176gat), .B(G204gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n680), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n677), .ZN(new_n687));
  AOI211_X1 g486(.A(KEYINPUT10), .B(new_n687), .C1(new_n673), .C2(new_n674), .ZN(new_n688));
  INV_X1    g487(.A(new_n679), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n668), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n681), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n684), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n667), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n606), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n473), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(new_n209), .ZN(G1324gat));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n396), .A2(new_n571), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT16), .B(G8gat), .ZN(new_n701));
  OR4_X1    g500(.A1(new_n699), .A2(new_n696), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n606), .A2(new_n695), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n704));
  INV_X1    g503(.A(new_n700), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT112), .B1(new_n696), .B2(new_n700), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(G8gat), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n701), .B1(new_n706), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n702), .B(new_n708), .C1(new_n709), .C2(new_n710), .ZN(G1325gat));
  NAND2_X1  g510(.A1(new_n548), .A2(new_n552), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n703), .A2(new_n213), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G15gat), .B1(new_n696), .B2(new_n555), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1326gat));
  NOR2_X1   g514(.A1(new_n696), .A2(new_n573), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT43), .B(G22gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  INV_X1    g517(.A(new_n645), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n694), .A2(new_n666), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n606), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n723), .A2(G29gat), .A3(new_n473), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n724), .A2(KEYINPUT45), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(KEYINPUT45), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n596), .A2(new_n605), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n645), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n601), .B(new_n603), .C1(new_n556), .C2(new_n594), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT44), .B1(new_n731), .B2(new_n719), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n720), .A2(new_n310), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n734), .A2(new_n473), .A3(new_n735), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n725), .B(new_n726), .C1(new_n736), .C2(new_n232), .ZN(G1328gat));
  NAND2_X1  g536(.A1(new_n705), .A2(new_n233), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT46), .B1(new_n723), .B2(new_n738), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n738), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n734), .A2(new_n700), .A3(new_n735), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n233), .ZN(G1329gat));
  NAND2_X1  g541(.A1(new_n251), .A2(new_n252), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n712), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n723), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n735), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n555), .A2(new_n744), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n730), .A2(new_n733), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g550(.A(new_n729), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n596), .B2(new_n605), .ZN(new_n753));
  NOR4_X1   g552(.A1(new_n753), .A2(new_n732), .A3(new_n573), .A4(new_n735), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT113), .B1(new_n754), .B2(new_n238), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n606), .A2(new_n238), .A3(new_n517), .A4(new_n722), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n754), .B2(new_n238), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OAI221_X1 g558(.A(new_n756), .B1(KEYINPUT113), .B2(KEYINPUT48), .C1(new_n754), .C2(new_n238), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1331gat));
  NOR3_X1   g560(.A1(new_n667), .A2(new_n310), .A3(new_n693), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n731), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n582), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT114), .B(G57gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1332gat));
  AOI21_X1  g565(.A(new_n700), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT115), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT116), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT117), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n769), .B(new_n772), .ZN(G1333gat));
  INV_X1    g572(.A(new_n555), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n648), .B1(new_n763), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n745), .A2(G71gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n763), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n517), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n310), .A2(new_n666), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n693), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n730), .A2(new_n733), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n473), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n731), .A2(new_n719), .A3(new_n781), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n731), .A2(KEYINPUT51), .A3(new_n719), .A4(new_n781), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n694), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n582), .A2(new_n609), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n785), .B1(new_n792), .B2(new_n793), .ZN(G1336gat));
  OAI21_X1  g593(.A(G92gat), .B1(new_n784), .B2(new_n700), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n700), .A2(G92gat), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n795), .B(new_n796), .C1(new_n792), .C2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n783), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n753), .A2(new_n732), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n610), .B1(new_n801), .B2(new_n705), .ZN(new_n802));
  AOI211_X1 g601(.A(new_n693), .B(new_n798), .C1(new_n788), .C2(new_n790), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT52), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(new_n804), .ZN(G1337gat));
  OAI21_X1  g604(.A(G99gat), .B1(new_n784), .B2(new_n555), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n745), .A2(G99gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n792), .B2(new_n807), .ZN(G1338gat));
  NAND4_X1  g607(.A1(new_n730), .A2(new_n733), .A3(new_n517), .A4(new_n783), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n573), .A2(G106gat), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n694), .B(new_n811), .C1(new_n789), .C2(new_n791), .ZN(new_n812));
  XNOR2_X1  g611(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n810), .B2(new_n812), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(G1339gat));
  NAND2_X1  g615(.A1(new_n695), .A2(new_n311), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n684), .B1(new_n680), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n678), .A2(new_n669), .A3(new_n679), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n690), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n822), .A3(KEYINPUT55), .ZN(new_n823));
  INV_X1    g622(.A(new_n686), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT55), .B1(new_n820), .B2(new_n822), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n282), .B1(new_n298), .B2(new_n285), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n289), .A2(new_n290), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n206), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n309), .A2(new_n829), .ZN(new_n830));
  NOR4_X1   g629(.A1(new_n645), .A2(new_n825), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n309), .B(new_n829), .C1(new_n686), .C2(new_n692), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n690), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n685), .B1(new_n690), .B2(KEYINPUT54), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n310), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n833), .B(new_n834), .C1(new_n839), .C2(new_n825), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n645), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n820), .A2(new_n822), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n835), .A2(new_n842), .B1(new_n302), .B2(new_n309), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n823), .A2(new_n824), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n833), .B1(new_n845), .B2(new_n834), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n832), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n666), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n818), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n517), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n705), .A2(new_n473), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n712), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n310), .ZN(new_n856));
  INV_X1    g655(.A(new_n834), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n844), .B2(new_n843), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n719), .B1(new_n858), .B2(new_n833), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n845), .A2(new_n834), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT119), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n831), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n817), .B1(new_n862), .B2(new_n666), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT120), .B1(new_n863), .B2(new_n573), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n849), .A2(new_n865), .A3(new_n517), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n853), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT121), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n853), .B(new_n870), .C1(new_n864), .C2(new_n866), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n310), .A2(G113gat), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n856), .B1(new_n873), .B2(new_n874), .ZN(G1340gat));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n868), .A2(new_n694), .A3(new_n871), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(G120gat), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n693), .A2(G120gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n854), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  AOI211_X1 g681(.A(KEYINPUT122), .B(new_n880), .C1(new_n877), .C2(G120gat), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(G1341gat));
  NAND3_X1  g683(.A1(new_n855), .A2(new_n400), .A3(new_n666), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n869), .A2(new_n872), .A3(new_n848), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n400), .ZN(G1342gat));
  NOR3_X1   g686(.A1(new_n849), .A2(new_n517), .A3(new_n745), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n700), .A2(new_n719), .ZN(new_n890));
  NOR4_X1   g689(.A1(new_n889), .A2(G134gat), .A3(new_n473), .A4(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT56), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n869), .A2(new_n872), .A3(new_n645), .ZN(new_n893));
  INV_X1    g692(.A(G134gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(G1343gat));
  NOR4_X1   g694(.A1(new_n849), .A2(new_n774), .A3(new_n473), .A4(new_n573), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n311), .A2(G141gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n700), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n849), .A2(new_n573), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n555), .A2(new_n851), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n831), .B1(new_n645), .B2(new_n860), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n817), .B1(new_n905), .B2(new_n666), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n517), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n904), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n903), .A2(new_n908), .A3(new_n310), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT58), .B1(new_n909), .B2(G141gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n900), .A2(new_n910), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n909), .A2(KEYINPUT123), .A3(G141gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT123), .B1(new_n909), .B2(G141gat), .ZN(new_n913));
  INV_X1    g712(.A(new_n904), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n901), .A2(new_n914), .A3(new_n899), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(G1344gat));
  INV_X1    g717(.A(G148gat), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n898), .A2(new_n919), .A3(new_n700), .A4(new_n694), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n903), .A2(new_n908), .ZN(new_n921));
  AOI211_X1 g720(.A(KEYINPUT59), .B(new_n919), .C1(new_n921), .C2(new_n694), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT57), .B1(new_n849), .B2(new_n573), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n902), .A3(new_n517), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n694), .A3(new_n914), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n923), .B1(new_n927), .B2(G148gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n920), .B1(new_n922), .B2(new_n928), .ZN(G1345gat));
  NOR2_X1   g728(.A1(new_n848), .A2(G155gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n898), .A2(new_n700), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n921), .A2(new_n666), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G155gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1346gat));
  NAND2_X1  g733(.A1(new_n921), .A2(new_n719), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G162gat), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n890), .A2(G162gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n898), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1347gat));
  NOR2_X1   g738(.A1(new_n700), .A2(new_n582), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n888), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G169gat), .B1(new_n942), .B2(new_n310), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n712), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n850), .A2(KEYINPUT120), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n865), .B1(new_n849), .B2(new_n517), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n310), .A2(G169gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(G1348gat));
  INV_X1    g748(.A(G176gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n942), .A2(new_n950), .A3(new_n694), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n947), .A2(new_n694), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n950), .ZN(G1349gat));
  NAND2_X1  g752(.A1(new_n666), .A2(new_n340), .ZN(new_n954));
  OR3_X1    g753(.A1(new_n941), .A2(KEYINPUT125), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT125), .B1(new_n941), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n947), .A2(new_n666), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G183gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g760(.A(G190gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n942), .A2(new_n962), .A3(new_n719), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n947), .B2(new_n719), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1351gat));
  AND2_X1   g767(.A1(new_n555), .A2(new_n940), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n901), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  OR3_X1    g770(.A1(new_n971), .A2(G197gat), .A3(new_n311), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n926), .A2(new_n969), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n310), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G197gat), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n975), .A2(new_n976), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n972), .B1(new_n978), .B2(new_n979), .ZN(G1352gat));
  NOR3_X1   g779(.A1(new_n971), .A2(G204gat), .A3(new_n693), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT62), .ZN(new_n982));
  OAI21_X1  g781(.A(G204gat), .B1(new_n973), .B2(new_n693), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1353gat));
  NAND3_X1  g783(.A1(new_n970), .A2(new_n371), .A3(new_n666), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n974), .A2(new_n666), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  AOI21_X1  g788(.A(G218gat), .B1(new_n970), .B2(new_n719), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT127), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n973), .A2(new_n372), .A3(new_n645), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(G1355gat));
endmodule


