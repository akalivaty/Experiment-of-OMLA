//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n193), .A2(new_n194), .A3(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT2), .B(G113), .Z(new_n197));
  XNOR2_X1  g011(.A(G116), .B(G119), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n196), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  OAI22_X1  g013(.A1(new_n195), .A2(new_n199), .B1(new_n198), .B2(new_n197), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(G107), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT4), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(G101), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(G101), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n212), .B(new_n203), .C1(new_n205), .C2(new_n206), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n211), .A2(new_n208), .A3(KEYINPUT4), .A4(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n200), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n197), .A2(new_n198), .A3(new_n196), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT67), .B1(new_n193), .B2(new_n194), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n202), .A2(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n206), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(G113), .C1(KEYINPUT5), .C2(new_n190), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n215), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT6), .ZN(new_n226));
  XNOR2_X1  g040(.A(G110), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n215), .A2(new_n224), .A3(new_n227), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT6), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n227), .B1(new_n215), .B2(new_n224), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT85), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G143), .ZN(new_n236));
  INV_X1    g050(.A(G143), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT0), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n239), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G143), .B(G146), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n241), .B2(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G125), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n237), .C2(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G128), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT66), .B1(new_n236), .B2(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n239), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n245), .A2(new_n253), .A3(G128), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n248), .B1(new_n255), .B2(G125), .ZN(new_n256));
  INV_X1    g070(.A(G224), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G953), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n256), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n231), .B2(new_n232), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n234), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n221), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n218), .A2(new_n223), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n227), .B(KEYINPUT8), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT7), .ZN(new_n271));
  OAI221_X1 g085(.A(new_n248), .B1(new_n271), .B2(new_n258), .C1(new_n255), .C2(G125), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n270), .A2(new_n230), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n259), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT87), .ZN(new_n275));
  AOI21_X1  g089(.A(G902), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n263), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G210), .B1(G237), .B2(G902), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n263), .A2(new_n278), .A3(new_n276), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n188), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G475), .ZN(new_n284));
  NOR2_X1   g098(.A1(G237), .A2(G953), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G214), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n237), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(G143), .A3(G214), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT88), .B1(new_n289), .B2(G131), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT17), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(G131), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n293));
  INV_X1    g107(.A(G131), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n287), .A2(new_n293), .A3(new_n294), .A4(new_n288), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G125), .B(G140), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT16), .ZN(new_n298));
  INV_X1    g112(.A(G125), .ZN(new_n299));
  OR3_X1    g113(.A1(new_n299), .A2(KEYINPUT16), .A3(G140), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n235), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n298), .A2(G146), .A3(new_n300), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n289), .A2(KEYINPUT17), .A3(G131), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n296), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n289), .A2(KEYINPUT18), .A3(G131), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT18), .A2(G131), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n287), .A2(new_n288), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n297), .B(new_n235), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G113), .B(G122), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(new_n204), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n305), .A2(new_n313), .A3(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G902), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n284), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT19), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n297), .B(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n303), .B1(new_n321), .B2(G146), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n292), .A2(new_n295), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(new_n290), .ZN(new_n324));
  INV_X1    g138(.A(new_n310), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n314), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n328));
  NOR2_X1   g142(.A1(G475), .A2(G902), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n328), .B1(new_n327), .B2(new_n329), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n327), .A2(KEYINPUT89), .A3(new_n328), .A4(new_n329), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n319), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n237), .A2(G128), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n242), .A2(G143), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(G134), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n340), .A3(G134), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G122), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G116), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n191), .A2(G122), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n202), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(G107), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n336), .A2(new_n337), .A3(new_n340), .A4(G134), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n342), .A2(new_n347), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT14), .A4(G107), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n344), .A2(KEYINPUT14), .A3(G107), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n347), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n339), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n339), .A2(new_n353), .A3(KEYINPUT90), .A4(new_n351), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n350), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT9), .B(G234), .Z(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT77), .ZN(new_n360));
  INV_X1    g174(.A(G953), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(G217), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n350), .A2(new_n364), .A3(new_n356), .A4(new_n357), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(KEYINPUT91), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n358), .A2(new_n367), .A3(new_n362), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n318), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G478), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n370), .A2(KEYINPUT15), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n369), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n361), .A2(G952), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(G234), .B2(G237), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(G234), .A2(G237), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(G902), .A3(G953), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT92), .ZN(new_n378));
  XOR2_X1   g192(.A(KEYINPUT21), .B(G898), .Z(new_n379));
  OAI21_X1  g193(.A(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT93), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n335), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n283), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT11), .ZN(new_n384));
  INV_X1    g198(.A(G134), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(G137), .ZN(new_n386));
  INV_X1    g200(.A(G137), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT11), .A3(G134), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(G137), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(KEYINPUT65), .A2(G131), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n391), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT1), .B1(new_n237), .B2(G146), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n397), .A2(G128), .B1(new_n236), .B2(new_n238), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n254), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n242), .B1(new_n236), .B2(KEYINPUT1), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n401), .A2(new_n245), .A3(KEYINPUT79), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n221), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT80), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT79), .B1(new_n401), .B2(new_n245), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n397), .A2(G128), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n399), .A3(new_n239), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n407), .A3(new_n254), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n221), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n396), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n213), .A2(KEYINPUT10), .A3(new_n220), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n252), .A2(new_n413), .A3(new_n254), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n252), .B2(new_n254), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n214), .A2(new_n247), .A3(new_n210), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n394), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n408), .A2(new_n409), .A3(new_n221), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n409), .B1(new_n408), .B2(new_n221), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n395), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n394), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n417), .A4(new_n416), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G140), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n361), .A2(G227), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n427), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n252), .A2(new_n254), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(new_n221), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n420), .B2(new_n421), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT12), .A3(new_n394), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT12), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n404), .B2(new_n410), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n435), .B1(new_n436), .B2(new_n423), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n411), .A2(new_n418), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n434), .A2(new_n437), .B1(new_n438), .B2(new_n423), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n429), .B1(new_n439), .B2(KEYINPUT82), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n436), .A2(new_n435), .A3(new_n423), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT12), .B1(new_n433), .B2(new_n394), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT82), .B(new_n424), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(G469), .B(new_n428), .C1(new_n440), .C2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n424), .B(new_n427), .C1(new_n441), .C2(new_n442), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n427), .B1(new_n419), .B2(new_n424), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n448), .B2(KEYINPUT83), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n450));
  AOI211_X1 g264(.A(new_n450), .B(new_n427), .C1(new_n419), .C2(new_n424), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n446), .B(new_n318), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(G469), .A2(G902), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n445), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G221), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n360), .B2(new_n318), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n454), .A2(KEYINPUT84), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT84), .B1(new_n454), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n383), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT94), .ZN(new_n461));
  XOR2_X1   g275(.A(G125), .B(G140), .Z(new_n462));
  NAND2_X1  g276(.A1(new_n242), .A2(G119), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n189), .A2(G128), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT24), .B(G110), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT75), .Z(new_n468));
  AOI21_X1  g282(.A(KEYINPUT73), .B1(new_n242), .B2(G119), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT23), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n470), .B2(new_n469), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT74), .B(G110), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI221_X1 g288(.A(new_n303), .B1(G146), .B2(new_n462), .C1(new_n468), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n302), .A2(new_n303), .ZN(new_n476));
  INV_X1    g290(.A(G110), .ZN(new_n477));
  OAI221_X1 g291(.A(new_n476), .B1(new_n477), .B2(new_n472), .C1(new_n465), .C2(new_n466), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT22), .B(G137), .ZN(new_n480));
  INV_X1    g294(.A(G234), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n455), .A2(new_n481), .A3(G953), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n480), .B(new_n482), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n475), .A2(new_n478), .A3(new_n483), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n318), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT25), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G217), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(G234), .B2(new_n318), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(G902), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT76), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n485), .A2(new_n486), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(G472), .A2(G902), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT26), .B(G101), .Z(new_n499));
  NAND2_X1  g313(.A1(new_n285), .A2(G210), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n390), .A2(new_n294), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n294), .B1(G134), .B2(new_n387), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n389), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n414), .B2(new_n415), .ZN(new_n509));
  INV_X1    g323(.A(new_n200), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n392), .A2(new_n393), .B1(new_n244), .B2(new_n246), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n255), .A2(new_n507), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n200), .B1(new_n519), .B2(new_n511), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT28), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n503), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n509), .A2(KEYINPUT30), .A3(new_n512), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n519), .B2(new_n511), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n200), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n513), .A3(new_n503), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT31), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT31), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n527), .A2(new_n530), .A3(new_n513), .A4(new_n503), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n498), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n527), .A2(new_n513), .ZN(new_n536));
  INV_X1    g350(.A(new_n503), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT29), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n513), .A2(new_n515), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT70), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n540), .A2(new_n522), .A3(new_n541), .A4(new_n503), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n430), .A2(KEYINPUT68), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n252), .A2(new_n413), .A3(new_n254), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n507), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n200), .B1(new_n546), .B2(new_n511), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT71), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n513), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n509), .A2(KEYINPUT71), .A3(new_n510), .A4(new_n512), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT28), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n518), .A2(new_n551), .A3(KEYINPUT29), .A4(new_n503), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n543), .A2(new_n552), .A3(new_n318), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n540), .A2(new_n522), .A3(new_n541), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n529), .B(new_n531), .C1(new_n555), .C2(new_n503), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT32), .A3(new_n498), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n535), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT72), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n535), .A2(new_n554), .A3(new_n557), .A4(KEYINPUT72), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n497), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n383), .B(new_n563), .C1(new_n458), .C2(new_n459), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n461), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(G101), .ZN(G3));
  NAND2_X1  g380(.A1(new_n454), .A2(new_n457), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT84), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n454), .A2(KEYINPUT84), .A3(new_n457), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n369), .A2(new_n370), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n369), .A2(KEYINPUT95), .A3(new_n370), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n366), .A2(new_n577), .A3(new_n368), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n363), .A2(KEYINPUT33), .A3(new_n365), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(G478), .A3(new_n318), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n335), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n281), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n278), .B1(new_n263), .B2(new_n276), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n187), .B(new_n381), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT96), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n335), .B1(new_n576), .B2(new_n581), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n589), .A2(new_n282), .A3(new_n590), .A4(new_n381), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G472), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n556), .B2(new_n318), .ZN(new_n594));
  INV_X1    g408(.A(new_n533), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n497), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n571), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT34), .B(G104), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G6));
  NAND2_X1  g415(.A1(new_n327), .A2(new_n329), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n330), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT97), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n606), .A3(new_n330), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n319), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n372), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n587), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n571), .A2(new_n598), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT35), .B(G107), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G9));
  NOR2_X1   g428(.A1(new_n484), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n479), .B(new_n615), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n489), .A2(new_n491), .B1(new_n494), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n597), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n461), .A2(new_n564), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT37), .B(G110), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G12));
  AOI21_X1  g435(.A(new_n617), .B1(new_n560), .B2(new_n561), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n378), .A2(G900), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n374), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(KEYINPUT98), .Z(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n608), .A2(new_n609), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n622), .A2(new_n571), .A3(new_n282), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G128), .ZN(G30));
  XNOR2_X1  g444(.A(new_n625), .B(KEYINPUT39), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n569), .B2(new_n570), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n535), .A2(new_n557), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n549), .A2(new_n537), .A3(new_n550), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n636), .A2(new_n528), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n637), .B2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n280), .A2(new_n281), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n335), .A2(new_n372), .ZN(new_n643));
  INV_X1    g457(.A(new_n617), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n188), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n634), .A2(new_n639), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n632), .A2(new_n633), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n237), .ZN(G45));
  NOR2_X1   g464(.A1(new_n584), .A2(new_n625), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n622), .A2(new_n571), .A3(new_n282), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  OAI21_X1  g467(.A(new_n318), .B1(new_n449), .B2(new_n451), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G469), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n457), .A3(new_n452), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n655), .A2(KEYINPUT100), .A3(new_n457), .A4(new_n452), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n562), .A2(new_n592), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT41), .B(G113), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G15));
  NAND3_X1  g477(.A1(new_n562), .A2(new_n611), .A3(new_n660), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G116), .ZN(G18));
  NAND4_X1  g479(.A1(new_n282), .A2(new_n457), .A3(new_n452), .A4(new_n655), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n382), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n622), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G119), .ZN(G21));
  NAND3_X1  g483(.A1(new_n282), .A2(new_n381), .A3(new_n643), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n658), .B2(new_n659), .ZN(new_n671));
  INV_X1    g485(.A(new_n498), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n518), .A2(new_n551), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n518), .A2(new_n551), .A3(KEYINPUT101), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n537), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n532), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n672), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n497), .A2(new_n679), .A3(new_n594), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n671), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G122), .ZN(G24));
  INV_X1    g496(.A(new_n666), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n679), .A2(new_n594), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n684), .B1(new_n685), .B2(new_n644), .ZN(new_n686));
  NOR4_X1   g500(.A1(new_n679), .A2(new_n617), .A3(new_n594), .A4(KEYINPUT102), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n651), .B(new_n683), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT103), .B(G125), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G27));
  AOI21_X1  g504(.A(KEYINPUT32), .B1(new_n556), .B2(new_n498), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n557), .B1(new_n691), .B2(KEYINPUT104), .ZN(new_n692));
  OR3_X1    g506(.A1(new_n533), .A2(KEYINPUT104), .A3(new_n534), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n554), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n497), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n567), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n280), .A2(new_n187), .A3(new_n281), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n651), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT42), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n567), .A2(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n589), .A2(new_n626), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n562), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n294), .ZN(G33));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n627), .B(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n562), .A3(new_n702), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT106), .B(G134), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G36));
  INV_X1    g526(.A(new_n631), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n428), .B1(new_n440), .B2(new_n444), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n446), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(new_n715), .B2(new_n714), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(KEYINPUT46), .A3(new_n453), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n452), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT46), .B1(new_n717), .B2(new_n453), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n457), .B(new_n713), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n582), .A2(new_n335), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(KEYINPUT43), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n582), .A2(new_n335), .B1(new_n724), .B2(KEYINPUT43), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n726), .B1(new_n727), .B2(new_n725), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n597), .A3(new_n644), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n698), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n722), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G137), .ZN(G39));
  OAI21_X1  g548(.A(new_n457), .B1(new_n719), .B2(new_n720), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT47), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n737), .B(new_n457), .C1(new_n719), .C2(new_n720), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n560), .A2(new_n561), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n739), .A2(new_n695), .A3(new_n703), .A4(new_n698), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n736), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G140), .ZN(G42));
  NAND3_X1  g556(.A1(new_n695), .A2(new_n457), .A3(new_n187), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n743), .A2(new_n642), .A3(new_n723), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n655), .A2(new_n452), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT49), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n635), .A3(new_n746), .A4(new_n638), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n562), .B(new_n660), .C1(new_n592), .C2(new_n611), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n609), .A2(new_n335), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n750), .B1(new_n587), .B2(new_n751), .ZN(new_n752));
  OR3_X1    g566(.A1(new_n587), .A2(new_n750), .A3(new_n751), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n571), .A2(new_n598), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n749), .A2(new_n668), .A3(new_n681), .A4(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n461), .A2(new_n564), .A3(new_n618), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n699), .A2(new_n626), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n622), .A2(new_n571), .A3(new_n372), .A4(new_n608), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n697), .B(new_n589), .C1(new_n686), .C2(new_n687), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n701), .A2(new_n710), .A3(new_n705), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n584), .A2(new_n587), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n571), .A2(new_n598), .A3(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n565), .A2(KEYINPUT108), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT108), .B1(new_n565), .B2(new_n765), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n757), .B(new_n763), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n644), .A2(new_n625), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n282), .A2(new_n643), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n639), .A2(new_n697), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n629), .A2(new_n652), .A3(new_n688), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT52), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n748), .B1(new_n768), .B2(new_n773), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n622), .A2(new_n667), .B1(new_n671), .B2(new_n680), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n619), .A2(new_n754), .A3(new_n775), .A4(new_n749), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n565), .A2(new_n765), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n565), .A2(KEYINPUT108), .A3(new_n765), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n772), .B(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n783), .A3(KEYINPUT53), .A4(new_n763), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n774), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(KEYINPUT110), .B(new_n748), .C1(new_n768), .C2(new_n773), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n774), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(KEYINPUT111), .B(new_n748), .C1(new_n768), .C2(new_n773), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n788), .B1(new_n792), .B2(KEYINPUT54), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  INV_X1    g608(.A(new_n728), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n795), .B2(new_n375), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n728), .A2(KEYINPUT112), .A3(new_n374), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n680), .A3(new_n699), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n736), .A2(new_n738), .ZN(new_n802));
  INV_X1    g616(.A(new_n745), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n456), .B1(new_n803), .B2(KEYINPUT114), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(KEYINPUT114), .B2(new_n803), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n800), .B(new_n801), .C1(new_n802), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT51), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n656), .A2(new_n698), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT115), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n810), .A2(new_n497), .A3(new_n375), .A4(new_n639), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n335), .A3(new_n576), .A4(new_n581), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n810), .B1(new_n796), .B2(new_n797), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n687), .B2(new_n686), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n642), .A2(new_n187), .A3(new_n656), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n798), .A2(new_n680), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n815), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n806), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n808), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n821), .B(new_n806), .C1(new_n807), .C2(KEYINPUT51), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n373), .B1(new_n811), .B2(new_n589), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n798), .A2(new_n683), .A3(new_n680), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(KEYINPUT117), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n696), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n813), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT48), .Z(new_n830));
  AOI21_X1  g644(.A(KEYINPUT117), .B1(new_n825), .B2(new_n826), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n823), .A2(new_n824), .A3(new_n827), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n793), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(G952), .A2(G953), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n747), .B1(new_n834), .B2(new_n835), .ZN(G75));
  NAND4_X1  g650(.A1(new_n790), .A2(G210), .A3(G902), .A4(new_n791), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n234), .A2(new_n262), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(new_n260), .ZN(new_n840));
  XOR2_X1   g654(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n837), .A2(new_n838), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n837), .B2(new_n838), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n361), .A2(G952), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G51));
  XOR2_X1   g660(.A(new_n453), .B(KEYINPUT57), .Z(new_n847));
  AND3_X1   g661(.A1(new_n790), .A2(KEYINPUT54), .A3(new_n791), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT54), .B1(new_n790), .B2(new_n791), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n449), .A2(new_n451), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n790), .A2(new_n791), .ZN(new_n853));
  OR3_X1    g667(.A1(new_n853), .A2(new_n318), .A3(new_n717), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n845), .B1(new_n852), .B2(new_n854), .ZN(G54));
  INV_X1    g669(.A(new_n845), .ZN(new_n856));
  NAND2_X1  g670(.A1(KEYINPUT58), .A2(G475), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT119), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n790), .A2(G902), .A3(new_n791), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n327), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT120), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n859), .A2(new_n864), .A3(new_n860), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n861), .B1(new_n863), .B2(new_n865), .ZN(G60));
  NAND2_X1  g680(.A1(G478), .A2(G902), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT59), .Z(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n580), .B1(new_n793), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n580), .A2(new_n869), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n848), .B2(new_n849), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n856), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n870), .A2(new_n873), .ZN(G63));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n875));
  NAND2_X1  g689(.A1(G217), .A2(G902), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT121), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT60), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n790), .A2(new_n791), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n496), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n616), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n856), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n875), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n792), .A2(new_n616), .A3(new_n878), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(KEYINPUT61), .A3(new_n856), .A4(new_n880), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(G66));
  AOI21_X1  g701(.A(new_n361), .B1(new_n379), .B2(G224), .ZN(new_n888));
  INV_X1    g702(.A(new_n781), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n361), .ZN(new_n890));
  INV_X1    g704(.A(G898), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n839), .B1(new_n891), .B2(G953), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n890), .B(new_n892), .ZN(G69));
  NAND2_X1  g707(.A1(new_n524), .A2(new_n526), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(new_n321), .Z(new_n895));
  AOI21_X1  g709(.A(new_n698), .B1(new_n584), .B2(new_n751), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n632), .A2(new_n562), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n733), .A2(new_n741), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n629), .A2(new_n688), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(new_n652), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n647), .A2(new_n648), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(KEYINPUT62), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n652), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n903), .B1(new_n904), .B2(new_n649), .ZN(new_n905));
  AOI211_X1 g719(.A(KEYINPUT122), .B(new_n898), .C1(new_n902), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n902), .A2(new_n905), .ZN(new_n908));
  INV_X1    g722(.A(new_n898), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n895), .B1(new_n911), .B2(G953), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n828), .A2(new_n770), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n721), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(KEYINPUT124), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n721), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n762), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n733), .A2(new_n741), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n361), .A4(new_n900), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n895), .B1(G900), .B2(G953), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n361), .B1(G227), .B2(G900), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT125), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n928));
  INV_X1    g742(.A(new_n925), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND4_X1   g744(.A1(new_n912), .A2(new_n922), .A3(new_n926), .A4(new_n930), .ZN(new_n931));
  AOI22_X1  g745(.A1(new_n912), .A2(new_n922), .B1(new_n930), .B2(new_n926), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(G72));
  NAND2_X1  g747(.A1(G472), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT63), .Z(new_n935));
  NAND3_X1  g749(.A1(new_n918), .A2(new_n919), .A3(new_n900), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n889), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n536), .B(KEYINPUT126), .Z(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n503), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n845), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n935), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n911), .B2(new_n781), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n938), .A2(new_n503), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n536), .A2(new_n537), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n945), .B2(new_n528), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n786), .A2(new_n787), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT127), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n947), .A2(KEYINPUT127), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(G57));
endmodule


