//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR2_X1   g0000(.A1(G50), .A2(G58), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n202), .A2(new_n205), .ZN(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT64), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT65), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n217), .B1(new_n203), .B2(new_n218), .C1(new_n204), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  NAND2_X1  g0028(.A1(new_n224), .A2(new_n203), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n216), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(new_n215), .B2(new_n214), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  NOR2_X1   g0046(.A1(new_n203), .A2(new_n204), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n205), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT67), .ZN(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G87), .B(G97), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT68), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n252), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(KEYINPUT10), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n232), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n224), .A2(KEYINPUT8), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G58), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n233), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n265), .A2(new_n267), .B1(G150), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n233), .B1(new_n201), .B2(new_n203), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n261), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(G50), .B1(new_n233), .B2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(G50), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n274), .A2(new_n261), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n279), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n222), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT71), .B1(new_n272), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n233), .A2(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n285), .A2(new_n266), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n260), .B1(new_n289), .B2(new_n270), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT71), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(new_n282), .A4(new_n280), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n284), .A2(new_n292), .A3(KEYINPUT9), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT72), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n284), .A2(new_n292), .A3(KEYINPUT72), .A4(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  AOI21_X1  g0099(.A(G1), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G1), .A3(G13), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n302), .A3(G274), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n223), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT3), .B(G33), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(new_n310), .A3(G222), .ZN(new_n311));
  OR2_X1    g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(G77), .A3(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  OAI211_X1 g0116(.A(G223), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n311), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n306), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G190), .ZN(new_n321));
  INV_X1    g0121(.A(G200), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n320), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT9), .B1(new_n284), .B2(new_n292), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n258), .B1(new_n297), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT73), .B1(new_n320), .B2(new_n322), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT73), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n317), .A2(new_n314), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n302), .B1(new_n330), .B2(new_n311), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n329), .B(G200), .C1(new_n331), .C2(new_n306), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n321), .A2(new_n258), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n333), .A2(new_n324), .A3(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n335), .A2(KEYINPUT74), .A3(new_n297), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT74), .B1(new_n335), .B2(new_n297), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n327), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n320), .A2(G169), .B1(new_n272), .B2(new_n283), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n331), .A2(G179), .A3(new_n306), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n303), .B1(new_n305), .B2(new_n219), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n315), .A2(new_n316), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G107), .ZN(new_n345));
  OAI21_X1  g0145(.A(G238), .B1(new_n315), .B2(new_n316), .ZN(new_n346));
  INV_X1    g0146(.A(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT69), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n347), .ZN(new_n349));
  NAND2_X1  g0149(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n350), .C1(new_n315), .C2(new_n316), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n345), .B1(new_n346), .B2(new_n347), .C1(new_n351), .C2(new_n225), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n343), .B1(new_n352), .B2(new_n319), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G190), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n265), .A2(new_n268), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n261), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n281), .A2(new_n260), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(G77), .A3(new_n276), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(G77), .B2(new_n279), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n354), .B(new_n363), .C1(new_n322), .C2(new_n353), .ZN(new_n364));
  INV_X1    g0164(.A(new_n363), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(G169), .B2(new_n353), .ZN(new_n366));
  INV_X1    g0166(.A(G179), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n353), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n338), .A2(new_n342), .A3(new_n364), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G232), .A2(G1698), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n312), .B2(new_n313), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G97), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT75), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(G33), .A3(G97), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n309), .A2(new_n310), .A3(G226), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n302), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n303), .B1(new_n305), .B2(new_n218), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT13), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n309), .A2(new_n310), .A3(G226), .ZN(new_n384));
  INV_X1    g0184(.A(new_n372), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n315), .B2(new_n316), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n375), .A3(new_n377), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n319), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT13), .ZN(new_n389));
  INV_X1    g0189(.A(new_n382), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n383), .A2(new_n391), .A3(G179), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n383), .A2(new_n391), .A3(KEYINPUT76), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n388), .A2(new_n394), .A3(new_n390), .A4(new_n389), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(G169), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(KEYINPUT77), .A2(KEYINPUT14), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n397), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n393), .A2(new_n395), .A3(G169), .A4(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n392), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n203), .A2(G20), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n402), .B1(new_n266), .B2(new_n204), .C1(new_n222), .C2(new_n288), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT11), .A3(new_n260), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n279), .A2(G68), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT12), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n360), .A2(G68), .A3(new_n276), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT11), .B1(new_n403), .B2(new_n260), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n383), .A2(new_n391), .A3(G190), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n413), .A2(new_n411), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n393), .A2(G200), .A3(new_n395), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G58), .A2(G68), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n233), .B1(new_n229), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G159), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n288), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT78), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(G58), .A2(G68), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G58), .A2(G68), .ZN(new_n426));
  OAI21_X1  g0226(.A(G20), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT78), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n427), .B(new_n428), .C1(new_n422), .C2(new_n288), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n312), .A2(new_n233), .A3(new_n313), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT7), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n312), .A2(KEYINPUT7), .A3(new_n233), .A4(new_n313), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n203), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n419), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT7), .B1(new_n344), .B2(new_n233), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n315), .A2(new_n316), .A3(new_n432), .A4(G20), .ZN(new_n438));
  OAI21_X1  g0238(.A(G68), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(KEYINPUT16), .A3(new_n429), .A4(new_n424), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(new_n440), .A3(new_n260), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n265), .A2(new_n276), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n360), .B1(new_n281), .B2(new_n285), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n349), .A2(G223), .A3(new_n350), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n223), .A2(new_n347), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n344), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G87), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n287), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n319), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n303), .B1(new_n305), .B2(new_n225), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(G169), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n446), .B1(new_n309), .B2(G223), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n455), .A2(new_n344), .B1(new_n287), .B2(new_n449), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n452), .B1(new_n456), .B2(new_n319), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n367), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n418), .B1(new_n444), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n444), .A2(new_n458), .A3(new_n418), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G190), .ZN(new_n463));
  AND4_X1   g0263(.A1(KEYINPUT79), .A2(new_n451), .A3(new_n463), .A4(new_n453), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT79), .B1(new_n457), .B2(G200), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n457), .A2(new_n463), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT17), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(KEYINPUT80), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n467), .A2(new_n444), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n441), .A2(new_n443), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n457), .A2(KEYINPUT79), .A3(new_n463), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n451), .A2(new_n453), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(new_n322), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(G190), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n471), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  NOR4_X1   g0280(.A1(new_n371), .A2(new_n417), .A3(new_n462), .A4(new_n480), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n299), .A2(G1), .ZN(new_n483));
  INV_X1    g0283(.A(new_n232), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n301), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G264), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n275), .A2(G45), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G274), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n484), .B2(new_n301), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(G257), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G294), .ZN(new_n498));
  INV_X1    g0298(.A(G250), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n498), .C1(new_n351), .C2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT88), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n309), .A2(new_n310), .A3(G250), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(KEYINPUT88), .A3(new_n497), .A4(new_n498), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n302), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n496), .B1(new_n505), .B2(KEYINPUT89), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT89), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n507), .B(new_n302), .C1(new_n502), .C2(new_n504), .ZN(new_n508));
  OAI21_X1  g0308(.A(G169), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n502), .A2(new_n504), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(new_n319), .B1(G264), .B2(new_n485), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G179), .A3(new_n494), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT87), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n233), .B(G87), .C1(new_n315), .C2(new_n316), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT85), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n310), .A2(new_n517), .A3(new_n233), .A4(G87), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G107), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G20), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT86), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT23), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n522), .A2(KEYINPUT23), .B1(G20), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n523), .B1(new_n522), .B2(KEYINPUT23), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT22), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n515), .A2(KEYINPUT85), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n513), .B(new_n514), .C1(new_n520), .C2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n519), .A2(new_n529), .A3(KEYINPUT87), .A4(new_n531), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT24), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n527), .A2(new_n528), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n531), .A2(new_n536), .A3(new_n524), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT87), .B1(new_n537), .B2(new_n519), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n533), .B(new_n260), .C1(new_n535), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n281), .A2(KEYINPUT25), .A3(new_n521), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT25), .B1(new_n281), .B2(new_n521), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n275), .A2(G33), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n261), .A2(new_n279), .A3(new_n543), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n541), .A2(new_n542), .B1(new_n544), .B2(new_n521), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n509), .A2(new_n512), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n261), .B1(new_n538), .B2(new_n514), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n513), .B1(new_n520), .B2(new_n532), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(KEYINPUT24), .A3(new_n534), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n545), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n510), .A2(new_n319), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n495), .B1(new_n552), .B2(new_n507), .ZN(new_n553));
  INV_X1    g0353(.A(new_n508), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n463), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n494), .A3(new_n486), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n322), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n547), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(KEYINPUT4), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n351), .B2(new_n219), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G283), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n347), .B1(new_n312), .B2(new_n313), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(G250), .ZN(new_n566));
  INV_X1    g0366(.A(new_n561), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n309), .A2(new_n310), .A3(new_n567), .A4(G244), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n562), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT82), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT82), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n562), .A2(new_n566), .A3(new_n571), .A4(new_n568), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n319), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n485), .A2(G257), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n574), .A2(new_n494), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n367), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT6), .ZN(new_n577));
  INV_X1    g0377(.A(G97), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n577), .A2(new_n578), .A3(G107), .ZN(new_n579));
  XNOR2_X1  g0379(.A(G97), .B(G107), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n579), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n581), .A2(new_n233), .B1(new_n204), .B2(new_n288), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n521), .B1(new_n433), .B2(new_n434), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n260), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n279), .A2(G97), .ZN(new_n585));
  INV_X1    g0385(.A(new_n544), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n585), .B1(new_n586), .B2(G97), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n573), .A2(new_n575), .ZN(new_n590));
  INV_X1    g0390(.A(G169), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n575), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n302), .B1(new_n569), .B2(KEYINPUT82), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(new_n572), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n588), .B1(new_n595), .B2(G190), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n590), .A2(G200), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n576), .A2(new_n592), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n360), .A2(G116), .A3(new_n543), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n281), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n259), .A2(new_n232), .B1(G20), .B2(new_n600), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n563), .B(new_n233), .C1(G33), .C2(new_n578), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n602), .A2(KEYINPUT20), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT20), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n599), .B(new_n601), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(G264), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n312), .A2(G303), .A3(new_n313), .ZN(new_n609));
  OAI21_X1  g0409(.A(G257), .B1(new_n315), .B2(new_n316), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n349), .A2(new_n350), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n319), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n485), .A2(G270), .B1(new_n493), .B2(new_n491), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n607), .B(KEYINPUT84), .C1(new_n615), .C2(new_n322), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n322), .B1(new_n613), .B2(new_n614), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n606), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(G190), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n616), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT19), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n375), .B2(new_n377), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n623), .A2(G20), .B1(G87), .B2(new_n208), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT83), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n625), .B(new_n622), .C1(new_n266), .C2(new_n578), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n310), .A2(new_n233), .A3(G68), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n622), .B1(new_n266), .B2(new_n578), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT83), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n624), .A2(new_n626), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n630), .A2(new_n260), .B1(new_n281), .B2(new_n355), .ZN(new_n631));
  OAI211_X1 g0431(.A(G244), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n632), .B(new_n526), .C1(new_n346), .C2(new_n611), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n319), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n483), .A2(G250), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n319), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(G274), .B2(new_n487), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G200), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n634), .A2(G190), .A3(new_n637), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n586), .A2(G87), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n631), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n378), .A2(KEYINPUT19), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n233), .B1(new_n449), .B2(new_n207), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n629), .A2(new_n627), .A3(new_n626), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n260), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n355), .A2(new_n281), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n586), .A2(new_n356), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n638), .A2(new_n591), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n634), .A2(new_n367), .A3(new_n637), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n613), .A2(new_n614), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(G169), .A3(new_n606), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT21), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n654), .A2(new_n606), .A3(KEYINPUT21), .A4(G169), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n613), .A2(new_n614), .A3(G179), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n606), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n621), .A2(new_n653), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n598), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n481), .A2(new_n559), .A3(new_n663), .ZN(G372));
  AND3_X1   g0464(.A1(new_n444), .A2(new_n418), .A3(new_n458), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(new_n459), .ZN(new_n666));
  INV_X1    g0466(.A(new_n412), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n416), .B2(new_n369), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n666), .B1(new_n668), .B2(new_n480), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT92), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n338), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g0471(.A(KEYINPUT92), .B(new_n327), .C1(new_n336), .C2(new_n337), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n341), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n576), .B(new_n588), .C1(new_n595), .C2(G169), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n675), .B2(new_n653), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n633), .A2(KEYINPUT90), .A3(new_n319), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT90), .B1(new_n633), .B2(new_n319), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n637), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n591), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT91), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n649), .A2(new_n651), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(KEYINPUT91), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n506), .A2(G190), .A3(new_n508), .ZN(new_n686));
  AOI21_X1  g0486(.A(G200), .B1(new_n511), .B2(new_n494), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n551), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n596), .A2(new_n597), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n509), .A2(new_n512), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n539), .A2(new_n546), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n661), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n675), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n631), .A2(new_n641), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n679), .A2(G200), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n695), .A2(new_n640), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(KEYINPUT26), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n685), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n481), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n674), .A2(new_n701), .ZN(G369));
  NAND3_X1  g0502(.A1(new_n275), .A2(new_n233), .A3(G13), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G213), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G343), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n559), .B1(new_n551), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n547), .A2(new_n708), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n621), .A2(new_n661), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n607), .A2(new_n709), .ZN(new_n714));
  MUX2_X1   g0514(.A(new_n713), .B(new_n661), .S(new_n714), .Z(new_n715));
  AND2_X1   g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n661), .A2(new_n709), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n559), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n547), .A2(new_n709), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n717), .A2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n212), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n230), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  INV_X1    g0529(.A(G330), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  INV_X1    g0531(.A(new_n638), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n552), .A2(new_n486), .A3(new_n659), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(new_n733), .B2(new_n590), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n654), .A2(new_n638), .A3(new_n367), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n595), .A2(new_n735), .A3(new_n511), .A4(KEYINPUT30), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n679), .A2(KEYINPUT93), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT93), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n739), .B(new_n637), .C1(new_n677), .C2(new_n678), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n590), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n615), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n556), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n708), .B1(new_n737), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(KEYINPUT31), .B(new_n708), .C1(new_n737), .C2(new_n744), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n663), .A2(new_n559), .A3(new_n709), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n730), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT29), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n699), .B2(new_n708), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT94), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n697), .B1(new_n558), .B2(new_n551), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n756), .B(new_n598), .C1(new_n547), .C2(new_n661), .ZN(new_n757));
  INV_X1    g0557(.A(new_n684), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n695), .A2(new_n640), .A3(new_n696), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(new_n592), .A3(KEYINPUT26), .A4(new_n576), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT26), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n675), .B2(new_n653), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(KEYINPUT29), .A3(new_n709), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n755), .A2(new_n765), .ZN(new_n766));
  OAI211_X1 g0566(.A(KEYINPUT94), .B(new_n752), .C1(new_n699), .C2(new_n708), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n751), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n729), .B1(new_n768), .B2(G1), .ZN(G364));
  XNOR2_X1  g0569(.A(new_n716), .B(KEYINPUT95), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n233), .A2(G13), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT96), .Z(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G45), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G1), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n724), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n770), .B(new_n776), .C1(G330), .C2(new_n715), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n212), .A2(G355), .A3(new_n310), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G116), .B2(new_n212), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n252), .A2(G45), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n310), .B(new_n723), .C1(new_n299), .C2(new_n231), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n232), .B1(G20), .B2(new_n591), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n775), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n233), .A2(new_n367), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n791), .A2(G190), .A3(new_n322), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n463), .A2(G179), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n233), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G68), .A2(new_n792), .B1(new_n795), .B2(G97), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT99), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n233), .A2(G179), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT98), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(KEYINPUT98), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G87), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G190), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n790), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n310), .B1(new_n806), .B2(new_n204), .C1(new_n222), .C2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n798), .A2(new_n463), .A3(G200), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(G107), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n790), .A2(G190), .A3(new_n322), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT97), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT32), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n798), .A2(new_n805), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n422), .ZN(new_n816));
  INV_X1    g0616(.A(new_n815), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n817), .A2(KEYINPUT32), .A3(G159), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n813), .A2(G58), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n797), .A2(new_n804), .A3(new_n811), .A4(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G329), .ZN(new_n821));
  INV_X1    g0621(.A(G322), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n344), .B1(new_n815), .B2(new_n821), .C1(new_n812), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT101), .ZN(new_n824));
  XOR2_X1   g0624(.A(KEYINPUT33), .B(G317), .Z(new_n825));
  OAI21_X1  g0625(.A(new_n792), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n823), .B(new_n827), .C1(G283), .C2(new_n810), .ZN(new_n828));
  INV_X1    g0628(.A(G303), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n802), .ZN(new_n830));
  INV_X1    g0630(.A(new_n806), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n795), .A2(G294), .B1(new_n831), .B2(G311), .ZN(new_n832));
  INV_X1    g0632(.A(G326), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n807), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT100), .Z(new_n835));
  OAI21_X1  g0635(.A(new_n820), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n789), .B1(new_n836), .B2(new_n786), .ZN(new_n837));
  INV_X1    g0637(.A(new_n785), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n715), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n777), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  NOR2_X1   g0641(.A1(new_n786), .A2(new_n783), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n776), .B1(new_n204), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n786), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n310), .B1(new_n817), .B2(G311), .ZN(new_n845));
  INV_X1    g0645(.A(G294), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n600), .B2(new_n806), .C1(new_n846), .C2(new_n812), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n809), .A2(new_n449), .ZN(new_n848));
  INV_X1    g0648(.A(new_n807), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(G303), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G283), .ZN(new_n851));
  INV_X1    g0651(.A(new_n792), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n850), .B1(new_n578), .B2(new_n794), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n847), .B(new_n853), .C1(G107), .C2(new_n803), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n849), .A2(G137), .B1(new_n831), .B2(G159), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n286), .B2(new_n852), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G143), .B2(new_n813), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT34), .Z(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n310), .B1(new_n815), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G68), .B2(new_n810), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n861), .B1(new_n224), .B2(new_n794), .C1(new_n802), .C2(new_n222), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT102), .Z(new_n863));
  AOI21_X1  g0663(.A(new_n854), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n364), .B1(new_n363), .B2(new_n709), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n370), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n370), .A2(new_n708), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n843), .B1(new_n844), .B2(new_n864), .C1(new_n869), .C2(new_n784), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n699), .A2(new_n708), .B1(new_n868), .B2(new_n867), .ZN(new_n872));
  INV_X1    g0672(.A(new_n698), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n688), .B(new_n689), .C1(new_n547), .C2(new_n661), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n874), .B2(new_n675), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n709), .B(new_n869), .C1(new_n875), .C2(new_n685), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n751), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT103), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n775), .B1(new_n877), .B2(new_n878), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n871), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  INV_X1    g0683(.A(new_n581), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(G116), .A3(new_n234), .A4(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT36), .Z(new_n888));
  NAND3_X1  g0688(.A1(new_n231), .A2(G77), .A3(new_n420), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n222), .A2(G68), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n275), .B(G13), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AOI221_X4 g0692(.A(new_n392), .B1(new_n414), .B2(new_n415), .C1(new_n398), .C2(new_n400), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n411), .A2(new_n709), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT104), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n401), .A2(new_n416), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT104), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(new_n894), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n416), .B(new_n895), .C1(new_n401), .C2(new_n411), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n691), .A2(new_n692), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n598), .A2(new_n662), .A3(new_n902), .A4(new_n688), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n747), .B(new_n748), .C1(new_n903), .C2(new_n708), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT40), .A4(new_n869), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  INV_X1    g0707(.A(new_n706), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n444), .B1(new_n458), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n909), .B2(KEYINPUT105), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n472), .A2(new_n478), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n909), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n910), .B(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n472), .A2(new_n706), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n480), .B2(new_n462), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT106), .ZN(new_n919));
  INV_X1    g0719(.A(new_n914), .ZN(new_n920));
  INV_X1    g0720(.A(new_n471), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n467), .B2(new_n444), .ZN(new_n922));
  INV_X1    g0722(.A(new_n469), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n472), .A2(new_n478), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n920), .B1(new_n925), .B2(new_n666), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n467), .A2(new_n444), .ZN(new_n927));
  INV_X1    g0727(.A(new_n454), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(G179), .B2(new_n475), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n929), .A2(new_n706), .B1(new_n441), .B2(new_n443), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n907), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n911), .A2(KEYINPUT37), .A3(new_n909), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n919), .B1(new_n934), .B2(KEYINPUT38), .ZN(new_n935));
  NOR4_X1   g0735(.A1(new_n926), .A2(new_n933), .A3(KEYINPUT106), .A4(new_n917), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n918), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n932), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT37), .B1(new_n911), .B2(new_n909), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n915), .A2(KEYINPUT38), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n917), .B1(new_n926), .B2(new_n933), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n943), .A2(new_n904), .A3(new_n869), .A4(new_n901), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT40), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n906), .A2(new_n937), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n946), .A2(new_n481), .A3(new_n904), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n946), .B1(new_n481), .B2(new_n904), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n947), .A2(new_n948), .A3(new_n730), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT38), .B1(new_n915), .B2(new_n940), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n926), .A2(new_n933), .A3(new_n917), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT39), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n412), .A2(new_n708), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n919), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n941), .A2(KEYINPUT106), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n955), .A2(new_n956), .B1(new_n917), .B2(new_n916), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n953), .B(new_n954), .C1(new_n957), .C2(KEYINPUT39), .ZN(new_n958));
  INV_X1    g0758(.A(new_n868), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n876), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n943), .A3(new_n901), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n462), .A2(new_n706), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n755), .A2(new_n481), .A3(new_n767), .A4(new_n765), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n674), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n963), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n949), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n275), .B2(new_n772), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n949), .A2(new_n966), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n892), .B1(new_n968), .B2(new_n969), .ZN(G367));
  OAI21_X1  g0770(.A(new_n787), .B1(new_n212), .B2(new_n355), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n723), .A2(new_n310), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n971), .B1(new_n972), .B2(new_n245), .ZN(new_n973));
  INV_X1    g0773(.A(G137), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n806), .A2(new_n222), .B1(new_n815), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n812), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n344), .B(new_n975), .C1(G150), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n803), .A2(G58), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n795), .A2(G68), .B1(new_n810), .B2(G77), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n792), .A2(G159), .B1(new_n849), .B2(G143), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n802), .A2(new_n600), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT46), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n813), .A2(G303), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G107), .A2(new_n795), .B1(new_n849), .B2(G311), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n792), .A2(G294), .B1(G97), .B2(new_n810), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n344), .B1(new_n806), .B2(new_n851), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G317), .B2(new_n817), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n981), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT47), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n776), .B(new_n973), .C1(new_n991), .C2(new_n786), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n695), .A2(new_n709), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n758), .B1(new_n995), .B2(new_n759), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n758), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n992), .B1(new_n997), .B2(new_n838), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n598), .B1(new_n589), .B2(new_n709), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT109), .B1(new_n675), .B2(new_n709), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT109), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n592), .A2(new_n1001), .A3(new_n576), .A4(new_n708), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n675), .B1(new_n1005), .B2(new_n902), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n709), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT42), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n1005), .B2(new_n719), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1004), .A2(KEYINPUT42), .A3(new_n559), .A4(new_n718), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n997), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1007), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT110), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1009), .A2(new_n1010), .B1(new_n1006), .B2(new_n709), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT110), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n1017), .A3(new_n1013), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1016), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1013), .B1(KEYINPUT43), .B2(new_n997), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AND3_X1   g0822(.A1(new_n1019), .A2(KEYINPUT111), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(KEYINPUT111), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1023), .A2(new_n1024), .B1(new_n717), .B2(new_n1005), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT111), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n717), .A2(new_n1005), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1019), .A2(KEYINPUT111), .A3(new_n1022), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n721), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT45), .B1(new_n721), .B2(new_n1004), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n719), .A2(new_n720), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1035), .A2(new_n1005), .A3(KEYINPUT44), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT44), .B1(new_n1035), .B2(new_n1005), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1033), .A2(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n717), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n712), .A2(new_n718), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n719), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n770), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n716), .A3(new_n719), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n768), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n724), .B(KEYINPUT41), .Z(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n774), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n998), .B1(new_n1032), .B2(new_n1049), .ZN(G387));
  INV_X1    g0850(.A(new_n1045), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n710), .A2(new_n711), .A3(new_n785), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n242), .A2(G45), .A3(new_n344), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n285), .B2(G50), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n265), .A2(KEYINPUT50), .A3(new_n222), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n247), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n726), .B1(new_n1057), .B2(new_n310), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n723), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n787), .B1(new_n212), .B2(new_n521), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n775), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n807), .A2(new_n422), .B1(new_n809), .B2(new_n578), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n310), .B1(new_n815), .B2(new_n286), .C1(new_n806), .C2(new_n203), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n265), .C2(new_n792), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n794), .A2(new_n355), .B1(new_n812), .B2(new_n222), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT112), .Z(new_n1066));
  NAND2_X1  g0866(.A1(new_n803), .A2(G77), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n802), .A2(new_n846), .B1(new_n851), .B2(new_n794), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n792), .A2(G311), .B1(G303), .B2(new_n831), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n822), .B2(new_n807), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G317), .B2(new_n813), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1069), .B1(new_n1072), .B2(KEYINPUT48), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT113), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(KEYINPUT48), .B2(new_n1072), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT49), .Z(new_n1076));
  OAI221_X1 g0876(.A(new_n344), .B1(new_n815), .B2(new_n833), .C1(new_n809), .C2(new_n600), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1068), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1061), .B1(new_n1078), .B2(new_n786), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1051), .A2(new_n774), .B1(new_n1052), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n768), .A2(new_n1051), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n724), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n768), .A2(new_n1051), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(G393));
  XNOR2_X1  g0884(.A(new_n1038), .B(new_n717), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n774), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n812), .A2(new_n422), .B1(new_n807), .B2(new_n286), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n794), .A2(new_n204), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n848), .B(new_n1089), .C1(G50), .C2(new_n792), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n803), .A2(G68), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n344), .B1(new_n817), .B2(G143), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n285), .B2(new_n806), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .A4(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n802), .A2(new_n851), .B1(new_n822), .B2(new_n815), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1096), .A2(KEYINPUT115), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(KEYINPUT115), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n310), .B1(new_n810), .B2(G107), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT116), .ZN(new_n1101));
  INV_X1    g0901(.A(G311), .ZN(new_n1102));
  INV_X1    g0902(.A(G317), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n812), .A2(new_n1102), .B1(new_n807), .B2(new_n1103), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n792), .A2(G303), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n795), .A2(G116), .B1(new_n831), .B2(G294), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1095), .B1(new_n1101), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n786), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n256), .A2(new_n972), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n788), .B1(new_n723), .B2(G97), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n776), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1112), .B(new_n1115), .C1(new_n1004), .C2(new_n838), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n724), .B1(new_n1081), .B2(new_n1040), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1085), .B1(new_n768), .B2(new_n1051), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1086), .B(new_n1116), .C1(new_n1117), .C2(new_n1118), .ZN(G390));
  INV_X1    g0919(.A(KEYINPUT39), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n943), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n937), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(new_n784), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n776), .B1(new_n285), .B2(new_n842), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1089), .B1(G68), .B2(new_n810), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1125), .B1(new_n521), .B2(new_n852), .C1(new_n851), .C2(new_n807), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n344), .B1(new_n812), .B2(new_n600), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n806), .A2(new_n578), .B1(new_n815), .B2(new_n846), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n802), .A2(new_n286), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT53), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT54), .B(G143), .Z(new_n1132));
  AOI22_X1  g0932(.A1(new_n831), .A2(new_n1132), .B1(new_n817), .B2(G125), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1133), .B(new_n310), .C1(new_n859), .C2(new_n812), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n852), .A2(new_n974), .B1(new_n222), .B2(new_n809), .ZN(new_n1135));
  INV_X1    g0935(.A(G128), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n794), .A2(new_n422), .B1(new_n807), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1129), .A2(new_n804), .B1(new_n1131), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1124), .B1(new_n1139), .B2(new_n844), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1123), .A2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n708), .B(new_n867), .C1(new_n757), .C2(new_n763), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n901), .B1(new_n1142), .B2(new_n868), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n954), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n937), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n954), .B1(new_n960), .B2(new_n901), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1122), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n904), .A2(G330), .A3(new_n869), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n901), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1150), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1145), .B(new_n1152), .C1(new_n1122), .C2(new_n1146), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n774), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT118), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT118), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1151), .A2(new_n1156), .A3(new_n774), .A4(new_n1153), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1141), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n481), .A2(new_n751), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n964), .A2(new_n674), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n960), .B1(new_n1163), .B2(new_n1150), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1142), .A2(new_n868), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1152), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1159), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1151), .A2(new_n1153), .A3(new_n1161), .A4(new_n1167), .ZN(new_n1170));
  AND4_X1   g0970(.A1(KEYINPUT117), .A2(new_n1169), .A3(new_n724), .A4(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n725), .B1(new_n1159), .B2(new_n1168), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT117), .B1(new_n1172), .B2(new_n1170), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1158), .B1(new_n1171), .B2(new_n1173), .ZN(G378));
  NAND3_X1  g0974(.A1(new_n671), .A2(new_n672), .A3(new_n342), .ZN(new_n1175));
  XOR2_X1   g0975(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1176), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n671), .A2(new_n672), .A3(new_n342), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n284), .A2(new_n292), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n908), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1182), .B(new_n1183), .Z(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1177), .A2(new_n1179), .A3(new_n1184), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n946), .B2(G330), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n901), .A2(new_n904), .A3(new_n869), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n945), .B1(new_n1190), .B2(new_n952), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1191), .B(G330), .C1(new_n957), .C2(new_n905), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1177), .A2(new_n1179), .A3(new_n1184), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1184), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n963), .B1(new_n1189), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT123), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1188), .A2(new_n946), .A3(G330), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1197), .A2(new_n1198), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1170), .A2(new_n1161), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(KEYINPUT123), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n725), .B1(new_n1209), .B2(new_n1204), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1203), .A2(new_n774), .A3(new_n1205), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G33), .A2(G41), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G50), .B(new_n1213), .C1(new_n344), .C2(new_n298), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n852), .A2(new_n578), .B1(new_n224), .B2(new_n809), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n344), .B(new_n298), .C1(new_n815), .C2(new_n851), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n812), .A2(new_n521), .B1(new_n806), .B2(new_n355), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n794), .A2(new_n203), .B1(new_n807), .B2(new_n600), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT119), .Z(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1220), .A3(new_n1067), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1214), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n803), .A2(new_n1132), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n812), .A2(new_n1136), .B1(new_n806), .B2(new_n974), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G150), .B2(new_n795), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n792), .A2(G132), .B1(new_n849), .B2(G125), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1228), .B(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(G124), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1213), .B1(new_n815), .B2(new_n1231), .C1(new_n809), .C2(new_n422), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1223), .B1(new_n1222), .B2(new_n1221), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n786), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n842), .A2(new_n222), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n775), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1195), .B2(new_n783), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1212), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1211), .A2(new_n1238), .ZN(G375));
  NAND2_X1  g1039(.A1(new_n813), .A2(G137), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G132), .A2(new_n849), .B1(new_n810), .B2(G58), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n792), .A2(new_n1132), .B1(new_n795), .B2(G50), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n310), .B1(new_n806), .B2(new_n286), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G128), .B2(new_n817), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n802), .A2(new_n422), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n802), .A2(new_n578), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n792), .A2(G116), .B1(new_n849), .B2(G294), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n795), .A2(new_n356), .B1(new_n810), .B2(G77), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n310), .B1(new_n976), .B2(G283), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G107), .A2(new_n831), .B1(new_n817), .B2(G303), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1245), .A2(new_n1246), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n786), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n776), .B1(new_n203), .B2(new_n842), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(new_n901), .C2(new_n784), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n774), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1168), .A2(new_n1048), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n964), .A2(new_n674), .A3(new_n1160), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1259), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(G381));
  NOR4_X1   g1065(.A1(G390), .A2(G396), .A3(G393), .A4(G384), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1264), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1172), .A2(new_n1170), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1158), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OR4_X1    g1070(.A1(G387), .A2(new_n1267), .A3(G375), .A4(new_n1270), .ZN(G407));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n707), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G375), .C2(new_n1272), .ZN(G409));
  NAND3_X1  g1073(.A1(new_n1211), .A2(G378), .A3(new_n1238), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1197), .A2(new_n1202), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1237), .B1(new_n1275), .B2(new_n774), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1206), .B2(new_n1047), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1269), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G213), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(G343), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1257), .A2(KEYINPUT60), .A3(new_n1262), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1283), .A2(new_n724), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1168), .A2(KEYINPUT60), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1263), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1259), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(G384), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1259), .B(new_n882), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1279), .A2(KEYINPUT63), .A3(new_n1282), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT125), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1281), .B1(new_n1274), .B2(new_n1278), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(KEYINPUT63), .A4(new_n1290), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1287), .A2(G384), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1289), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1281), .A2(G2897), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G2897), .B(new_n1281), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1297), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(G390), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT124), .B1(G387), .B2(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(G393), .B(new_n840), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n766), .A2(new_n767), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n878), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n1085), .B2(new_n1051), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1258), .B1(new_n1312), .B2(new_n1047), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(new_n1031), .A3(new_n1025), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(new_n998), .A3(G390), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G390), .B1(new_n1314), .B2(new_n998), .ZN(new_n1317));
  OAI22_X1  g1117(.A1(new_n1307), .A2(new_n1309), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1317), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1320), .A2(KEYINPUT124), .A3(new_n1315), .A4(new_n1308), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1318), .A2(new_n1319), .A3(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1279), .A2(new_n1282), .A3(new_n1290), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1305), .B(new_n1322), .C1(new_n1324), .C2(KEYINPUT63), .ZN(new_n1325));
  XOR2_X1   g1125(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n1293), .B2(new_n1303), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT62), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1323), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1293), .A2(KEYINPUT62), .A3(new_n1290), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1327), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1318), .A2(KEYINPUT127), .A3(new_n1321), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI22_X1  g1136(.A1(new_n1296), .A2(new_n1325), .B1(new_n1331), .B2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(G375), .A2(new_n1269), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1338), .B(new_n1274), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1270), .B1(new_n1211), .B2(new_n1238), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1211), .A2(G378), .A3(new_n1238), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1290), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1332), .ZN(G402));
endmodule


