//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(G43gat), .B(G50gat), .Z(new_n204));
  NOR2_X1   g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT89), .B(G36gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n204), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n205), .B(KEYINPUT14), .ZN(new_n213));
  INV_X1    g012(.A(new_n209), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n213), .B1(G29gat), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(KEYINPUT15), .A3(new_n204), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT17), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G1gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  MUX2_X1   g022(.A(G1gat), .B(new_n222), .S(new_n223), .Z(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(G8gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n225), .B(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n228), .A2(KEYINPUT91), .A3(new_n219), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT91), .B1(new_n228), .B2(new_n219), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n203), .B(new_n226), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT18), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n228), .A2(new_n219), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n228), .A2(new_n219), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(KEYINPUT91), .A3(new_n219), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n203), .B(KEYINPUT13), .Z(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT92), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT92), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n229), .A2(new_n230), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n242), .B(new_n239), .C1(new_n243), .C2(new_n233), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT11), .ZN(new_n247));
  INV_X1    g046(.A(G169gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G197gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n232), .A2(new_n245), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n232), .B2(new_n245), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n202), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n232), .A2(new_n245), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n251), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n232), .A2(new_n245), .A3(new_n252), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(KEYINPUT93), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G155gat), .B(G162gat), .ZN(new_n262));
  INV_X1    g061(.A(G141gat), .ZN(new_n263));
  INV_X1    g062(.A(G148gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G155gat), .ZN(new_n266));
  INV_X1    g065(.A(G162gat), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT2), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n262), .A2(new_n265), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n271), .A3(new_n269), .ZN(new_n272));
  AND2_X1   g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g077(.A(G134gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT67), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G134gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n282), .A3(G127gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n284));
  INV_X1    g083(.A(G127gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(G134gat), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G120gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G113gat), .ZN(new_n291));
  INV_X1    g090(.A(G113gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G120gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n294), .A2(new_n298), .A3(new_n295), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(KEYINPUT75), .B(KEYINPUT3), .Z(new_n301));
  NAND3_X1  g100(.A1(new_n270), .A2(new_n276), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n278), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n297), .A2(new_n276), .A3(new_n270), .A4(new_n299), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT4), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n283), .A2(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n294), .A2(new_n298), .A3(new_n295), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n270), .A2(new_n276), .ZN(new_n312));
  XOR2_X1   g111(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n313));
  NAND4_X1  g112(.A1(new_n311), .A2(KEYINPUT78), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n277), .A2(new_n309), .A3(new_n310), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT78), .B1(new_n316), .B2(new_n313), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n303), .B(new_n306), .C1(new_n315), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n307), .A2(new_n313), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n311), .A2(KEYINPUT4), .A3(new_n312), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n319), .A2(new_n303), .A3(new_n304), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT5), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n277), .B1(new_n309), .B2(new_n310), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n324), .B2(new_n305), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT0), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT77), .ZN(new_n329));
  XOR2_X1   g128(.A(G57gat), .B(G85gat), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n328), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n330), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n326), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT6), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT79), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n318), .A2(new_n326), .ZN(new_n341));
  INV_X1    g140(.A(new_n336), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(new_n346), .A3(new_n338), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n336), .B1(new_n318), .B2(new_n326), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT80), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n340), .A2(new_n345), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT81), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n348), .B(new_n344), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n340), .A4(new_n347), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n341), .A2(KEYINPUT6), .A3(new_n342), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G22gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  AND2_X1   g157(.A1(G211gat), .A2(G218gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(G211gat), .A2(G218gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n363));
  INV_X1    g162(.A(G197gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(G204gat), .ZN(new_n365));
  INV_X1    g164(.A(G204gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(G197gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(G197gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n364), .A2(G204gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT70), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n359), .A2(KEYINPUT22), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n362), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  AOI211_X1 g174(.A(new_n361), .B(new_n373), .C1(new_n368), .C2(new_n371), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n358), .B(new_n277), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n302), .A2(new_n358), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n372), .A2(new_n362), .A3(new_n374), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT70), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT70), .B1(new_n369), .B2(new_n370), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n361), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n378), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G228gat), .ZN(new_n385));
  INV_X1    g184(.A(G233gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n278), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n377), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n358), .B1(new_n375), .B2(new_n376), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n301), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n391), .A2(new_n277), .B1(new_n392), .B2(new_n378), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n357), .B(new_n389), .C1(new_n393), .C2(new_n387), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n383), .B2(new_n379), .ZN(new_n395));
  INV_X1    g194(.A(new_n301), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n277), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n387), .B1(new_n397), .B2(new_n384), .ZN(new_n398));
  INV_X1    g197(.A(new_n389), .ZN(new_n399));
  OAI21_X1  g198(.A(G22gat), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XOR2_X1   g202(.A(G78gat), .B(G106gat), .Z(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT82), .ZN(new_n405));
  XOR2_X1   g204(.A(KEYINPUT31), .B(G50gat), .Z(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n401), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n407), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n394), .B(new_n400), .C1(new_n402), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT23), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n414), .A2(G169gat), .A3(G176gat), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n415), .B2(KEYINPUT64), .ZN(new_n416));
  INV_X1    g215(.A(G176gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n248), .A2(new_n417), .A3(KEYINPUT23), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT23), .B1(new_n248), .B2(new_n417), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT64), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(G183gat), .A2(G190gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n416), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT25), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n414), .B1(G169gat), .B2(G176gat), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n418), .A2(new_n430), .A3(KEYINPUT25), .A4(new_n412), .ZN(new_n431));
  AND3_X1   g230(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n423), .B2(new_n422), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n423), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT65), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT26), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(new_n248), .A3(new_n417), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n413), .B1(new_n443), .B2(KEYINPUT65), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n437), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(G183gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT27), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT27), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G183gat), .ZN(new_n449));
  INV_X1    g248(.A(G190gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT28), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT27), .B(G183gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(KEYINPUT28), .A3(new_n450), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n445), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n445), .B2(new_n456), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n436), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n300), .ZN(new_n461));
  INV_X1    g260(.A(G227gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n386), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n436), .B(new_n311), .C1(new_n458), .C2(new_n459), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT34), .ZN(new_n467));
  XOR2_X1   g266(.A(G15gat), .B(G43gat), .Z(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n464), .B1(new_n461), .B2(new_n465), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n470), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n465), .ZN(new_n478));
  AOI221_X4 g277(.A(new_n475), .B1(new_n473), .B2(new_n470), .C1(new_n478), .C2(new_n463), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n467), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n463), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT32), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n472), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n470), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT34), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n466), .B(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n474), .A2(new_n476), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n411), .A2(new_n480), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G226gat), .A2(G233gat), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n460), .B2(new_n358), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n445), .A2(new_n456), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n412), .B1(new_n418), .B2(new_n420), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n433), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT25), .B1(new_n495), .B2(new_n421), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n496), .B2(new_n434), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n497), .A2(KEYINPUT72), .A3(new_n491), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT72), .B1(new_n497), .B2(new_n491), .ZN(new_n499));
  OAI22_X1  g298(.A1(new_n492), .A2(KEYINPUT71), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n434), .B1(new_n427), .B2(new_n428), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n493), .A2(KEYINPUT66), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n445), .A2(new_n456), .A3(new_n457), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n490), .B1(new_n504), .B2(KEYINPUT29), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT71), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n392), .B1(new_n500), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT29), .B1(new_n436), .B2(new_n493), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT73), .B1(new_n509), .B2(new_n491), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT73), .ZN(new_n511));
  INV_X1    g310(.A(new_n493), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(new_n501), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n511), .B(new_n490), .C1(new_n513), .C2(KEYINPUT29), .ZN(new_n514));
  INV_X1    g313(.A(new_n392), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n460), .A2(new_n491), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n510), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G8gat), .B(G36gat), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT74), .ZN(new_n519));
  XOR2_X1   g318(.A(G64gat), .B(G92gat), .Z(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AND4_X1   g320(.A1(KEYINPUT30), .A2(new_n508), .A3(new_n517), .A4(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n517), .ZN(new_n523));
  INV_X1    g322(.A(new_n499), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n497), .A2(KEYINPUT72), .A3(new_n491), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n505), .A2(new_n506), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n523), .B1(new_n529), .B2(new_n392), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT30), .B1(new_n530), .B2(new_n521), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n508), .A2(new_n517), .A3(new_n521), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n522), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n356), .A2(new_n489), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n411), .A2(new_n480), .A3(new_n488), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n343), .A2(new_n338), .A3(new_n337), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n355), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n348), .A2(KEYINPUT87), .A3(KEYINPUT6), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n534), .A2(KEYINPUT35), .B1(new_n533), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT37), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n508), .A2(new_n545), .A3(new_n517), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n510), .A2(new_n514), .A3(new_n392), .A4(new_n516), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n547), .A2(KEYINPUT37), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n515), .B1(new_n500), .B2(new_n507), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n521), .A2(KEYINPUT38), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n546), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n532), .A2(new_n539), .A3(new_n536), .A4(new_n538), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT88), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n546), .A2(new_n550), .A3(new_n551), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n532), .ZN(new_n558));
  INV_X1    g357(.A(new_n521), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n546), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n530), .A2(new_n545), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT38), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n554), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT86), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n521), .B1(new_n508), .B2(new_n517), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n532), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n508), .A2(new_n517), .A3(new_n521), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT30), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT85), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT40), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n573));
  INV_X1    g372(.A(new_n313), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n307), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(new_n314), .A3(new_n308), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n304), .B1(new_n576), .B2(new_n303), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT39), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n307), .A2(new_n323), .A3(new_n304), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(KEYINPUT84), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(KEYINPUT84), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n336), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n577), .A2(new_n578), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n572), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n577), .A2(new_n581), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n577), .A2(new_n578), .ZN(new_n586));
  INV_X1    g385(.A(new_n572), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n585), .A2(new_n336), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(new_n588), .A3(new_n343), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n564), .B1(new_n570), .B2(new_n590), .ZN(new_n591));
  AOI211_X1 g390(.A(KEYINPUT86), .B(new_n589), .C1(new_n567), .C2(new_n569), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n563), .B(new_n411), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n486), .B1(new_n484), .B2(new_n487), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n477), .A2(new_n467), .A3(new_n479), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT36), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n480), .A2(new_n488), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n356), .A2(new_n533), .ZN(new_n600));
  INV_X1    g399(.A(new_n411), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n544), .B1(new_n593), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n261), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT8), .ZN(new_n607));
  AND2_X1   g406(.A1(G99gat), .A2(G106gat), .ZN(new_n608));
  OAI221_X1 g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .C1(G85gat), .C2(G92gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(G99gat), .B(G106gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n220), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n219), .A2(new_n611), .B1(KEYINPUT41), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  NOR2_X1   g417(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n616), .B(new_n617), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(KEYINPUT41), .B2(new_n614), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G134gat), .B(G162gat), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G57gat), .B(G64gat), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G71gat), .B(G78gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G127gat), .B(G155gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n633), .B(KEYINPUT94), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n228), .B1(KEYINPUT21), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  XOR2_X1   g445(.A(G183gat), .B(G211gat), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n645), .B2(new_n646), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n611), .B(new_n633), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n642), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(G230gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n386), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n652), .A2(new_n659), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n660), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n658), .B1(new_n654), .B2(new_n655), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n668), .B2(new_n661), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n667), .A2(KEYINPUT95), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT95), .B1(new_n667), .B2(new_n669), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n628), .A2(new_n651), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n604), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n356), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  INV_X1    g476(.A(new_n674), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n533), .ZN(new_n679));
  INV_X1    g478(.A(G8gat), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT42), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  MUX2_X1   g482(.A(KEYINPUT42), .B(new_n681), .S(new_n683), .Z(G1325gat));
  NOR2_X1   g483(.A1(new_n594), .A2(new_n595), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n678), .A2(G15gat), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G15gat), .B1(new_n678), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n601), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  AND3_X1   g494(.A1(new_n620), .A2(new_n622), .A3(new_n626), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n626), .B1(new_n620), .B2(new_n622), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n672), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n651), .A2(new_n699), .ZN(new_n700));
  NOR4_X1   g499(.A1(new_n261), .A2(new_n603), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n208), .A3(new_n675), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n543), .A2(new_n533), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT97), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n591), .A2(new_n592), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n558), .A2(new_n562), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n540), .A2(new_n568), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n557), .B1(new_n711), .B2(new_n555), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n411), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n602), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n544), .A2(KEYINPUT97), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n708), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT98), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .A4(new_n628), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT44), .B1(new_n603), .B2(new_n698), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n593), .A2(new_n602), .B1(new_n544), .B2(KEYINPUT97), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n698), .B1(new_n722), .B2(new_n708), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n717), .B1(new_n723), .B2(new_n718), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n257), .A2(new_n258), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n725), .A2(new_n727), .A3(new_n700), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n675), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n703), .B1(new_n730), .B2(new_n208), .ZN(G1328gat));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n570), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n214), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n701), .A2(new_n570), .A3(new_n209), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT99), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n733), .B(new_n737), .C1(new_n735), .C2(new_n734), .ZN(G1329gat));
  INV_X1    g537(.A(G43gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n701), .A2(new_n739), .A3(new_n685), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT101), .Z(new_n741));
  INV_X1    g540(.A(new_n690), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n700), .A2(new_n727), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n742), .B(new_n743), .C1(new_n721), .C2(new_n724), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n744), .A2(KEYINPUT100), .A3(G43gat), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT100), .B1(new_n744), .B2(G43gat), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n741), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n739), .B1(new_n728), .B2(new_n599), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n740), .A2(KEYINPUT47), .ZN(new_n749));
  OAI22_X1  g548(.A1(new_n747), .A2(KEYINPUT47), .B1(new_n748), .B2(new_n749), .ZN(G1330gat));
  NAND3_X1  g549(.A1(new_n728), .A2(G50gat), .A3(new_n601), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n701), .A2(new_n601), .ZN(new_n752));
  INV_X1    g551(.A(G50gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n751), .A2(KEYINPUT48), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT48), .B1(new_n751), .B2(new_n754), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(G1331gat));
  INV_X1    g556(.A(new_n651), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n727), .A2(new_n758), .A3(new_n698), .A4(new_n672), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n708), .B2(new_n722), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n675), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g561(.A(new_n570), .B(KEYINPUT102), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  AND2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n766), .B2(new_n765), .ZN(G1333gat));
  AOI21_X1  g568(.A(G71gat), .B1(new_n760), .B2(new_n685), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n742), .A2(G71gat), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n760), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT103), .B(KEYINPUT50), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n760), .A2(new_n601), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g575(.A1(new_n758), .A2(new_n726), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n716), .A2(KEYINPUT51), .A3(new_n628), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT104), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT104), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n723), .A2(new_n780), .A3(KEYINPUT51), .A4(new_n777), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n716), .A2(new_n628), .A3(new_n777), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n779), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(G85gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n785), .A2(new_n786), .A3(new_n675), .A4(new_n672), .ZN(new_n787));
  INV_X1    g586(.A(new_n777), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n725), .A2(new_n699), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n675), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n787), .B1(new_n791), .B2(new_n786), .ZN(G1336gat));
  INV_X1    g591(.A(G92gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n789), .B2(new_n570), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n784), .A2(new_n778), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n763), .A2(G92gat), .A3(new_n699), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(KEYINPUT106), .B(KEYINPUT52), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n788), .A2(new_n699), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n764), .B(new_n800), .C1(new_n721), .C2(new_n724), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n799), .B1(new_n801), .B2(G92gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT107), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT105), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n785), .A2(new_n804), .A3(new_n796), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n785), .B2(new_n796), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n802), .B(new_n803), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n785), .A2(new_n796), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT105), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n805), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n803), .B1(new_n812), .B2(new_n802), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n798), .B1(new_n809), .B2(new_n813), .ZN(G1337gat));
  NOR2_X1   g613(.A1(new_n686), .A2(G99gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n785), .A2(new_n672), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n789), .A2(new_n742), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G99gat), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n817), .A2(new_n818), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n816), .B1(new_n820), .B2(new_n821), .ZN(G1338gat));
  NAND2_X1  g621(.A1(new_n789), .A2(new_n601), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n699), .A2(G106gat), .A3(new_n411), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT53), .B1(new_n785), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n823), .A2(G106gat), .B1(new_n795), .B2(new_n825), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(G1339gat));
  NAND3_X1  g629(.A1(new_n654), .A2(new_n655), .A3(new_n658), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n660), .A2(KEYINPUT54), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n666), .B1(new_n668), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(KEYINPUT55), .A3(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n667), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n834), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n257), .B2(new_n258), .ZN(new_n841));
  INV_X1    g640(.A(new_n243), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n203), .B1(new_n842), .B2(new_n226), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n243), .A2(new_n233), .A3(new_n239), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n250), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n258), .A2(new_n672), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n698), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n839), .A2(new_n667), .A3(new_n835), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n628), .A2(new_n258), .A3(new_n845), .A4(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n758), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR4_X1   g650(.A1(new_n628), .A2(new_n726), .A3(new_n651), .A4(new_n672), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n356), .A3(new_n535), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n763), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n292), .A3(new_n726), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT109), .ZN(new_n859));
  INV_X1    g658(.A(new_n855), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n260), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n859), .B1(new_n861), .B2(G113gat), .ZN(new_n862));
  AOI211_X1 g661(.A(KEYINPUT109), .B(new_n292), .C1(new_n860), .C2(new_n260), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(G1340gat));
  NAND3_X1  g663(.A1(new_n857), .A2(new_n290), .A3(new_n672), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n672), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT111), .B1(new_n866), .B2(G120gat), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n868), .B(new_n290), .C1(new_n860), .C2(new_n672), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n865), .B1(new_n867), .B2(new_n869), .ZN(G1341gat));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n651), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n286), .A2(new_n287), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT112), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n871), .B(new_n873), .ZN(G1342gat));
  NOR2_X1   g673(.A1(new_n698), .A2(new_n570), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n854), .A2(new_n280), .A3(new_n282), .A4(new_n875), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT56), .Z(new_n877));
  OAI21_X1  g676(.A(G134gat), .B1(new_n855), .B2(new_n698), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1343gat));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT117), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n763), .A2(new_n675), .A3(new_n596), .A4(new_n598), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n411), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n836), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n889), .B1(new_n255), .B2(new_n259), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n698), .B1(new_n890), .B2(new_n847), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n758), .B1(new_n891), .B2(new_n850), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n884), .B1(new_n892), .B2(new_n852), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n883), .B1(new_n853), .B2(new_n411), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n882), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n263), .B1(new_n895), .B2(new_n726), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n881), .B1(new_n896), .B2(new_n880), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n898), .B(new_n675), .C1(new_n851), .C2(new_n852), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n690), .A2(new_n601), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n849), .B1(new_n253), .B2(new_n254), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n628), .B1(new_n903), .B2(new_n846), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n849), .B1(new_n696), .B2(new_n697), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n258), .A2(new_n845), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n651), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n852), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n898), .B1(new_n910), .B2(new_n675), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n902), .A2(new_n911), .A3(new_n764), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n260), .A2(new_n263), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT116), .Z(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n902), .A2(new_n911), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n916), .A2(new_n917), .A3(new_n763), .A4(new_n914), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n261), .B(new_n882), .C1(new_n893), .C2(new_n894), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n263), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n897), .A2(new_n915), .B1(new_n920), .B2(new_n880), .ZN(G1344gat));
  NAND3_X1  g720(.A1(new_n912), .A2(new_n264), .A3(new_n672), .ZN(new_n922));
  XNOR2_X1  g721(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n261), .A2(new_n673), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n883), .B(new_n601), .C1(new_n892), .C2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT57), .B1(new_n853), .B2(new_n411), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n672), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n882), .B(KEYINPUT119), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n923), .B1(new_n929), .B2(G148gat), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT59), .B(new_n264), .C1(new_n895), .C2(new_n672), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n922), .B1(new_n930), .B2(new_n931), .ZN(G1345gat));
  NAND3_X1  g731(.A1(new_n912), .A2(new_n266), .A3(new_n758), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n895), .A2(new_n758), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n266), .ZN(G1346gat));
  AOI21_X1  g734(.A(new_n267), .B1(new_n895), .B2(new_n628), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n875), .A2(new_n267), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n902), .A2(new_n911), .A3(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n939));
  OR3_X1    g738(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n936), .B2(new_n938), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1347gat));
  NOR2_X1   g741(.A1(new_n763), .A2(new_n535), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n910), .A2(new_n356), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n910), .A2(KEYINPUT121), .A3(new_n356), .A4(new_n943), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n726), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n248), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n356), .A2(new_n570), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n853), .A2(new_n535), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(G169gat), .A3(new_n260), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(G1348gat));
  NAND2_X1  g754(.A1(new_n951), .A2(new_n672), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G176gat), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n946), .A2(new_n417), .A3(new_n672), .A4(new_n947), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT123), .Z(G1349gat));
  NAND2_X1  g759(.A1(new_n951), .A2(new_n758), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT124), .B1(new_n961), .B2(G183gat), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n853), .A2(new_n675), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n963), .A2(new_n454), .A3(new_n758), .A4(new_n943), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g765(.A(new_n450), .B1(new_n951), .B2(new_n628), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT61), .Z(new_n968));
  NAND4_X1  g767(.A1(new_n946), .A2(new_n450), .A3(new_n628), .A4(new_n947), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1351gat));
  NOR2_X1   g769(.A1(new_n742), .A2(new_n950), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n925), .A2(new_n260), .A3(new_n926), .A4(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n364), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n974), .B1(new_n973), .B2(new_n972), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n900), .A2(new_n763), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n726), .A2(new_n364), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(G1352gat));
  NOR3_X1   g780(.A1(new_n979), .A2(G204gat), .A3(new_n699), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT62), .ZN(new_n983));
  INV_X1    g782(.A(new_n971), .ZN(new_n984));
  OAI21_X1  g783(.A(G204gat), .B1(new_n927), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1353gat));
  OR3_X1    g785(.A1(new_n979), .A2(G211gat), .A3(new_n651), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n925), .A2(new_n758), .A3(new_n926), .A4(new_n971), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  NAND4_X1  g790(.A1(new_n925), .A2(new_n628), .A3(new_n926), .A4(new_n971), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G218gat), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n698), .A2(G218gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n979), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(KEYINPUT127), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n997));
  OAI211_X1 g796(.A(new_n993), .B(new_n997), .C1(new_n979), .C2(new_n994), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n996), .A2(new_n998), .ZN(G1355gat));
endmodule


