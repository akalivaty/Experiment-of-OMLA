//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G58), .A3(G68), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n216), .B1(new_n203), .B2(new_n217), .C1(new_n206), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n209), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n209), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT66), .Z(new_n230));
  AOI21_X1  g0030(.A(new_n225), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n246), .B(KEYINPUT69), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n226), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G50), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n255), .A2(new_n256), .B1(new_n227), .B2(G68), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n227), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n203), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n253), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT11), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n261), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n253), .B1(new_n264), .B2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n266));
  OR3_X1    g0066(.A1(new_n266), .A2(KEYINPUT12), .A3(G68), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT12), .B1(new_n266), .B2(G68), .ZN(new_n268));
  AOI22_X1  g0068(.A1(G68), .A2(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n262), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT14), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G226), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(G1698), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n278), .B1(new_n273), .B2(new_n205), .C1(new_n279), .C2(new_n235), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n285), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(G238), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n283), .B1(new_n282), .B2(new_n289), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n271), .B(G169), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  INV_X1    g0094(.A(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n290), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n293), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n271), .B1(new_n296), .B2(G169), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n270), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n291), .A2(new_n292), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n270), .B1(new_n300), .B2(G190), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT73), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n296), .B2(G200), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n302), .B(G200), .C1(new_n291), .C2(new_n292), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n301), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n276), .A2(G222), .A3(new_n277), .ZN(new_n309));
  INV_X1    g0109(.A(G223), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n309), .B1(new_n203), .B2(new_n276), .C1(new_n279), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n281), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n286), .B1(G226), .B2(new_n288), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n254), .A2(G150), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G58), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT8), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n319), .B(new_n320), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n317), .B1(new_n321), .B2(new_n258), .C1(new_n202), .C2(new_n227), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n322), .A2(new_n253), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n265), .A2(G50), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(G50), .B2(new_n266), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT9), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n316), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n326), .A2(KEYINPUT9), .B1(new_n314), .B2(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT10), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n329), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT71), .B(G179), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n314), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  AOI211_X1 g0139(.A(new_n338), .B(new_n326), .C1(new_n339), .C2(new_n314), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n276), .A2(G232), .A3(new_n277), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT72), .B(G107), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n342), .B1(new_n344), .B2(new_n276), .C1(new_n279), .C2(new_n212), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n281), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n286), .B1(G244), .B2(new_n288), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G200), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n252), .A2(new_n226), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT8), .B(G58), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n354), .A2(new_n258), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n350), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n265), .A2(G77), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(G77), .B2(new_n266), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n349), .B(new_n359), .C1(new_n315), .C2(new_n348), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(new_n348), .B2(new_n339), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n346), .A2(new_n336), .A3(new_n347), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n308), .A2(new_n335), .A3(new_n341), .A4(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n286), .B1(G232), .B2(new_n288), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT74), .B(G33), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n274), .B1(new_n367), .B2(new_n272), .ZN(new_n368));
  MUX2_X1   g0168(.A(G223), .B(G226), .S(G1698), .Z(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(new_n369), .B1(G33), .B2(G87), .ZN(new_n370));
  INV_X1    g0170(.A(new_n281), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n372), .A2(KEYINPUT77), .A3(G190), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n368), .A2(new_n369), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n286), .ZN(new_n378));
  INV_X1    g0178(.A(new_n288), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n235), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n374), .B1(new_n381), .B2(new_n315), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n373), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n321), .A2(new_n265), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n321), .B2(new_n266), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n227), .B(new_n274), .C1(new_n367), .C2(new_n272), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT7), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT74), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(G33), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT3), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(new_n227), .A4(new_n274), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n389), .A2(G68), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G58), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n211), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n254), .A2(G159), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n350), .B1(new_n396), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n275), .A2(new_n227), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n394), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n390), .A2(G33), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n272), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(KEYINPUT3), .A2(G33), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n394), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n211), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n403), .B1(new_n414), .B2(new_n402), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n387), .B1(new_n405), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n385), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n385), .A2(KEYINPUT17), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(G68), .B1(new_n388), .B2(KEYINPUT7), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n408), .A2(new_n409), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n412), .B1(new_n424), .B2(KEYINPUT3), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n394), .B1(new_n425), .B2(new_n227), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n404), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n415), .A3(new_n253), .ZN(new_n428));
  INV_X1    g0228(.A(new_n387), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT75), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n416), .A2(KEYINPUT75), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n372), .A2(G169), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n372), .B2(new_n336), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT18), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT76), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n432), .A2(new_n433), .A3(new_n439), .A4(new_n435), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n437), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n422), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n365), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n371), .B(G250), .C1(G1), .C2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n281), .A2(new_n284), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n445), .A2(G1), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n272), .B1(new_n408), .B2(new_n409), .ZN(new_n452));
  OAI211_X1 g0252(.A(G238), .B(new_n277), .C1(new_n452), .C2(new_n412), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n424), .A2(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n368), .A2(G244), .A3(G1698), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n368), .A2(KEYINPUT79), .A3(G244), .A4(G1698), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n451), .B1(new_n460), .B2(new_n371), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n339), .ZN(new_n462));
  INV_X1    g0262(.A(new_n354), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n266), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n425), .A2(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G68), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT19), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n344), .A2(new_n213), .A3(new_n205), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n227), .B1(new_n273), .B2(new_n205), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n258), .A2(KEYINPUT19), .A3(new_n205), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n464), .B1(new_n472), .B2(new_n253), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n264), .A2(G33), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n350), .A2(new_n266), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n462), .B(new_n478), .C1(new_n337), .C2(new_n461), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n475), .A2(new_n213), .ZN(new_n480));
  AOI211_X1 g0280(.A(new_n464), .B(new_n480), .C1(new_n472), .C2(new_n253), .ZN(new_n481));
  OAI211_X1 g0281(.A(G190), .B(new_n451), .C1(new_n460), .C2(new_n371), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n458), .A2(new_n459), .ZN(new_n483));
  INV_X1    g0283(.A(new_n455), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n450), .B1(new_n485), .B2(new_n281), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n481), .B(new_n482), .C1(new_n486), .C2(new_n383), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n217), .A2(G1698), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT4), .B1(new_n368), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n276), .A2(KEYINPUT4), .A3(G244), .A4(new_n277), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n281), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT5), .B(G41), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n448), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n496), .A2(new_n284), .A3(new_n281), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n371), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(G257), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G169), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n336), .B2(new_n501), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT6), .B1(new_n207), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n507), .A2(new_n227), .B1(new_n203), .B2(new_n255), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n344), .B1(new_n411), .B2(new_n413), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n253), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n266), .A2(G97), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n476), .B2(G97), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT78), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n510), .A2(KEYINPUT78), .A3(new_n512), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n501), .A2(G190), .ZN(new_n518));
  AOI21_X1  g0318(.A(G200), .B1(new_n494), .B2(new_n500), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n516), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  AND4_X1   g0320(.A1(new_n479), .A2(new_n487), .A3(new_n514), .A4(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n498), .A2(new_n218), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n368), .A2(G250), .A3(new_n277), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n424), .A2(G294), .ZN(new_n524));
  OAI211_X1 g0324(.A(G257), .B(G1698), .C1(new_n452), .C2(new_n412), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n497), .B(new_n522), .C1(new_n526), .C2(new_n281), .ZN(new_n527));
  OR3_X1    g0327(.A1(new_n527), .A2(KEYINPUT84), .A3(G200), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT84), .B1(new_n527), .B2(G200), .ZN(new_n529));
  INV_X1    g0329(.A(new_n527), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n528), .B(new_n529), .C1(G190), .C2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n213), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n276), .A2(new_n227), .A3(G87), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n465), .A2(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT23), .B1(new_n343), .B2(new_n227), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n424), .A2(new_n227), .A3(G116), .ZN(new_n537));
  OR3_X1    g0337(.A1(new_n227), .A2(KEYINPUT23), .A3(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT24), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n539), .B(new_n540), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT24), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n535), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n350), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n266), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT25), .B1(new_n549), .B2(new_n206), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n476), .A2(G107), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n531), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n521), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n522), .B1(new_n526), .B2(new_n281), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n447), .A2(new_n448), .A3(new_n495), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n294), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(G169), .B2(new_n527), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n543), .A2(KEYINPUT24), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n546), .B1(new_n545), .B2(new_n535), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n253), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n564), .B2(new_n553), .ZN(new_n565));
  OAI211_X1 g0365(.A(G257), .B(new_n277), .C1(new_n452), .C2(new_n412), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT80), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT80), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n368), .A2(new_n568), .A3(G257), .A4(new_n277), .ZN(new_n569));
  INV_X1    g0369(.A(new_n276), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G303), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n368), .A2(G264), .A3(G1698), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n567), .A2(new_n569), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n281), .ZN(new_n574));
  INV_X1    g0374(.A(G270), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n559), .B1(new_n575), .B2(new_n498), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT82), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n491), .B(new_n227), .C1(G33), .C2(new_n205), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n253), .C1(new_n227), .C2(G116), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT20), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT81), .B1(new_n582), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n475), .A2(G116), .ZN(new_n587));
  INV_X1    g0387(.A(G116), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n266), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT81), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n582), .A2(new_n591), .A3(new_n583), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n578), .A2(G169), .A3(new_n580), .A4(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n576), .B1(new_n573), .B2(new_n281), .ZN(new_n596));
  OAI21_X1  g0396(.A(G169), .B1(new_n586), .B2(new_n593), .ZN(new_n597));
  OAI211_X1 g0397(.A(KEYINPUT82), .B(new_n579), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n294), .B(new_n576), .C1(new_n573), .C2(new_n281), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n594), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n578), .A2(new_n315), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n586), .A2(new_n593), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n596), .B2(new_n383), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n565), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n444), .A2(new_n557), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g0407(.A(new_n607), .B(KEYINPUT85), .Z(G372));
  NAND2_X1  g0408(.A1(new_n435), .A2(new_n430), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT18), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n363), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n306), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(new_n299), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n611), .B1(new_n614), .B2(new_n421), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n340), .B1(new_n615), .B2(new_n335), .ZN(new_n616));
  INV_X1    g0416(.A(new_n444), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n530), .A2(new_n339), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n618), .B(new_n560), .C1(new_n548), .C2(new_n554), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT87), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT87), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n565), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT86), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n601), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n595), .A2(new_n598), .A3(new_n600), .A4(KEYINPUT86), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n557), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n479), .A2(new_n487), .A3(new_n513), .A4(new_n503), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n630), .A2(KEYINPUT26), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n516), .A2(new_n517), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n479), .A2(new_n487), .A3(new_n503), .A4(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n479), .B1(new_n633), .B2(KEYINPUT26), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n616), .B1(new_n617), .B2(new_n636), .ZN(G369));
  NAND3_X1  g0437(.A1(new_n264), .A2(new_n227), .A3(G13), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT88), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT89), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n642));
  INV_X1    g0442(.A(G213), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n603), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n625), .A2(new_n626), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n601), .ZN(new_n650));
  INV_X1    g0450(.A(new_n605), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n649), .B1(new_n652), .B2(new_n648), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n555), .A2(new_n647), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n565), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n556), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n619), .B2(new_n647), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n620), .A2(new_n622), .A3(new_n647), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n601), .A2(new_n647), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n657), .A2(new_n663), .A3(new_n556), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n660), .A2(new_n661), .A3(new_n664), .ZN(G399));
  INV_X1    g0465(.A(new_n222), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n230), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n468), .A2(G116), .ZN(new_n669));
  INV_X1    g0469(.A(new_n667), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G1), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  INV_X1    g0473(.A(new_n647), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n633), .A2(KEYINPUT26), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n479), .B1(new_n630), .B2(KEYINPUT26), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n521), .B(new_n556), .C1(new_n565), .C2(new_n601), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT29), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n674), .B1(new_n629), .B2(new_n635), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(KEYINPUT29), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT91), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n596), .A2(G179), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n526), .A2(new_n281), .ZN(new_n685));
  INV_X1    g0485(.A(new_n522), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(new_n494), .A4(new_n500), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NOR4_X1   g0488(.A1(new_n684), .A2(new_n461), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n461), .A2(new_n687), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT30), .B1(new_n690), .B2(new_n599), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n596), .A2(new_n337), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n461), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n696), .A3(new_n461), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n527), .B1(new_n494), .B2(new_n500), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n647), .B1(new_n692), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n683), .B1(new_n700), .B2(KEYINPUT31), .ZN(new_n701));
  INV_X1    g0501(.A(new_n687), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n486), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n688), .B1(new_n703), .B2(new_n684), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n690), .A2(KEYINPUT30), .A3(new_n599), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n698), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n696), .B1(new_n693), .B2(new_n461), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n704), .B(new_n705), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n674), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(KEYINPUT91), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n606), .A2(new_n521), .A3(new_n556), .A4(new_n647), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n701), .A2(new_n711), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n682), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n673), .B1(new_n717), .B2(G1), .ZN(G364));
  AND2_X1   g0518(.A1(new_n227), .A2(G13), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n264), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n667), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n655), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n653), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT92), .Z(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n226), .B1(G20), .B2(new_n339), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n570), .A2(new_n666), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G355), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G116), .B2(new_n222), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n368), .A2(new_n666), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n445), .B2(new_n230), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n246), .A2(G45), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n227), .A2(G190), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n337), .A2(new_n383), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n227), .A2(new_n315), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n337), .A2(new_n383), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(G311), .A2(new_n741), .B1(new_n744), .B2(G322), .ZN(new_n745));
  INV_X1    g0545(.A(G326), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n227), .A2(new_n383), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n337), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n315), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n745), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G294), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n383), .A2(G179), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n742), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G303), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n570), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(new_n739), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n739), .A2(new_n752), .ZN(new_n764));
  INV_X1    g0564(.A(G329), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n762), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n751), .A2(new_n757), .A3(new_n761), .A4(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT94), .ZN(new_n768));
  INV_X1    g0568(.A(new_n748), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n768), .B1(new_n769), .B2(new_n315), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n748), .A2(KEYINPUT94), .A3(G190), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(G317), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n773), .A2(G68), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n755), .A2(new_n205), .ZN(new_n778));
  INV_X1    g0578(.A(new_n762), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(G107), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  OAI21_X1  g0581(.A(KEYINPUT32), .B1(new_n764), .B2(new_n781), .ZN(new_n782));
  OR3_X1    g0582(.A1(new_n764), .A2(KEYINPUT32), .A3(new_n781), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n276), .B1(new_n759), .B2(new_n213), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(KEYINPUT93), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n785), .A2(KEYINPUT93), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(new_n750), .C2(new_n256), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n397), .A2(new_n743), .B1(new_n740), .B2(new_n203), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n784), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n767), .A2(new_n776), .B1(new_n777), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n728), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n722), .B1(new_n730), .B2(new_n738), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT96), .ZN(new_n794));
  INV_X1    g0594(.A(new_n727), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n653), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n724), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  OR2_X1    g0598(.A1(new_n647), .A2(new_n359), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n612), .B1(new_n799), .B2(new_n360), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n674), .A2(new_n363), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n681), .B(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(new_n715), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n722), .B1(new_n803), .B2(new_n715), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n722), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n728), .A2(new_n725), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n203), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G137), .A2(new_n749), .B1(new_n741), .B2(G159), .ZN(new_n811));
  INV_X1    g0611(.A(G143), .ZN(new_n812));
  INV_X1    g0612(.A(G150), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(new_n812), .B2(new_n743), .C1(new_n772), .C2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT98), .Z(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT34), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n779), .A2(G68), .ZN(new_n818));
  INV_X1    g0618(.A(G132), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n256), .B2(new_n759), .C1(new_n819), .C2(new_n764), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n425), .B(new_n820), .C1(G58), .C2(new_n754), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n816), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G303), .A2(new_n749), .B1(new_n741), .B2(G116), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n772), .B2(new_n763), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT97), .Z(new_n825));
  NOR2_X1   g0625(.A1(new_n762), .A2(new_n213), .ZN(new_n826));
  INV_X1    g0626(.A(new_n764), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(G311), .B2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n828), .B(new_n570), .C1(new_n206), .C2(new_n759), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n778), .B(new_n829), .C1(G294), .C2(new_n744), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n792), .B1(new_n822), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n726), .ZN(new_n833));
  INV_X1    g0633(.A(new_n802), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n810), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n806), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  INV_X1    g0637(.A(new_n507), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n838), .A2(KEYINPUT35), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(KEYINPUT35), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n839), .A2(G116), .A3(new_n228), .A4(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT36), .Z(new_n842));
  OAI211_X1 g0642(.A(new_n230), .B(G77), .C1(new_n397), .C2(new_n211), .ZN(new_n843));
  INV_X1    g0643(.A(new_n201), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G68), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n264), .B(G13), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n719), .A2(new_n264), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n801), .B(KEYINPUT99), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n681), .B2(new_n802), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n674), .A2(new_n270), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n307), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n851), .B1(new_n299), .B2(new_n306), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT100), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n427), .A2(new_n253), .ZN(new_n858));
  INV_X1    g0658(.A(new_n402), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT16), .B1(new_n396), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n429), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n646), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n861), .A2(new_n646), .A3(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n861), .A2(new_n435), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n417), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT37), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT37), .B1(new_n385), .B2(new_n416), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n432), .A2(new_n433), .A3(new_n646), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n436), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n431), .B(new_n387), .C1(new_n405), .C2(new_n415), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT75), .B1(new_n428), .B2(new_n429), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n439), .B1(new_n876), .B2(new_n435), .ZN(new_n877));
  AND4_X1   g0677(.A1(new_n439), .A2(new_n432), .A3(new_n433), .A4(new_n435), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT76), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n421), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n866), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n873), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n443), .A2(new_n866), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n869), .B2(new_n872), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT102), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT102), .B(new_n887), .C1(new_n881), .C2(new_n882), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n885), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n887), .B1(new_n881), .B2(new_n882), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT102), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n889), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(KEYINPUT103), .A3(new_n885), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n857), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n610), .A2(new_n645), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT104), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n872), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n870), .A2(KEYINPUT104), .A3(new_n436), .A4(new_n871), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n871), .A2(new_n417), .A3(new_n609), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n871), .B1(new_n422), .B2(new_n611), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n884), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n894), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n891), .B2(KEYINPUT39), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n299), .A2(new_n674), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n900), .A2(new_n901), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n680), .B(new_n444), .C1(KEYINPUT29), .C2(new_n681), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n616), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n915), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n700), .B2(KEYINPUT31), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n709), .A2(KEYINPUT105), .A3(new_n710), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n713), .A2(new_n712), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n855), .A2(new_n834), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n897), .A2(KEYINPUT103), .A3(new_n885), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT103), .B1(new_n897), .B2(new_n885), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT40), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT106), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT106), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n909), .B2(new_n894), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n930), .A2(new_n931), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n924), .A2(new_n444), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  INV_X1    g0740(.A(G330), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n848), .B1(new_n918), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT107), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n943), .A2(new_n944), .B1(new_n918), .B2(new_n942), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n847), .B1(new_n945), .B2(new_n946), .ZN(G367));
  NOR2_X1   g0747(.A1(new_n242), .A2(new_n735), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n729), .B1(new_n222), .B2(new_n354), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n722), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n740), .A2(new_n763), .B1(new_n344), .B2(new_n755), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n773), .A2(G294), .B1(KEYINPUT110), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(G311), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n750), .A2(new_n953), .B1(new_n760), .B2(new_n743), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n827), .A2(G317), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n955), .B(new_n425), .C1(new_n205), .C2(new_n762), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n759), .A2(new_n588), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT46), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n954), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n952), .B(new_n959), .C1(KEYINPUT110), .C2(new_n951), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n773), .A2(G159), .B1(new_n201), .B2(new_n741), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT111), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n755), .A2(new_n211), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n827), .A2(G137), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n276), .B1(new_n759), .B2(new_n397), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n762), .A2(new_n203), .ZN(new_n967));
  NOR4_X1   g0767(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G143), .A2(new_n749), .B1(new_n744), .B2(G150), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n963), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n961), .A2(new_n962), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n960), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT47), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n950), .B1(new_n973), .B2(new_n728), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n647), .A2(new_n481), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(new_n479), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n479), .A3(new_n487), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n974), .B1(new_n795), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n980));
  INV_X1    g0780(.A(new_n978), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT43), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n632), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n514), .B(new_n520), .C1(new_n984), .C2(new_n647), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n674), .A2(new_n503), .A3(new_n632), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n664), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(KEYINPUT42), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT108), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n514), .B1(new_n988), .B2(new_n619), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n989), .A2(KEYINPUT42), .B1(new_n993), .B2(new_n647), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n980), .B(new_n983), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n660), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n992), .A2(new_n982), .A3(new_n981), .A4(new_n994), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n987), .A4(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n998), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n995), .A2(new_n1000), .B1(new_n660), .B2(new_n988), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n664), .A2(new_n661), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n988), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT44), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n664), .A2(new_n661), .A3(new_n987), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT45), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n1005), .A2(new_n1007), .A3(new_n997), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n997), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n664), .B1(new_n659), .B2(new_n663), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n654), .A2(KEYINPUT109), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n717), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n667), .B(KEYINPUT41), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n721), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n979), .B1(new_n1002), .B2(new_n1017), .ZN(G387));
  NAND2_X1  g0818(.A1(new_n717), .A2(new_n1013), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1014), .A2(new_n716), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n667), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1013), .A2(new_n721), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n238), .A2(new_n445), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1023), .A2(new_n734), .B1(new_n669), .B2(new_n731), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n352), .A2(new_n256), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n445), .B1(new_n211), .B2(new_n203), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1026), .A2(new_n669), .A3(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1024), .A2(new_n1028), .B1(G107), .B2(new_n222), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n807), .B1(new_n1029), .B2(new_n729), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n772), .A2(new_n321), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G50), .A2(new_n744), .B1(new_n741), .B2(G68), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n781), .B2(new_n750), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n759), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G77), .A2(new_n1034), .B1(new_n779), .B2(G97), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n827), .A2(G150), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n463), .A2(new_n754), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n368), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1031), .A2(new_n1033), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(G322), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n772), .A2(new_n953), .B1(new_n1040), .B2(new_n750), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT112), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT112), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G303), .A2(new_n741), .B1(new_n744), .B2(G317), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1034), .A2(G294), .B1(new_n754), .B2(G283), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT49), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n762), .A2(new_n588), .B1(new_n764), .B2(new_n746), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1052), .A2(new_n368), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1039), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1030), .B1(new_n659), .B2(new_n795), .C1(new_n1054), .C2(new_n792), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1022), .A2(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1021), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(G393));
  OAI21_X1  g0858(.A(new_n667), .B1(new_n1010), .B2(new_n1019), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1019), .B2(new_n1010), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n729), .B1(new_n205), .B2(new_n222), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n735), .A2(new_n250), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n722), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n773), .A2(new_n201), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n826), .B(new_n425), .C1(G77), .C2(new_n754), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n759), .A2(new_n211), .B1(new_n764), .B2(new_n812), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT113), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n741), .A2(new_n352), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1064), .A2(new_n1065), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G150), .A2(new_n749), .B1(new_n744), .B2(G159), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G317), .A2(new_n749), .B1(new_n744), .B2(G311), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n759), .A2(new_n763), .B1(new_n764), .B2(new_n1040), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n570), .B1(new_n762), .B2(new_n206), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(G116), .C2(new_n754), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n756), .B2(new_n740), .C1(new_n772), .C2(new_n760), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1070), .A2(new_n1072), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1063), .B1(new_n1079), .B2(new_n728), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n987), .B2(new_n795), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1010), .B2(new_n720), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1060), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(new_n913), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n912), .B1(new_n856), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n308), .A2(new_n851), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n854), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(KEYINPUT114), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n853), .B2(new_n854), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n849), .B1(new_n679), .B2(new_n802), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n913), .B(new_n910), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n855), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n714), .A2(new_n1096), .A3(G330), .A4(new_n802), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1086), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n941), .B1(new_n922), .B2(new_n923), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n444), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n916), .A2(new_n1100), .A3(new_n616), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n714), .A2(G330), .A3(new_n802), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n855), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(new_n925), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n850), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n941), .B(new_n834), .C1(new_n922), .C2(new_n923), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1094), .B(new_n1097), .C1(new_n1108), .C2(new_n1092), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1101), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1098), .B(new_n1110), .C1(new_n1111), .C2(new_n1104), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1110), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1086), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1104), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1112), .A2(new_n1116), .A3(new_n667), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n570), .B1(new_n827), .B2(G125), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n781), .B2(new_n755), .C1(new_n844), .C2(new_n762), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  NAND3_X1  g0920(.A1(new_n1034), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n759), .B2(new_n813), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n741), .A2(new_n1120), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1124), .B1(new_n819), .B2(new_n743), .C1(new_n1125), .C2(new_n750), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1119), .B(new_n1126), .C1(G137), .C2(new_n773), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G68), .A2(new_n779), .B1(new_n827), .B2(G294), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT115), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n570), .B1(new_n759), .B2(new_n213), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1128), .B1(new_n203), .B2(new_n755), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n741), .A2(G97), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n588), .B2(new_n743), .C1(new_n763), .C2(new_n750), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(new_n343), .C2(new_n773), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n728), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n807), .B1(new_n321), .B2(new_n808), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n912), .B2(new_n833), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n721), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1117), .A2(new_n1140), .ZN(G378));
  INV_X1    g0941(.A(G41), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n425), .A2(new_n1142), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n206), .A2(new_n743), .B1(new_n740), .B2(new_n354), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G116), .C2(new_n749), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n779), .A2(G58), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n203), .B2(new_n759), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n964), .B(new_n1147), .C1(G283), .C2(new_n827), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1145), .B(new_n1148), .C1(new_n205), .C2(new_n772), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT58), .ZN(new_n1150));
  AOI21_X1  g0950(.A(G50), .B1(new_n273), .B2(new_n1142), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1149), .A2(new_n1150), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n749), .A2(G125), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n744), .A2(G128), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1034), .A2(new_n1120), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n754), .A2(G150), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n773), .A2(G132), .B1(G137), .B2(new_n741), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(KEYINPUT116), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(KEYINPUT116), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1157), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT59), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n273), .B(new_n1142), .C1(new_n762), .C2(new_n781), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G124), .B2(new_n827), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1152), .B1(new_n1150), .B2(new_n1149), .C1(new_n1165), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n728), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n807), .B1(new_n844), .B2(new_n808), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n335), .A2(new_n341), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n326), .A2(new_n645), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1170), .B(new_n1171), .C1(new_n1178), .C2(new_n726), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT119), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n941), .B1(new_n936), .B2(new_n933), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n926), .B1(new_n893), .B2(new_n898), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1182), .B2(KEYINPUT40), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT120), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(KEYINPUT120), .B(new_n1181), .C1(new_n1182), .C2(KEYINPUT40), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n1186), .A3(new_n1178), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1183), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1178), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(KEYINPUT120), .A3(new_n1189), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1187), .A2(new_n915), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n915), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1180), .B1(new_n1193), .B2(new_n721), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1101), .B1(new_n1139), .B2(new_n1110), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT57), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n915), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1187), .A2(new_n915), .A3(new_n1190), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n916), .A2(new_n1100), .A3(new_n616), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(new_n1112), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1200), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n667), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1194), .B1(new_n1197), .B2(new_n1206), .ZN(G375));
  NAND3_X1  g1007(.A1(new_n1107), .A2(new_n1109), .A3(new_n1101), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1113), .A2(new_n1208), .A3(new_n1016), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1102), .A2(new_n855), .B1(new_n1099), .B2(new_n925), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1097), .A2(new_n1094), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1092), .B1(new_n1099), .B2(new_n802), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1210), .A2(new_n850), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n721), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n807), .B1(new_n211), .B2(new_n808), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n759), .A2(new_n205), .B1(new_n764), .B2(new_n760), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1216), .A2(new_n276), .A3(new_n967), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1037), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n750), .A2(new_n756), .B1(new_n344), .B2(new_n740), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G283), .C2(new_n744), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n773), .A2(G116), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G137), .A2(new_n744), .B1(new_n741), .B2(G150), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n819), .B2(new_n750), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1146), .B1(new_n1125), .B2(new_n764), .C1(new_n781), .C2(new_n759), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n368), .B1(new_n755), .B2(new_n256), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n773), .A2(new_n1120), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1220), .A2(new_n1221), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n725), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1215), .B1(new_n792), .B2(new_n1228), .C1(new_n1092), .C2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1214), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1209), .A2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT121), .ZN(G381));
  NOR2_X1   g1034(.A1(G393), .A2(G396), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n836), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT122), .Z(new_n1237));
  NOR4_X1   g1037(.A1(new_n1237), .A2(G387), .A3(G390), .A4(G381), .ZN(new_n1238));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1200), .A2(new_n721), .A3(new_n1201), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1180), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n670), .B1(new_n1193), .B2(new_n1204), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1200), .A2(new_n1196), .A3(new_n1201), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1202), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1242), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1238), .A2(new_n1239), .A3(new_n1246), .ZN(G407));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1239), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G407), .B(G213), .C1(G343), .C2(new_n1248), .ZN(G409));
  INV_X1    g1049(.A(KEYINPUT123), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT60), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1213), .B2(new_n1203), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1213), .A2(new_n1203), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n667), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n1101), .A4(new_n1109), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1250), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1208), .B1(new_n1110), .B2(new_n1251), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1258), .A2(KEYINPUT123), .A3(new_n667), .A4(new_n1255), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1260), .B2(new_n1232), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n836), .B(new_n1231), .C1(new_n1257), .C2(new_n1259), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n643), .A2(G343), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1117), .A2(new_n1140), .A3(new_n1179), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1193), .B2(new_n721), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1193), .A2(new_n1016), .A3(new_n1196), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1264), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1263), .B(new_n1268), .C1(new_n1246), .C2(new_n1239), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT62), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G375), .A2(G378), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1263), .A4(new_n1268), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1264), .A2(G2897), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1264), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(KEYINPUT124), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1275), .B1(new_n1263), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1275), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(new_n1261), .A2(new_n1262), .A3(new_n1280), .A4(new_n1277), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1191), .A2(new_n1192), .A3(new_n1195), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n667), .B(new_n1205), .C1(new_n1283), .C2(KEYINPUT57), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1239), .B1(new_n1284), .B2(new_n1194), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1276), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1282), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1270), .A2(new_n1273), .A3(new_n1274), .A4(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1057), .A2(new_n797), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1235), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(KEYINPUT125), .B(new_n979), .C1(new_n1002), .C2(new_n1017), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  AND3_X1   g1093(.A1(G390), .A2(G387), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G390), .B1(G387), .B2(new_n1293), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1291), .B(new_n1292), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1083), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(G390), .A2(G387), .A3(new_n1297), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1299), .B(new_n1300), .C1(new_n1235), .C2(new_n1290), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1289), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1302), .B1(new_n1269), .B2(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1271), .A2(KEYINPUT63), .A3(new_n1263), .A4(new_n1268), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1305), .A2(new_n1274), .A3(new_n1306), .A4(new_n1288), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1303), .A2(new_n1307), .ZN(G405));
  INV_X1    g1108(.A(KEYINPUT127), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1263), .A2(new_n1309), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1302), .B(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1271), .A2(new_n1248), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1311), .B(new_n1312), .ZN(G402));
endmodule


