//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT3), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n192), .B2(G104), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n190), .A2(KEYINPUT82), .A3(G107), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(new_n195), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n190), .A2(G107), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n192), .A2(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(G101), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT2), .B(G113), .ZN(new_n205));
  OR2_X1    g019(.A1(KEYINPUT66), .A2(G116), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT66), .A2(G116), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(G119), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(G116), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n206), .A2(new_n209), .A3(G119), .A4(new_n207), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT89), .B(KEYINPUT5), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(G116), .ZN(new_n218));
  OAI21_X1  g032(.A(G113), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n212), .A2(new_n213), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(new_n217), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n192), .A2(KEYINPUT3), .A3(G104), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(new_n192), .B2(G104), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n197), .B(new_n198), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n229), .A3(G101), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n212), .A2(new_n205), .A3(new_n213), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(new_n214), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n223), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n212), .A2(new_n205), .A3(new_n213), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n215), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n236), .A2(KEYINPUT88), .A3(new_n230), .A4(new_n228), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n222), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n188), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n238), .B2(KEYINPUT90), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT90), .ZN(new_n243));
  AOI211_X1 g057(.A(new_n243), .B(new_n222), .C1(new_n234), .C2(new_n237), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n240), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n234), .A2(new_n237), .ZN(new_n246));
  INV_X1    g060(.A(new_n222), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n243), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n238), .A2(KEYINPUT90), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n249), .A2(new_n188), .A3(new_n250), .A4(new_n241), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G143), .B(G146), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n263), .A2(KEYINPUT91), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(KEYINPUT91), .ZN(new_n265));
  INV_X1    g079(.A(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n267));
  OAI22_X1  g081(.A1(new_n267), .A2(new_n253), .B1(new_n255), .B2(G128), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT65), .B1(new_n261), .B2(new_n267), .ZN(new_n270));
  AND4_X1   g084(.A1(KEYINPUT65), .A2(new_n267), .A3(new_n253), .A4(new_n255), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n264), .B(new_n265), .C1(G125), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G224), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G953), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n273), .B(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n245), .A2(new_n251), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G210), .B1(G237), .B2(G902), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n239), .B(KEYINPUT8), .Z(new_n279));
  AND2_X1   g093(.A1(new_n220), .A2(KEYINPUT5), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n215), .B(new_n204), .C1(new_n280), .C2(new_n219), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n203), .B1(new_n221), .B2(new_n214), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT7), .B1(new_n274), .B2(G953), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n273), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n263), .B1(new_n272), .B2(G125), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n283), .B(new_n285), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n238), .A2(new_n239), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n277), .A2(new_n278), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n278), .B1(new_n277), .B2(new_n289), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n187), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT92), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G953), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n295), .A2(G952), .ZN(new_n296));
  NAND2_X1  g110(.A1(G234), .A2(G237), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT21), .B(G898), .Z(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(G902), .A3(G953), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  INV_X1    g116(.A(G237), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n303), .A2(new_n295), .A3(G214), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT93), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(G143), .ZN(new_n306));
  INV_X1    g120(.A(G131), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT93), .B(G143), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n306), .B(new_n307), .C1(new_n304), .C2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n304), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n303), .A2(new_n295), .A3(G214), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(KEYINPUT93), .B2(new_n252), .ZN(new_n312));
  OAI21_X1  g126(.A(G131), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT17), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n309), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G125), .B(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT16), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n254), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n317), .A2(G146), .A3(new_n320), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT17), .B(G131), .C1(new_n310), .C2(new_n312), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n315), .A2(new_n322), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G113), .B(G122), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(new_n190), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT80), .B1(new_n330), .B2(G146), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n316), .A2(new_n332), .A3(new_n254), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n254), .B2(new_n316), .ZN(new_n335));
  NAND2_X1  g149(.A1(KEYINPUT94), .A2(KEYINPUT18), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(G131), .B(new_n337), .C1(new_n310), .C2(new_n312), .ZN(new_n338));
  OAI221_X1 g152(.A(new_n306), .B1(new_n307), .B2(new_n336), .C1(new_n304), .C2(new_n308), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n325), .A2(new_n327), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n327), .B1(new_n325), .B2(new_n340), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n302), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G475), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT20), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n309), .A2(new_n313), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n323), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n316), .B(KEYINPUT19), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n254), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n317), .A2(KEYINPUT79), .A3(new_n320), .A4(G146), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n347), .A2(new_n349), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n340), .ZN(new_n354));
  INV_X1    g168(.A(new_n327), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n341), .ZN(new_n357));
  NOR2_X1   g171(.A1(G475), .A2(G902), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n346), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n358), .ZN(new_n360));
  AOI211_X1 g174(.A(KEYINPUT20), .B(new_n360), .C1(new_n356), .C2(new_n341), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n345), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT95), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT95), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n345), .B(new_n364), .C1(new_n359), .C2(new_n361), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT13), .B1(new_n266), .B2(G143), .ZN(new_n366));
  INV_X1    g180(.A(G134), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G128), .B(G143), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n206), .A2(new_n207), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G122), .ZN(new_n372));
  INV_X1    g186(.A(G122), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G116), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n192), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n192), .B1(new_n372), .B2(new_n374), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n370), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT9), .B(G234), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(G217), .A3(new_n295), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n371), .A2(KEYINPUT14), .A3(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G107), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n372), .A2(new_n374), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT96), .B(G134), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n369), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n375), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n378), .B(new_n382), .C1(new_n388), .C2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT97), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n385), .A2(KEYINPUT14), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n375), .B(new_n390), .C1(new_n395), .C2(new_n384), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n378), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n381), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n396), .A2(KEYINPUT97), .A3(new_n378), .A4(new_n382), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT15), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G478), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n400), .A2(new_n302), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n400), .B2(new_n302), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AND4_X1   g219(.A1(new_n301), .A2(new_n363), .A3(new_n365), .A4(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT92), .B(new_n187), .C1(new_n290), .C2(new_n291), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n294), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G234), .ZN(new_n409));
  OAI21_X1  g223(.A(G217), .B1(new_n409), .B2(G902), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT74), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT23), .B1(new_n266), .B2(G119), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT76), .B1(new_n210), .B2(G128), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n412), .B(new_n413), .Z(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G110), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT77), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n322), .A2(new_n323), .ZN(new_n418));
  XOR2_X1   g232(.A(G119), .B(G128), .Z(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT75), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT24), .B(G110), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n417), .B(new_n418), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n349), .A2(new_n352), .A3(new_n334), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(KEYINPUT78), .A3(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(G110), .B2(new_n414), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT78), .B1(new_n420), .B2(new_n421), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT22), .B(G137), .ZN(new_n429));
  INV_X1    g243(.A(G221), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n430), .A2(new_n409), .A3(G953), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n429), .B(new_n431), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n422), .A2(new_n427), .A3(new_n432), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT25), .ZN(new_n436));
  AOI21_X1  g250(.A(G902), .B1(new_n436), .B2(KEYINPUT81), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n411), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n439), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n434), .A2(new_n441), .A3(new_n435), .A4(new_n437), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n434), .A2(new_n435), .ZN(new_n444));
  AOI21_X1  g258(.A(G902), .B1(new_n409), .B2(G217), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT72), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n450));
  INV_X1    g264(.A(G137), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(G134), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT64), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n367), .B2(G137), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n454), .B2(KEYINPUT11), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT64), .B1(new_n451), .B2(G134), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT11), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n307), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n367), .A2(G137), .ZN(new_n460));
  OAI21_X1  g274(.A(G131), .B1(new_n460), .B2(new_n452), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n267), .A2(new_n253), .A3(new_n255), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT65), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n261), .A2(KEYINPUT65), .A3(new_n267), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n268), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n450), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n272), .A2(KEYINPUT69), .A3(new_n461), .A4(new_n459), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT68), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n257), .B(new_n470), .C1(new_n260), .C2(new_n261), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n455), .A2(new_n307), .A3(new_n458), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n307), .B1(new_n455), .B2(new_n458), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n471), .B(new_n472), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n468), .A2(new_n469), .A3(new_n475), .A4(new_n233), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT70), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n468), .A2(new_n469), .A3(new_n475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT30), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n455), .A2(new_n458), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G131), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n459), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n254), .A2(G143), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n252), .A2(G146), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n259), .B(new_n258), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n257), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n272), .A2(new_n461), .A3(new_n459), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n233), .B1(new_n480), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT26), .B(G101), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n303), .A2(new_n295), .A3(G210), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n478), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n449), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n480), .A2(new_n490), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n236), .ZN(new_n501));
  INV_X1    g315(.A(new_n496), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n462), .A2(new_n467), .ZN(new_n503));
  INV_X1    g317(.A(new_n471), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n470), .B1(new_n486), .B2(new_n257), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n503), .A2(KEYINPUT69), .B1(new_n506), .B2(new_n483), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n507), .A2(new_n477), .A3(new_n233), .A4(new_n468), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n476), .A2(KEYINPUT70), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n501), .A2(new_n502), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT28), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n233), .A2(new_n489), .ZN(new_n514));
  INV_X1    g328(.A(new_n475), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n233), .B1(new_n487), .B2(new_n489), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n508), .B2(new_n509), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n518), .B2(new_n513), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n496), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n497), .A2(new_n498), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n499), .A2(new_n512), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT32), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT73), .B1(new_n519), .B2(new_n496), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT28), .B1(new_n478), .B2(new_n517), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT73), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n502), .A4(new_n516), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n500), .A2(new_n236), .B1(new_n508), .B2(new_n509), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n496), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n529), .A2(new_n532), .A3(new_n533), .A4(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n516), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n479), .A2(new_n236), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n510), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n538), .B1(new_n540), .B2(KEYINPUT28), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n496), .A2(new_n533), .ZN(new_n542));
  AOI21_X1  g356(.A(G902), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G472), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n448), .B1(new_n528), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n430), .B1(new_n380), .B2(new_n302), .ZN(new_n547));
  INV_X1    g361(.A(G469), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(new_n302), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n203), .B2(new_n467), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n272), .A2(KEYINPUT83), .A3(new_n199), .A4(new_n202), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n203), .A2(new_n467), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n554), .A2(KEYINPUT12), .A3(new_n483), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT12), .B1(new_n554), .B2(new_n483), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT86), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n483), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(KEYINPUT12), .A3(new_n483), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n204), .A2(KEYINPUT10), .A3(new_n272), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n472), .A2(new_n471), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n231), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n551), .A2(new_n552), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT84), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT84), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n551), .A2(new_n552), .A3(new_n571), .A4(new_n568), .ZN(new_n572));
  AOI211_X1 g386(.A(new_n483), .B(new_n567), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G140), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n295), .A2(G227), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n574), .B(new_n575), .Z(new_n576));
  OAI21_X1  g390(.A(KEYINPUT87), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n570), .A2(new_n572), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n473), .A2(new_n474), .ZN(new_n579));
  INV_X1    g393(.A(new_n567), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT87), .ZN(new_n582));
  INV_X1    g396(.A(new_n576), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n564), .A2(new_n577), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n567), .B1(new_n570), .B2(new_n572), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(new_n579), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n576), .B1(new_n587), .B2(new_n573), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n549), .B1(new_n589), .B2(new_n548), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT85), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n555), .A2(new_n556), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n573), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n560), .A2(new_n562), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n581), .A2(KEYINPUT85), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n576), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n587), .A2(new_n573), .A3(new_n576), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(G469), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n547), .B1(new_n590), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n408), .A2(new_n546), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND2_X1  g417(.A1(new_n522), .A2(new_n302), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n604), .A2(G472), .B1(new_n523), .B2(new_n522), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n585), .A2(new_n588), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n548), .A3(new_n302), .ZN(new_n607));
  INV_X1    g421(.A(new_n549), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n600), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n547), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n605), .A2(new_n447), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n187), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n277), .A2(new_n289), .ZN(new_n613));
  INV_X1    g427(.A(new_n278), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n277), .A2(new_n278), .A3(new_n289), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n396), .A2(new_n378), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n381), .A2(KEYINPUT98), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n397), .A2(KEYINPUT98), .A3(new_n381), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n400), .A2(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G478), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n400), .A2(new_n302), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n624), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n365), .B2(new_n363), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n617), .A2(new_n301), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n611), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND2_X1  g448(.A1(new_n615), .A2(new_n616), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n301), .A3(new_n187), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n359), .B2(new_n361), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n327), .B1(new_n353), .B2(new_n340), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n358), .B1(new_n342), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT20), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n357), .A2(new_n346), .A3(new_n358), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(KEYINPUT99), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n405), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n345), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n611), .A2(new_n636), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT100), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT35), .B(G107), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n433), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT101), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n428), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n445), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n443), .A2(new_n657), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n449), .B(new_n498), .C1(new_n534), .C2(new_n502), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT72), .B1(new_n511), .B2(KEYINPUT31), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n496), .A2(new_n519), .B1(new_n497), .B2(new_n498), .ZN(new_n662));
  AOI21_X1  g476(.A(G902), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(G472), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n524), .B(new_n658), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT102), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n604), .A2(G472), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n667), .A2(new_n668), .A3(new_n524), .A4(new_n658), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n601), .A2(new_n406), .A3(new_n294), .A4(new_n407), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT37), .B(G110), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  AND3_X1   g488(.A1(new_n609), .A2(new_n617), .A3(new_n610), .ZN(new_n675));
  INV_X1    g489(.A(new_n527), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n526), .B1(new_n522), .B2(new_n523), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n545), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n298), .B1(G900), .B2(new_n300), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n638), .A2(new_n643), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n647), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n675), .A2(new_n678), .A3(new_n658), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NAND2_X1  g497(.A1(new_n609), .A2(new_n610), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n679), .B(KEYINPUT39), .Z(new_n685));
  OR2_X1    g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n535), .A2(new_n502), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n689), .B(new_n302), .C1(new_n502), .C2(new_n540), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G472), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n528), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n290), .A2(new_n291), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT38), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT38), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n635), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n363), .A2(new_n365), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n646), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n697), .A2(new_n612), .A3(new_n658), .A4(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n687), .A2(new_n688), .A3(new_n692), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  NAND2_X1  g516(.A1(new_n626), .A2(new_n628), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n698), .A2(new_n703), .A3(new_n679), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n675), .A2(new_n678), .A3(new_n658), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  INV_X1    g520(.A(new_n636), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n678), .A3(new_n447), .A4(new_n630), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n586), .A2(new_n579), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n583), .B1(new_n709), .B2(new_n581), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n582), .B1(new_n581), .B2(new_n583), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n557), .A2(new_n563), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n710), .B1(new_n713), .B2(new_n584), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n714), .B2(G902), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n610), .A3(new_n607), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT103), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n715), .A2(new_n718), .A3(new_n610), .A4(new_n607), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n708), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT41), .B(G113), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  NAND3_X1  g537(.A1(new_n717), .A2(new_n707), .A3(new_n719), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n678), .A2(new_n447), .A3(new_n648), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n726), .B1(new_n724), .B2(new_n725), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  NOR2_X1   g545(.A1(new_n589), .A2(new_n548), .ZN(new_n732));
  AOI211_X1 g546(.A(G469), .B(G902), .C1(new_n585), .C2(new_n588), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n610), .A2(new_n734), .A3(new_n406), .A4(new_n617), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n525), .A2(new_n527), .B1(G472), .B2(new_n544), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n440), .A2(new_n442), .B1(new_n445), .B2(new_n656), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  AND3_X1   g554(.A1(new_n717), .A2(new_n707), .A3(new_n719), .ZN(new_n741));
  INV_X1    g555(.A(new_n699), .ZN(new_n742));
  INV_X1    g556(.A(new_n523), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n511), .B(new_n498), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n541), .A2(new_n502), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n667), .A2(new_n447), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n667), .A2(new_n447), .A3(KEYINPUT105), .A4(new_n747), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n741), .A2(new_n742), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT106), .B(G122), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G24));
  NAND3_X1  g569(.A1(new_n734), .A2(new_n610), .A3(new_n617), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n667), .A2(new_n704), .A3(new_n747), .A4(new_n658), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n328), .ZN(G27));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n600), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n598), .B1(new_n596), .B2(new_n576), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT107), .A3(G469), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n590), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n610), .A2(new_n187), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n635), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n678), .A2(new_n765), .A3(new_n447), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n704), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n760), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n765), .A2(new_n767), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n546), .A3(KEYINPUT42), .A4(new_n704), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  XNOR2_X1  g588(.A(new_n681), .B(KEYINPUT108), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n367), .ZN(G36));
  OAI21_X1  g591(.A(G469), .B1(new_n763), .B2(KEYINPUT45), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT109), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n780), .B(G469), .C1(new_n763), .C2(KEYINPUT45), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n763), .A2(KEYINPUT45), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n608), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n607), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n778), .A2(KEYINPUT109), .B1(KEYINPUT45), .B2(new_n763), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n549), .B1(new_n786), .B2(new_n781), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n610), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(new_n685), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n605), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n703), .A2(new_n363), .A3(new_n365), .ZN(new_n793));
  XNOR2_X1  g607(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n795), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(new_n658), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n615), .A2(new_n187), .A3(new_n616), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n798), .B2(new_n799), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n791), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NOR2_X1   g618(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n805));
  NAND2_X1  g619(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n789), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n610), .B(new_n806), .C1(new_n785), .C2(new_n788), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n678), .A2(new_n447), .A3(new_n769), .A4(new_n801), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NOR2_X1   g626(.A1(G952), .A2(G953), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT120), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n678), .A2(new_n447), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n698), .A2(new_n629), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n363), .A2(new_n405), .A3(new_n365), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n818), .A2(new_n301), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n294), .A2(new_n820), .A3(new_n407), .ZN(new_n821));
  OAI22_X1  g635(.A1(new_n671), .A2(new_n817), .B1(new_n821), .B2(new_n611), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n816), .B1(new_n822), .B2(new_n672), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n408), .A2(new_n601), .A3(new_n666), .A4(new_n669), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n294), .A2(new_n820), .A3(new_n407), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n667), .A2(new_n524), .A3(new_n447), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n684), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(new_n602), .A3(KEYINPUT113), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n716), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n406), .A3(new_n617), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n678), .A2(new_n658), .ZN(new_n833));
  OAI22_X1  g647(.A1(new_n708), .A2(new_n720), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n724), .A2(new_n699), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(new_n752), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n345), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n403), .A3(new_n404), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n644), .A2(new_n838), .A3(new_n839), .A4(new_n679), .ZN(new_n840));
  INV_X1    g654(.A(new_n404), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n400), .A2(new_n302), .A3(new_n402), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n345), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT114), .B1(new_n680), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n801), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n678), .A2(new_n846), .A3(new_n601), .A4(new_n658), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n664), .B1(new_n522), .B2(new_n302), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n746), .A3(new_n737), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n765), .A3(new_n767), .A4(new_n704), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n847), .B(new_n850), .C1(new_n768), .C2(new_n775), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n770), .B2(new_n772), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n830), .A2(new_n730), .A3(new_n836), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n758), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n682), .A3(new_n705), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n737), .A2(new_n610), .A3(new_n679), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n765), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n693), .A2(new_n612), .A3(new_n699), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n692), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n857), .B1(new_n765), .B2(new_n856), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT52), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n678), .A2(new_n601), .A3(new_n617), .A4(new_n658), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n758), .B1(new_n864), .B2(new_n681), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  INV_X1    g680(.A(new_n861), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n692), .A3(new_n858), .A4(new_n859), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n865), .A2(new_n866), .A3(new_n868), .A4(new_n705), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n815), .B1(new_n853), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n863), .A2(new_n869), .ZN(new_n872));
  INV_X1    g686(.A(new_n720), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n736), .A2(new_n631), .A3(new_n448), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n873), .A2(new_n874), .B1(new_n735), .B2(new_n738), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n736), .A2(new_n448), .A3(new_n649), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT104), .B1(new_n741), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n875), .B(new_n753), .C1(new_n877), .C2(new_n727), .ZN(new_n878));
  INV_X1    g692(.A(new_n851), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n773), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n865), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n815), .B1(new_n882), .B2(KEYINPUT52), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n872), .A2(new_n881), .A3(new_n830), .A4(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n885));
  AND3_X1   g699(.A1(new_n871), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n815), .B1(new_n865), .B2(new_n866), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n872), .A2(new_n881), .A3(new_n830), .A4(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n887), .B1(new_n871), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n298), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n767), .A2(new_n797), .A3(new_n734), .A4(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT118), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT48), .B1(new_n894), .B2(new_n817), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n893), .B(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT48), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n546), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n797), .A2(new_n892), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n750), .B2(new_n751), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n617), .A3(new_n831), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n295), .A2(G952), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n528), .A2(new_n691), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n715), .A2(new_n607), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(new_n298), .ZN(new_n907));
  AND4_X1   g721(.A1(new_n447), .A2(new_n905), .A3(new_n907), .A4(new_n767), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n908), .B2(new_n630), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n900), .A2(new_n903), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n698), .A2(new_n703), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n897), .A2(new_n849), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n697), .A2(new_n831), .A3(new_n612), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n902), .A2(new_n914), .B1(KEYINPUT117), .B2(KEYINPUT50), .ZN(new_n915));
  NOR2_X1   g729(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI211_X1 g731(.A(KEYINPUT117), .B(KEYINPUT50), .C1(new_n902), .C2(new_n914), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n733), .B1(new_n787), .B2(KEYINPUT46), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n547), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n807), .A2(new_n805), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n809), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n906), .A2(new_n610), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n801), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n902), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n919), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n911), .B1(new_n931), .B2(KEYINPUT51), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n913), .B(KEYINPUT51), .C1(new_n917), .C2(new_n918), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n925), .B1(new_n808), .B2(new_n809), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n934), .B2(KEYINPUT119), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n933), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n814), .B1(new_n891), .B2(new_n939), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n448), .A2(new_n766), .A3(new_n793), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT112), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n942), .A2(new_n697), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n734), .B(KEYINPUT49), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n905), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT121), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n907), .A2(new_n767), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(new_n447), .A3(new_n905), .A4(new_n912), .ZN(new_n950));
  INV_X1    g764(.A(new_n849), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n894), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n916), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n902), .A2(new_n914), .ZN(new_n954));
  AND2_X1   g768(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n915), .A2(new_n916), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n934), .B2(new_n929), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT51), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n910), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n933), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n930), .B1(new_n927), .B2(new_n936), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n934), .A2(KEYINPUT119), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n966), .A2(new_n886), .A3(new_n890), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n948), .B(new_n945), .C1(new_n967), .C2(new_n814), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n947), .A2(new_n968), .ZN(G75));
  NOR2_X1   g783(.A1(new_n295), .A2(G952), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n302), .B1(new_n871), .B2(new_n884), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT56), .B1(new_n972), .B2(G210), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n245), .A2(new_n251), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(new_n276), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT55), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n971), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n973), .B2(new_n977), .ZN(G51));
  NAND3_X1  g793(.A1(new_n972), .A2(new_n781), .A3(new_n786), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT123), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n871), .A2(new_n884), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(new_n885), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n549), .B(KEYINPUT122), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT57), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n606), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n970), .B1(new_n981), .B2(new_n986), .ZN(G54));
  NAND2_X1  g801(.A1(KEYINPUT58), .A2(G475), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT124), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n972), .A2(new_n357), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n357), .B1(new_n972), .B2(new_n989), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n990), .A2(new_n991), .A3(new_n970), .ZN(G60));
  INV_X1    g806(.A(new_n891), .ZN(new_n993));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT59), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n623), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n623), .A2(new_n995), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n971), .B1(new_n983), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(G63));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT60), .Z(new_n1001));
  NAND3_X1  g815(.A1(new_n982), .A2(new_n656), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n982), .A2(new_n1001), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n971), .B(new_n1002), .C1(new_n1003), .C2(new_n444), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT61), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(G66));
  AOI21_X1  g820(.A(new_n295), .B1(new_n299), .B2(G224), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n830), .A2(new_n730), .A3(new_n836), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n295), .ZN(new_n1009));
  INV_X1    g823(.A(G898), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n974), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1009), .B(new_n1011), .ZN(G69));
  NAND2_X1  g826(.A1(G900), .A2(G953), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n791), .A2(new_n546), .A3(new_n859), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n776), .B(new_n855), .C1(new_n770), .C2(new_n772), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n803), .A2(new_n1014), .A3(new_n811), .A4(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1013), .B1(new_n1016), .B2(G953), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n500), .B(KEYINPUT125), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(new_n350), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n701), .A2(new_n705), .A3(new_n865), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT62), .Z(new_n1021));
  NAND2_X1  g835(.A1(new_n818), .A2(new_n819), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT126), .ZN(new_n1023));
  OR4_X1    g837(.A1(new_n817), .A2(new_n686), .A3(new_n1023), .A4(new_n801), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1021), .A2(new_n803), .A3(new_n811), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1019), .A2(G953), .ZN(new_n1026));
  AOI22_X1  g840(.A1(new_n1017), .A2(new_n1019), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n295), .B1(G227), .B2(G900), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(G72));
  NAND2_X1  g843(.A1(G472), .A2(G902), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT63), .Z(new_n1031));
  OAI21_X1  g845(.A(new_n1031), .B1(new_n1025), .B2(new_n1008), .ZN(new_n1032));
  INV_X1    g846(.A(new_n689), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1031), .B1(new_n1016), .B2(new_n1008), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1035), .A2(new_n496), .A3(new_n534), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n871), .A2(new_n889), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n511), .A2(KEYINPUT127), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n536), .B(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1037), .A2(new_n1031), .A3(new_n1039), .ZN(new_n1040));
  AND4_X1   g854(.A1(new_n971), .A2(new_n1034), .A3(new_n1036), .A4(new_n1040), .ZN(G57));
endmodule


