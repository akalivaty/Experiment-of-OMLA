//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n210));
  NAND4_X1  g0010(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n212), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  NOR4_X1   g0024(.A1(new_n215), .A2(new_n217), .A3(new_n221), .A4(new_n224), .ZN(G361));
  XOR2_X1   g0025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT67), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT68), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT69), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n231), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G68), .ZN(new_n242));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n240), .B(new_n247), .ZN(G351));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n219), .A2(G33), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT15), .B(G87), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(KEYINPUT70), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n220), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n262), .A2(new_n219), .A3(G1), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n255), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n260), .A2(new_n263), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(G77), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(G274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n279), .A2(G244), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G232), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(G238), .A3(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G107), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n281), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n287));
  AOI211_X1 g0087(.A(new_n276), .B(new_n280), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n269), .B1(new_n288), .B2(G190), .ZN(new_n289));
  INV_X1    g0089(.A(G200), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n288), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n293), .B(new_n269), .C1(G169), .C2(new_n288), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g0095(.A(new_n295), .B(KEYINPUT71), .Z(new_n296));
  INV_X1    g0096(.A(G226), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n275), .B1(new_n278), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n281), .A2(G223), .A3(G1698), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n281), .A2(new_n282), .ZN(new_n300));
  INV_X1    g0100(.A(G222), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n299), .B1(new_n261), .B2(new_n281), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n298), .B1(new_n302), .B2(new_n287), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n265), .A2(G50), .A3(new_n267), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n251), .A2(G150), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n249), .B2(new_n253), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n219), .B1(new_n201), .B2(new_n241), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n260), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n263), .A2(new_n241), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n305), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n304), .A2(G200), .B1(new_n311), .B2(KEYINPUT9), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n305), .A2(new_n309), .A3(new_n310), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n303), .A2(G190), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT10), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n312), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n304), .A2(G179), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n313), .B1(new_n303), .B2(G169), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n296), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n243), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n261), .B2(new_n253), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n328), .A2(new_n260), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(KEYINPUT11), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n262), .A2(G1), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G20), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(G68), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT12), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n329), .A2(KEYINPUT11), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n265), .A2(G68), .A3(new_n267), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n330), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT72), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n281), .A2(G232), .A3(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G97), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(new_n300), .C2(new_n297), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n287), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n276), .B1(G238), .B2(new_n279), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT13), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT13), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n346), .A3(new_n343), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(G169), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n292), .B2(new_n348), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n349), .B1(new_n348), .B2(G169), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n338), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n290), .B1(new_n345), .B2(new_n347), .ZN(new_n354));
  INV_X1    g0154(.A(G190), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  OR3_X1    g0156(.A1(new_n338), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G33), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT3), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT3), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G33), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n359), .A2(new_n361), .A3(G226), .A4(G1698), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n359), .A2(new_n361), .A3(G223), .A4(new_n282), .ZN(new_n363));
  INV_X1    g0163(.A(G87), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(new_n363), .C1(new_n358), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n287), .ZN(new_n366));
  INV_X1    g0166(.A(G232), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n275), .B1(new_n367), .B2(new_n278), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(new_n355), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n287), .B2(new_n365), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(G200), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n249), .B1(new_n266), .B2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n265), .A2(new_n373), .B1(new_n263), .B2(new_n249), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n281), .B2(G20), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n360), .A2(G33), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n358), .A2(KEYINPUT3), .ZN(new_n378));
  OAI211_X1 g0178(.A(KEYINPUT7), .B(new_n219), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(KEYINPUT73), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT73), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(new_n375), .C1(new_n281), .C2(G20), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(G68), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G58), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n243), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n201), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n251), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT16), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n281), .A2(new_n375), .A3(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n359), .A2(new_n361), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n392), .B2(new_n219), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n260), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n372), .B(new_n374), .C1(new_n390), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n383), .A2(new_n389), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n258), .A2(new_n220), .A3(new_n259), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n243), .B1(new_n376), .B2(new_n379), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(new_n388), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT74), .B(KEYINPUT17), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n408), .A2(new_n374), .A3(new_n372), .A4(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n400), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n374), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n403), .B2(new_n407), .ZN(new_n414));
  INV_X1    g0214(.A(G169), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n371), .A2(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n366), .A2(G179), .A3(new_n369), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT18), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n418), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n374), .B1(new_n396), .B2(new_n390), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n326), .A2(new_n353), .A3(new_n357), .A4(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n380), .A2(G107), .A3(new_n382), .ZN(new_n427));
  INV_X1    g0227(.A(G97), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n285), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n429), .A2(new_n204), .B1(KEYINPUT75), .B2(KEYINPUT6), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n429), .A2(new_n204), .ZN(new_n431));
  NOR2_X1   g0231(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(KEYINPUT6), .B2(new_n428), .ZN(new_n433));
  OAI211_X1 g0233(.A(G20), .B(new_n430), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n251), .A2(G77), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n427), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n260), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n263), .A2(new_n428), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT76), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n266), .A2(G33), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n265), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n441), .B2(G97), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n359), .A2(new_n361), .A3(G244), .A4(new_n282), .ZN(new_n443));
  NOR2_X1   g0243(.A1(KEYINPUT77), .A2(KEYINPUT4), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n444), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n281), .A2(G244), .A3(new_n282), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n281), .A2(G250), .A3(G1698), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n445), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n287), .ZN(new_n451));
  OR2_X1    g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  NAND2_X1  g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n266), .A2(G45), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(G257), .A3(new_n274), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n452), .B2(new_n453), .ZN(new_n459));
  INV_X1    g0259(.A(G274), .ZN(new_n460));
  INV_X1    g0260(.A(new_n220), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(new_n273), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n451), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n437), .A2(new_n442), .B1(new_n415), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT78), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n450), .A2(new_n468), .A3(new_n287), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n450), .B2(new_n287), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n464), .A2(G179), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT79), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n451), .A2(KEYINPUT78), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n450), .A2(new_n468), .A3(new_n287), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n474), .A2(KEYINPUT79), .A3(new_n475), .A4(new_n472), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n467), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT80), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(new_n475), .A3(new_n472), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT79), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n476), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n467), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n437), .A2(new_n442), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n466), .A2(new_n355), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n469), .A2(new_n470), .A3(new_n464), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n290), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n441), .A2(G87), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n281), .A2(new_n219), .A3(G68), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT19), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n219), .B1(new_n340), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(G87), .B2(new_n205), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n253), .B2(new_n428), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(new_n260), .B1(new_n263), .B2(new_n254), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n455), .A2(KEYINPUT81), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT81), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(new_n266), .A3(G45), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n501), .A2(G250), .A3(new_n274), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n456), .A2(new_n274), .A3(G274), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n500), .A3(new_n505), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n359), .A2(new_n361), .A3(G238), .A4(new_n282), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G116), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT83), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n281), .A2(new_n512), .A3(G244), .A4(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n359), .A2(new_n361), .A3(G244), .A4(G1698), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT83), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n506), .A2(new_n508), .B1(new_n516), .B2(new_n274), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n499), .B1(new_n518), .B2(G190), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(G200), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n292), .ZN(new_n521));
  INV_X1    g0321(.A(new_n254), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n441), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n517), .A2(new_n415), .B1(new_n523), .B2(new_n498), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n479), .A2(new_n485), .A3(new_n490), .A4(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n359), .A2(new_n361), .A3(new_n219), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n281), .A2(new_n529), .A3(new_n219), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n510), .A2(G20), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n219), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n285), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n531), .A2(new_n532), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n532), .B1(new_n531), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n260), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n263), .A2(new_n285), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n541), .B(KEYINPUT25), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n441), .B2(G107), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n359), .A2(new_n361), .A3(G257), .A4(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n359), .A2(new_n361), .A3(G250), .A4(new_n282), .ZN(new_n545));
  AND2_X1   g0345(.A1(KEYINPUT85), .A2(G294), .ZN(new_n546));
  NOR2_X1   g0346(.A1(KEYINPUT85), .A2(G294), .ZN(new_n547));
  OAI21_X1  g0347(.A(G33), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n287), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n459), .A2(new_n287), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G264), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n552), .A3(new_n463), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n287), .A2(new_n549), .B1(new_n551), .B2(G264), .ZN(new_n555));
  AOI21_X1  g0355(.A(G200), .B1(new_n555), .B2(new_n463), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n540), .B(new_n543), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n415), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n292), .A3(new_n463), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n540), .B2(new_n543), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT86), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n540), .A2(new_n543), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n560), .A3(new_n559), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT86), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(new_n557), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n404), .A2(G116), .A3(new_n332), .A4(new_n440), .ZN(new_n569));
  INV_X1    g0369(.A(G116), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n263), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(G20), .B1(G33), .B2(G283), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n358), .A2(G97), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n572), .A2(new_n573), .B1(G20), .B2(new_n570), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n260), .A2(KEYINPUT20), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT20), .B1(new_n260), .B2(new_n574), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n569), .B(new_n571), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n359), .A2(new_n361), .A3(G264), .A4(G1698), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n359), .A2(new_n361), .A3(G257), .A4(new_n282), .ZN(new_n580));
  INV_X1    g0380(.A(G303), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n281), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n582), .A2(new_n287), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n457), .A2(G270), .A3(new_n274), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n463), .ZN(new_n585));
  OAI21_X1  g0385(.A(G200), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT84), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n578), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n551), .A2(G270), .B1(new_n462), .B2(new_n459), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n582), .A2(new_n287), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n290), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT84), .B1(new_n591), .B2(new_n577), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n583), .A2(new_n585), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G190), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n588), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n589), .A2(new_n590), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n577), .A2(new_n596), .A3(G169), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n596), .A2(new_n292), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n577), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n577), .A2(new_n596), .A3(KEYINPUT21), .A4(G169), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n568), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n426), .A2(new_n526), .A3(new_n605), .ZN(G372));
  INV_X1    g0406(.A(new_n412), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n357), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n353), .B2(new_n294), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(new_n424), .ZN(new_n610));
  INV_X1    g0410(.A(new_n320), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n324), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n521), .A2(new_n524), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n525), .A2(new_n615), .A3(new_n483), .A4(new_n467), .ZN(new_n616));
  INV_X1    g0416(.A(new_n525), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n479), .B2(new_n485), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n614), .B(new_n616), .C1(new_n618), .C2(new_n615), .ZN(new_n619));
  INV_X1    g0419(.A(new_n603), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n558), .B1(new_n620), .B2(new_n565), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT87), .B1(new_n526), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n483), .A2(new_n484), .A3(new_n467), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n484), .B1(new_n483), .B2(new_n467), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n489), .A2(new_n290), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n626), .A2(new_n486), .A3(new_n487), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n525), .A4(new_n621), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n619), .B1(new_n623), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n613), .B1(new_n426), .B2(new_n631), .ZN(G369));
  NAND2_X1  g0432(.A1(new_n331), .A2(new_n219), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(G213), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n577), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n604), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n595), .A2(new_n639), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n620), .A3(new_n641), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(G330), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n564), .A2(new_n638), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n563), .A2(new_n567), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n562), .A2(new_n638), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n620), .A2(new_n638), .ZN(new_n652));
  INV_X1    g0452(.A(new_n638), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n568), .A2(new_n652), .B1(new_n562), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(G399));
  INV_X1    g0455(.A(new_n222), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G41), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n266), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n204), .A2(new_n364), .A3(new_n570), .ZN(new_n660));
  INV_X1    g0460(.A(new_n657), .ZN(new_n661));
  OAI22_X1  g0461(.A1(new_n659), .A2(new_n660), .B1(new_n218), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT28), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n630), .A2(new_n623), .ZN(new_n664));
  INV_X1    g0464(.A(new_n619), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT29), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n653), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n471), .A2(new_n465), .ZN(new_n669));
  AOI21_X1  g0469(.A(G179), .B1(new_n589), .B2(new_n590), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n517), .A2(new_n553), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n464), .B1(new_n287), .B2(new_n450), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(new_n555), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(KEYINPUT30), .A3(new_n518), .A4(new_n600), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n515), .A2(new_n513), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n510), .A3(new_n509), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n287), .ZN(new_n679));
  INV_X1    g0479(.A(new_n506), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n507), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n593), .A2(new_n679), .A3(G179), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n673), .A2(new_n555), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n676), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n672), .A2(new_n675), .A3(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n685), .A2(KEYINPUT31), .A3(new_n638), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT31), .B1(new_n685), .B2(new_n638), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n563), .A2(new_n604), .A3(new_n567), .A4(new_n653), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n526), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n525), .A2(new_n483), .A3(new_n467), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n692), .A2(KEYINPUT26), .B1(new_n521), .B2(new_n524), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n615), .B(new_n525), .C1(new_n624), .C2(new_n625), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n693), .B(new_n694), .C1(new_n526), .C2(new_n622), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT29), .B1(new_n696), .B2(new_n638), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n668), .A2(new_n691), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n663), .B1(new_n699), .B2(G1), .ZN(G364));
  NAND2_X1  g0500(.A1(new_n642), .A2(new_n644), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT89), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n262), .A2(new_n271), .A3(G20), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT90), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n659), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n704), .A2(new_n645), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G13), .A2(G33), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n701), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n219), .A2(new_n292), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(G190), .A3(G200), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G50), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n355), .A2(G179), .A3(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n219), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n428), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n714), .A2(new_n355), .A3(G200), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n219), .A2(G179), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(G190), .A3(G200), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n725), .A2(new_n243), .B1(new_n727), .B2(new_n364), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n355), .A3(G200), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n724), .B(new_n728), .C1(G107), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G190), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G159), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT32), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n714), .A2(G190), .A3(new_n290), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n281), .B1(new_n737), .B2(new_n384), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n714), .A2(new_n732), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n738), .B1(G77), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n721), .A2(new_n731), .A3(new_n736), .A4(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n725), .ZN(new_n743));
  XNOR2_X1  g0543(.A(KEYINPUT33), .B(G317), .ZN(new_n744));
  INV_X1    g0544(.A(new_n737), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n743), .A2(new_n744), .B1(new_n745), .B2(G322), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT94), .Z(new_n747));
  OAI21_X1  g0547(.A(new_n392), .B1(new_n727), .B2(new_n581), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT92), .Z(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n720), .A2(G326), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n733), .A2(KEYINPUT93), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n733), .A2(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G329), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n730), .A2(G283), .ZN(new_n757));
  INV_X1    g0557(.A(new_n723), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n546), .A2(new_n547), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n758), .A2(new_n760), .B1(new_n740), .B2(G311), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n751), .A2(new_n756), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n742), .B1(new_n750), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n220), .B1(G20), .B2(new_n415), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n656), .A2(new_n392), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n766), .A2(G355), .B1(new_n570), .B2(new_n656), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n247), .A2(new_n271), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n656), .A2(new_n281), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G45), .B2(new_n218), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n712), .A2(new_n764), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n708), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n713), .A2(new_n765), .A3(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n709), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(G396));
  NAND2_X1  g0576(.A1(new_n269), .A2(new_n638), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n291), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n294), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n294), .A2(new_n638), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n631), .B2(new_n638), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n291), .A2(new_n294), .A3(new_n653), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n631), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n707), .B1(new_n784), .B2(new_n691), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n691), .B2(new_n784), .ZN(new_n786));
  INV_X1    g0586(.A(new_n727), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n392), .B1(new_n787), .B2(G50), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n788), .B1(new_n384), .B2(new_n723), .C1(new_n243), .C2(new_n729), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n745), .A2(G143), .B1(new_n740), .B2(G159), .ZN(new_n790));
  INV_X1    g0590(.A(G150), .ZN(new_n791));
  INV_X1    g0591(.A(G137), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n790), .B1(new_n791), .B2(new_n725), .C1(new_n719), .C2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT34), .Z(new_n794));
  AOI211_X1 g0594(.A(new_n789), .B(new_n794), .C1(G132), .C2(new_n755), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n281), .B1(new_n740), .B2(G116), .ZN(new_n796));
  INV_X1    g0596(.A(G294), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n797), .B2(new_n737), .C1(new_n754), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n729), .A2(new_n364), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n724), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n285), .B2(new_n727), .C1(new_n802), .C2(new_n725), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n799), .B(new_n803), .C1(G303), .C2(new_n720), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n764), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n764), .A2(new_n710), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n708), .B1(new_n261), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n781), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n805), .B(new_n807), .C1(new_n808), .C2(new_n711), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n786), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G384));
  NOR3_X1   g0611(.A1(new_n220), .A2(new_n219), .A3(new_n570), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n430), .B1(new_n431), .B2(new_n433), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT35), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT36), .ZN(new_n817));
  OR3_X1    g0617(.A1(new_n218), .A2(new_n261), .A3(new_n385), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n266), .B(G13), .C1(new_n818), .C2(new_n242), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n426), .B1(new_n668), .B2(new_n697), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n612), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n402), .B1(new_n405), .B2(new_n388), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n395), .A2(new_n823), .A3(new_n260), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n636), .B1(new_n824), .B2(new_n374), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n412), .B2(new_n424), .ZN(new_n826));
  INV_X1    g0626(.A(new_n397), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n418), .A2(new_n636), .B1(new_n374), .B2(new_n824), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT37), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT95), .B1(new_n414), .B2(new_n418), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT95), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n420), .A2(new_n421), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n636), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n421), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n836), .A3(new_n397), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n829), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n826), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n826), .A2(KEYINPUT38), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n338), .A2(new_n638), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n357), .A2(new_n353), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n338), .B(new_n638), .C1(new_n351), .C2(new_n352), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n783), .B1(new_n664), .B2(new_n665), .ZN(new_n848));
  INV_X1    g0648(.A(new_n780), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n843), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT39), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT96), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n826), .A2(new_n838), .A3(new_n852), .A4(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n842), .A2(KEYINPUT96), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n397), .B1(new_n414), .B2(new_n418), .ZN(new_n855));
  INV_X1    g0655(.A(new_n835), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT37), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n837), .B2(new_n833), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n856), .B1(new_n412), .B2(new_n424), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT38), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n851), .B(new_n853), .C1(new_n854), .C2(new_n860), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n353), .A2(new_n638), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(new_n843), .C2(new_n851), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n424), .A2(new_n636), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n850), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n822), .B(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT97), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n526), .A2(new_n689), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n685), .A2(new_n638), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT31), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n685), .A2(KEYINPUT31), .A3(new_n638), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n868), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n688), .B(KEYINPUT97), .C1(new_n526), .C2(new_n689), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n781), .B1(new_n845), .B2(new_n846), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n853), .B1(new_n854), .B2(new_n860), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT40), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT40), .B1(new_n841), .B2(new_n842), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n881), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n875), .A2(new_n876), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n426), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n883), .A2(new_n885), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n886), .A2(new_n887), .A3(new_n702), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n867), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(G1), .B1(new_n262), .B2(G20), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n867), .B2(new_n888), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n820), .B1(new_n889), .B2(new_n891), .ZN(G367));
  INV_X1    g0692(.A(new_n769), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n235), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n772), .B1(new_n222), .B2(new_n254), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n707), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n720), .A2(G143), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n739), .A2(new_n241), .B1(new_n733), .B2(new_n792), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n392), .B(new_n898), .C1(G150), .C2(new_n745), .ZN(new_n899));
  AOI22_X1  g0699(.A1(G159), .A2(new_n743), .B1(new_n730), .B2(G77), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n758), .A2(G68), .B1(new_n787), .B2(G58), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n897), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT105), .ZN(new_n903));
  XNOR2_X1  g0703(.A(KEYINPUT104), .B(G317), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n392), .B1(new_n733), .B2(new_n904), .C1(new_n428), .C2(new_n729), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n720), .A2(G311), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n787), .A2(G116), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT46), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n737), .A2(new_n581), .B1(new_n739), .B2(new_n802), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(G107), .B2(new_n758), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n909), .B(new_n911), .C1(new_n759), .C2(new_n725), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n902), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT47), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n896), .B1(new_n914), .B2(new_n764), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n499), .A2(new_n638), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n525), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n614), .A2(new_n916), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n712), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n706), .A2(new_n266), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n645), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT101), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n647), .B(new_n648), .C1(new_n620), .C2(new_n638), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT100), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n568), .A2(new_n652), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT101), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n930), .B2(new_n645), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n924), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n927), .A2(new_n924), .A3(new_n931), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n699), .A2(new_n935), .A3(KEYINPUT102), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT102), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n927), .A2(new_n924), .A3(new_n931), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(new_n932), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n939), .B2(new_n698), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n486), .A2(new_n638), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n628), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n483), .A2(new_n467), .A3(new_n638), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n654), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(KEYINPUT45), .A3(new_n654), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(KEYINPUT44), .A3(new_n948), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT44), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n946), .B2(new_n654), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n951), .A2(new_n955), .A3(new_n651), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n651), .B1(new_n951), .B2(new_n955), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT103), .B1(new_n941), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n956), .A2(new_n957), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT103), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(new_n936), .A3(new_n940), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n699), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n657), .B(KEYINPUT41), .Z(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n922), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n946), .A2(new_n929), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT42), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n947), .A2(new_n565), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n479), .A2(new_n485), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n969), .B1(new_n653), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n917), .A2(new_n918), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT98), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT99), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n973), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n651), .A2(new_n947), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n981), .A2(new_n985), .A3(new_n983), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n920), .B1(new_n967), .B2(new_n989), .ZN(G387));
  XNOR2_X1  g0790(.A(new_n657), .B(KEYINPUT109), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n941), .B(new_n991), .C1(new_n699), .C2(new_n935), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n720), .A2(G159), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n737), .A2(new_n241), .B1(new_n739), .B2(new_n243), .ZN(new_n994));
  INV_X1    g0794(.A(new_n733), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n392), .B(new_n994), .C1(G150), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n727), .A2(new_n261), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G97), .B2(new_n730), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n723), .A2(new_n254), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n250), .B2(new_n743), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n993), .A2(new_n996), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(G322), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n719), .A2(new_n1002), .B1(new_n798), .B2(new_n725), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1003), .A2(KEYINPUT107), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n737), .A2(new_n904), .B1(new_n739), .B2(new_n581), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT107), .B2(new_n1003), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT48), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n758), .A2(G283), .B1(new_n787), .B2(new_n760), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT108), .Z(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT49), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n281), .B1(new_n995), .B2(G326), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n570), .C2(new_n729), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1013), .A2(KEYINPUT49), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1001), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n764), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n649), .A2(new_n712), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n766), .A2(new_n660), .B1(new_n285), .B2(new_n656), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n231), .A2(new_n271), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n249), .A2(G50), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  AOI211_X1 g0825(.A(G45), .B(new_n660), .C1(G68), .C2(G77), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n769), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1021), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n708), .B1(new_n1029), .B2(new_n772), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1019), .A2(new_n1020), .A3(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n992), .B(new_n1031), .C1(new_n939), .C2(new_n921), .ZN(G393));
  INV_X1    g0832(.A(new_n991), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n941), .B2(new_n958), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n963), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n947), .A2(new_n712), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n772), .B1(new_n428), .B2(new_n222), .C1(new_n240), .C2(new_n893), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n707), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n720), .A2(G317), .B1(G311), .B2(new_n745), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT52), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n392), .B1(new_n733), .B2(new_n1002), .C1(new_n797), .C2(new_n739), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n725), .A2(new_n581), .B1(new_n729), .B2(new_n285), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n723), .A2(new_n570), .B1(new_n727), .B2(new_n802), .ZN(new_n1043));
  OR3_X1    g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n719), .A2(new_n791), .B1(new_n734), .B2(new_n737), .ZN(new_n1045));
  XOR2_X1   g0845(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n740), .A2(new_n250), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n392), .B1(new_n995), .B2(G143), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n725), .A2(new_n241), .B1(new_n727), .B2(new_n243), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n800), .B(new_n1051), .C1(G77), .C2(new_n758), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1040), .A2(new_n1044), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1038), .B1(new_n1054), .B2(new_n764), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n960), .A2(new_n922), .B1(new_n1036), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT111), .B1(new_n1035), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT111), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1056), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n963), .C2(new_n1034), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1057), .A2(new_n1060), .ZN(G390));
  OAI22_X1  g0861(.A1(new_n243), .A2(new_n729), .B1(new_n727), .B2(new_n364), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n754), .A2(new_n797), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n723), .A2(new_n261), .B1(new_n725), .B2(new_n285), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n392), .B1(new_n739), .B2(new_n428), .C1(new_n570), .C2(new_n737), .ZN(new_n1065));
  OR4_X1    g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n719), .A2(new_n802), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n755), .A2(G125), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT54), .B(G143), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n739), .A2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n392), .B(new_n1070), .C1(G132), .C2(new_n745), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n730), .A2(G50), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G159), .A2(new_n758), .B1(new_n743), .B2(G137), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(new_n1071), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n727), .A2(new_n791), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(G128), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n719), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1066), .A2(new_n1067), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n764), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n708), .B1(new_n249), .B2(new_n806), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n861), .B1(new_n843), .B2(new_n851), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1081), .B(new_n1082), .C1(new_n1084), .C2(new_n711), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n862), .B(new_n853), .C1(new_n854), .C2(new_n860), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n847), .B(KEYINPUT112), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n695), .A2(new_n653), .A3(new_n779), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n780), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n690), .A2(new_n847), .A3(G330), .A4(new_n808), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n780), .B1(new_n631), .B2(new_n783), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n863), .B1(new_n1093), .B2(new_n847), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1091), .B(new_n1092), .C1(new_n1094), .C2(new_n1084), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n783), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n849), .B1(new_n666), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n847), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n862), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1090), .B1(new_n1099), .B2(new_n1083), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n875), .A2(new_n876), .A3(G330), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n877), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1095), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1085), .B1(new_n1104), .B2(new_n921), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1091), .B1(new_n1094), .B2(new_n1084), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n877), .A3(new_n1102), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1098), .B1(new_n691), .B2(new_n781), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1093), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT112), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n847), .B(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1101), .B2(new_n781), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1092), .A2(new_n780), .A3(new_n1088), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT113), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1115), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1110), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n426), .A2(new_n1101), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n821), .A2(new_n612), .A3(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1107), .A2(new_n1119), .A3(new_n1095), .A4(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1122), .A2(new_n991), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1104), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1105), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(G378));
  AOI21_X1  g0927(.A(new_n708), .B1(new_n241), .B2(new_n806), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n725), .A2(new_n428), .B1(new_n729), .B2(new_n384), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n997), .B(new_n1129), .C1(G68), .C2(new_n758), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n281), .A2(G41), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n739), .B2(new_n254), .C1(new_n285), .C2(new_n737), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n755), .B2(G283), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1130), .B(new_n1133), .C1(new_n570), .C2(new_n719), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT58), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n737), .A2(new_n1078), .B1(new_n739), .B2(new_n792), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G132), .B2(new_n743), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1069), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n758), .A2(G150), .B1(new_n787), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(G125), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1137), .B(new_n1139), .C1(new_n1140), .C2(new_n719), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT115), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1144), .A2(G124), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(G124), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n995), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1147), .A2(new_n358), .A3(new_n270), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1143), .B(new_n1148), .C1(new_n734), .C2(new_n729), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n241), .B1(G33), .B2(G41), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1135), .B1(new_n1142), .B2(new_n1149), .C1(new_n1131), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1151), .A2(KEYINPUT116), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(KEYINPUT116), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n764), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n311), .A2(new_n636), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n325), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1155), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n320), .A2(new_n324), .A3(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1159), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1157), .B1(new_n320), .B2(new_n324), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1155), .B(new_n323), .C1(new_n317), .C2(new_n319), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1160), .A2(new_n1164), .A3(KEYINPUT117), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT117), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1128), .B1(new_n1152), .B2(new_n1154), .C1(new_n1168), .C2(new_n711), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT118), .Z(new_n1170));
  NAND2_X1  g0970(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n883), .B2(G330), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n702), .B(new_n1167), .C1(new_n880), .C2(new_n882), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n866), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n883), .A2(G330), .A3(new_n1168), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n850), .A2(new_n864), .A3(new_n865), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n702), .B1(new_n880), .B2(new_n882), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(new_n1176), .C1(new_n1177), .C2(new_n1171), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT119), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT119), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1174), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1170), .B1(new_n1183), .B2(new_n922), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT113), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1186), .A2(new_n1116), .B1(new_n1109), .B2(new_n1093), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1121), .B1(new_n1104), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT120), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT120), .B1(new_n1192), .B2(new_n1176), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1188), .B(KEYINPUT57), .C1(new_n1191), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n991), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1184), .B1(new_n1189), .B2(new_n1195), .ZN(G375));
  INV_X1    g0996(.A(new_n1121), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1187), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n1124), .A3(new_n966), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n708), .B1(new_n243), .B2(new_n806), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n725), .A2(new_n570), .B1(new_n727), .B2(new_n428), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n999), .B(new_n1201), .C1(G77), .C2(new_n730), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n392), .B1(new_n739), .B2(new_n285), .C1(new_n802), .C2(new_n737), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n755), .B2(G303), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n797), .C2(new_n719), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT121), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n720), .A2(G132), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n723), .A2(new_n241), .B1(new_n729), .B2(new_n384), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n725), .A2(new_n1069), .B1(new_n727), .B2(new_n734), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n755), .A2(G128), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n281), .B1(new_n737), .B2(new_n792), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G150), .B2(new_n740), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1207), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1206), .A2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT122), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(KEYINPUT122), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n764), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1200), .B1(new_n1216), .B2(new_n1218), .C1(new_n1087), .C2(new_n711), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n1187), .B2(new_n921), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1199), .A2(new_n1221), .ZN(G381));
  AND3_X1   g1022(.A1(new_n981), .A2(new_n985), .A3(new_n983), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n985), .B1(new_n981), .B2(new_n983), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n698), .B1(new_n959), .B2(new_n962), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n921), .B1(new_n1226), .B2(new_n965), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1225), .A2(new_n1227), .B1(new_n919), .B2(new_n915), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT123), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT123), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1126), .B(new_n1184), .C1(new_n1189), .C2(new_n1195), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .ZN(G407));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G343), .C2(new_n1234), .ZN(G409));
  INV_X1    g1037(.A(KEYINPUT60), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1198), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n991), .A3(new_n1124), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT124), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1198), .B2(new_n1238), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1187), .A2(KEYINPUT124), .A3(KEYINPUT60), .A4(new_n1197), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n810), .B1(new_n1244), .B2(new_n1220), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G384), .B(new_n1221), .C1(new_n1246), .C2(new_n1240), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n637), .A2(G213), .A3(G2897), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1245), .A2(new_n1247), .A3(new_n1249), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n922), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1126), .A2(new_n1169), .A3(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1180), .A2(new_n1182), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n966), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1255), .A2(new_n1257), .B1(G213), .B2(new_n637), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G375), .A2(G378), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G390), .A2(new_n1228), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1229), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT125), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(G393), .B(new_n775), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT125), .B1(G390), .B2(new_n1228), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1268), .A2(new_n1265), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1248), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1261), .A2(new_n1270), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1260), .A2(new_n1252), .A3(new_n1251), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1271), .A2(new_n1258), .A3(new_n1280), .A4(new_n1259), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .A4(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1263), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(G387), .A2(new_n1229), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1264), .B1(G387), .B2(new_n1229), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1265), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n1283), .A2(new_n1284), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1266), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1282), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1276), .A2(new_n1289), .ZN(G405));
  OAI211_X1 g1090(.A(new_n991), .B(new_n1194), .C1(new_n1256), .C2(KEYINPUT57), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1126), .B1(new_n1291), .B2(new_n1184), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT126), .B1(new_n1235), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1259), .A2(new_n1294), .A3(new_n1234), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1271), .A3(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1248), .B1(new_n1235), .B2(new_n1292), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1293), .A2(new_n1298), .A3(new_n1295), .A4(new_n1271), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1300), .A2(new_n1288), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1288), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(G402));
endmodule


