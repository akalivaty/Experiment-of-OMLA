//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n207), .A2(new_n208), .B1(G155gat), .B2(G162gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G141gat), .B(G148gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(G155gat), .B2(G162gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n206), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT2), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT76), .B1(new_n216), .B2(new_n217), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n215), .B(new_n218), .C1(new_n205), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G211gat), .A2(G218gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G211gat), .A2(G218gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(G197gat), .A2(G204gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G197gat), .A2(G204gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(G197gat), .B(G204gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n229), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT73), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n230), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  OAI211_X1 g036(.A(KEYINPUT73), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n222), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n212), .A2(new_n220), .A3(new_n240), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n242), .A2(new_n243), .B1(new_n236), .B2(new_n238), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n204), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT79), .ZN(new_n246));
  INV_X1    g045(.A(new_n243), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n247), .B1(new_n230), .B2(new_n234), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n221), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT78), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n242), .A2(new_n243), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT78), .B(new_n221), .C1(new_n248), .C2(KEYINPUT3), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n252), .A2(new_n255), .A3(new_n203), .A4(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n245), .A2(new_n246), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n246), .B1(new_n245), .B2(new_n257), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n202), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT79), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n257), .ZN(new_n263));
  INV_X1    g062(.A(new_n202), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(G22gat), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n260), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n260), .B2(new_n265), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n254), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT23), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT65), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n279));
  INV_X1    g078(.A(new_n278), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT23), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n277), .A2(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  AND2_X1   g083(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT64), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n287), .B2(new_n289), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT25), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n289), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n295), .B(new_n296), .C1(G183gat), .C2(G190gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT66), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT23), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n282), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n297), .A2(new_n301), .A3(KEYINPUT25), .A4(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n278), .B1(new_n305), .B2(new_n281), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n298), .A2(new_n300), .A3(new_n305), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT67), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n298), .A2(new_n300), .A3(new_n309), .A4(new_n305), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  INV_X1    g111(.A(G190gat), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT28), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT27), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  AND4_X1   g117(.A1(KEYINPUT28), .A2(new_n316), .A3(new_n318), .A4(new_n313), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n287), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n294), .A2(new_n304), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n310), .ZN(new_n325));
  INV_X1    g124(.A(new_n306), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n287), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n312), .A2(KEYINPUT28), .A3(new_n313), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT25), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n278), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT65), .B1(new_n278), .B2(KEYINPUT23), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n302), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n296), .B1(G183gat), .B2(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n295), .A2(KEYINPUT64), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(new_n290), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n335), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n303), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT29), .B1(new_n334), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n272), .B(new_n324), .C1(new_n344), .C2(new_n323), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n323), .B1(new_n321), .B2(new_n243), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n321), .A2(new_n348), .A3(new_n323), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n345), .B1(new_n350), .B2(new_n272), .ZN(new_n351));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(G64gat), .B(G92gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n321), .A2(new_n243), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n322), .ZN(new_n358));
  INV_X1    g157(.A(new_n349), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n348), .B1(new_n321), .B2(new_n323), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n254), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n354), .A3(new_n345), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n356), .A2(new_n363), .A3(KEYINPUT30), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n362), .A2(new_n365), .A3(new_n354), .A4(new_n345), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT40), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT39), .ZN(new_n370));
  INV_X1    g169(.A(G113gat), .ZN(new_n371));
  INV_X1    g170(.A(G120gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G113gat), .A2(G120gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT69), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT1), .ZN(new_n377));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT69), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n379), .A3(new_n374), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n376), .A2(new_n377), .A3(new_n378), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(KEYINPUT68), .ZN(new_n382));
  INV_X1    g181(.A(G127gat), .ZN(new_n383));
  OR3_X1    g182(.A1(new_n383), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n373), .A2(new_n377), .A3(new_n374), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n381), .A2(new_n386), .A3(new_n220), .A4(new_n212), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n381), .A2(new_n386), .B1(new_n220), .B2(new_n212), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n387), .B(KEYINPUT4), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n381), .A2(new_n386), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n250), .A2(new_n242), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n370), .B(new_n392), .C1(new_n396), .C2(new_n390), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n370), .A3(new_n390), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n369), .B1(new_n397), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n390), .B1(new_n388), .B2(new_n391), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT5), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n388), .A2(KEYINPUT4), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n387), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n407), .A2(new_n395), .A3(new_n409), .A4(new_n389), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n393), .A2(KEYINPUT5), .A3(new_n389), .A4(new_n395), .ZN(new_n412));
  INV_X1    g211(.A(new_n402), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n404), .A2(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n397), .A2(new_n403), .A3(new_n369), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n271), .B1(new_n368), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n358), .B(new_n272), .C1(new_n359), .C2(new_n360), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT37), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n323), .B1(new_n321), .B2(new_n237), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n322), .B1(new_n334), .B2(new_n343), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n254), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n424), .A2(new_n420), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT38), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n427), .B(new_n355), .C1(new_n351), .C2(KEYINPUT37), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n412), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n402), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n414), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT6), .A4(new_n413), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n363), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT81), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n351), .A2(KEYINPUT37), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n355), .B1(new_n351), .B2(KEYINPUT37), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT38), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n429), .A2(new_n435), .A3(KEYINPUT81), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n418), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n394), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n321), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n334), .A2(new_n343), .A3(new_n394), .ZN(new_n445));
  INV_X1    g244(.A(G227gat), .ZN(new_n446));
  INV_X1    g245(.A(G233gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT70), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(G15gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G43gat), .ZN(new_n455));
  INV_X1    g254(.A(G15gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n453), .B(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(G43gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n451), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n444), .A2(new_n445), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT34), .B1(new_n463), .B2(new_n448), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n448), .B1(new_n444), .B2(new_n445), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n449), .A2(KEYINPUT32), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n460), .B1(new_n449), .B2(new_n450), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n465), .A2(new_n466), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT34), .B(new_n448), .C1(new_n444), .C2(new_n445), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n468), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n468), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT72), .B1(new_n477), .B2(KEYINPUT36), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT72), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT36), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n479), .B(new_n480), .C1(new_n475), .C2(new_n476), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT71), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(new_n483), .A3(KEYINPUT36), .ZN(new_n484));
  INV_X1    g283(.A(new_n474), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n469), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n470), .A3(new_n474), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(KEYINPUT36), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT71), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n433), .A2(new_n434), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n367), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n367), .A2(KEYINPUT77), .A3(new_n493), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n271), .A3(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n442), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n260), .A2(new_n265), .ZN(new_n500));
  INV_X1    g299(.A(new_n267), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n260), .A2(new_n265), .A3(new_n267), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n502), .A3(new_n503), .A4(new_n488), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n494), .A2(new_n504), .A3(KEYINPUT35), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(KEYINPUT82), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT82), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n477), .B2(new_n270), .ZN(new_n508));
  AOI221_X4 g307(.A(new_n495), .B1(new_n433), .B2(new_n434), .C1(new_n364), .C2(new_n366), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT77), .B1(new_n367), .B2(new_n493), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n506), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT83), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(KEYINPUT83), .A3(KEYINPUT35), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n499), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT16), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(G1gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(G1gat), .B2(new_n517), .ZN(new_n520));
  INV_X1    g319(.A(G8gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT85), .B(G50gat), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n458), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n524), .A2(new_n525), .B1(new_n528), .B2(KEYINPUT86), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530));
  OR2_X1    g329(.A1(G43gat), .A2(G50gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(G43gat), .A2(G50gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n529), .B(new_n534), .C1(KEYINPUT86), .C2(new_n528), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n528), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n533), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n536), .B1(new_n535), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n522), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n522), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n535), .A2(new_n540), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT18), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(KEYINPUT87), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(KEYINPUT87), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT18), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n522), .A2(new_n540), .A3(new_n535), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n544), .B(KEYINPUT13), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT12), .ZN(new_n562));
  AND4_X1   g361(.A1(new_n550), .A2(new_n552), .A3(new_n556), .A4(new_n562), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n551), .A2(KEYINPUT18), .B1(new_n554), .B2(new_n555), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n564), .B2(new_n550), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n516), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT89), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT7), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n570), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n574), .B1(new_n568), .B2(new_n569), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G99gat), .B(G106gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n577), .A3(new_n575), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n546), .A2(new_n582), .B1(KEYINPUT41), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n541), .A2(new_n542), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT90), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n581), .B(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n584), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT91), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n595), .B(new_n584), .C1(new_n585), .C2(new_n587), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n591), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n594), .B1(new_n591), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G57gat), .B(G64gat), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G71gat), .B(G78gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n606));
  XOR2_X1   g405(.A(G127gat), .B(G155gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n545), .B1(KEYINPUT21), .B2(new_n605), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT88), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n610), .A2(new_n616), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n603), .B(new_n604), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n581), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n605), .A2(new_n579), .A3(new_n580), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n582), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n622), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n626), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(new_n622), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(KEYINPUT92), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT92), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n627), .A2(new_n628), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n621), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n630), .A2(new_n622), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n634), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n620), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n567), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n493), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n368), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  OAI21_X1  g452(.A(G8gat), .B1(new_n653), .B2(new_n367), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n652), .ZN(new_n655));
  MUX2_X1   g454(.A(new_n652), .B(new_n655), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g455(.A(G15gat), .B1(new_n653), .B2(new_n492), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n647), .A2(new_n456), .A3(new_n477), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(G1326gat));
  NOR3_X1   g458(.A1(new_n516), .A2(new_n566), .A3(new_n270), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n646), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  NOR3_X1   g462(.A1(new_n600), .A2(new_n619), .A3(new_n645), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n567), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n537), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n665), .A2(KEYINPUT93), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT93), .B1(new_n665), .B2(new_n666), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n667), .A2(KEYINPUT45), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT45), .B1(new_n667), .B2(new_n668), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n619), .B(KEYINPUT94), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n566), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n645), .B(KEYINPUT95), .Z(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n504), .A2(KEYINPUT82), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n477), .A2(new_n270), .A3(new_n507), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n496), .A2(new_n497), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT35), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n513), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n505), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n515), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n442), .A2(new_n492), .A3(new_n498), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n600), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n677), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(KEYINPUT96), .B(KEYINPUT44), .C1(new_n516), .C2(new_n600), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n516), .A2(KEYINPUT97), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n684), .A2(new_n685), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT97), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n691), .A2(new_n694), .A3(new_n687), .A4(new_n599), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n676), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(new_n648), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT98), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n671), .B1(new_n699), .B2(new_n700), .ZN(G1328gat));
  NOR3_X1   g500(.A1(new_n665), .A2(G36gat), .A3(new_n367), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT46), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n696), .A2(new_n368), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G36gat), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(G1329gat));
  NOR2_X1   g507(.A1(new_n492), .A2(new_n458), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n567), .A2(new_n477), .A3(new_n664), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n696), .A2(new_n709), .B1(new_n710), .B2(new_n458), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g511(.A(new_n523), .B1(new_n696), .B2(new_n271), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n660), .A2(new_n523), .A3(new_n664), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n714), .B1(new_n713), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1331gat));
  AND2_X1   g518(.A1(new_n691), .A2(new_n694), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n675), .A2(new_n674), .A3(new_n620), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT100), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n493), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT101), .B(G57gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1332gat));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n720), .A2(KEYINPUT102), .A3(new_n722), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n367), .B(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n728), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n734), .B(new_n735), .Z(G1333gat));
  INV_X1    g535(.A(new_n492), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n728), .A2(G71gat), .A3(new_n737), .A4(new_n729), .ZN(new_n738));
  INV_X1    g537(.A(G71gat), .ZN(new_n739));
  INV_X1    g538(.A(new_n477), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n723), .B2(new_n740), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n738), .A2(KEYINPUT50), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT50), .B1(new_n738), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(G1334gat));
  AND2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n271), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G78gat), .ZN(new_n747));
  INV_X1    g546(.A(G78gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n748), .A3(new_n271), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n674), .A2(new_n619), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n645), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n690), .B2(new_n695), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(new_n648), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n686), .A2(new_n751), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n756), .A2(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(KEYINPUT51), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n686), .A2(new_n751), .B1(new_n756), .B2(KEYINPUT51), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n645), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n648), .A2(new_n568), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n754), .A2(new_n568), .B1(new_n762), .B2(new_n763), .ZN(G1336gat));
  AOI21_X1  g563(.A(new_n569), .B1(new_n753), .B2(new_n368), .ZN(new_n765));
  INV_X1    g564(.A(new_n675), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n732), .A2(G92gat), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n766), .B(new_n767), .C1(new_n760), .C2(new_n761), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n690), .A2(new_n695), .ZN(new_n772));
  INV_X1    g571(.A(new_n752), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n731), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n768), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n771), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n569), .B1(new_n753), .B2(new_n731), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n780), .A2(KEYINPUT105), .A3(new_n777), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n770), .B1(new_n779), .B2(new_n781), .ZN(G1337gat));
  AND2_X1   g581(.A1(new_n753), .A2(new_n737), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT106), .B(G99gat), .Z(new_n784));
  NAND2_X1  g583(.A1(new_n477), .A2(new_n784), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n783), .A2(new_n784), .B1(new_n762), .B2(new_n785), .ZN(G1338gat));
  INV_X1    g585(.A(new_n760), .ZN(new_n787));
  INV_X1    g586(.A(new_n761), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n675), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(G106gat), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(new_n790), .A3(new_n271), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n753), .B2(new_n271), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT53), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n790), .A3(new_n271), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n753), .A2(new_n271), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n790), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(G1339gat));
  INV_X1    g597(.A(new_n645), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n566), .A2(new_n619), .A3(new_n600), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT107), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n544), .B1(new_n543), .B2(new_n547), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n554), .A2(new_n555), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n561), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT108), .B(new_n561), .C1(new_n802), .C2(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n564), .A2(new_n550), .A3(new_n562), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n645), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n637), .A2(new_n621), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n812), .A2(new_n813), .A3(new_n629), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n634), .B1(new_n629), .B2(new_n813), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n811), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n629), .A2(new_n813), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n637), .B2(new_n621), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n815), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n643), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n810), .B1(new_n566), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT110), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n815), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n824), .A2(new_n811), .B1(new_n635), .B2(new_n642), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(new_n820), .C1(new_n563), .C2(new_n565), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n810), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n600), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n825), .A2(new_n599), .A3(new_n820), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n809), .A2(new_n808), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n832), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n643), .A2(new_n817), .A3(new_n820), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n834), .A2(KEYINPUT109), .A3(new_n599), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n829), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n801), .B1(new_n839), .B2(new_n673), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n493), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n678), .A2(new_n679), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n731), .ZN(new_n844));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n674), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n800), .B(KEYINPUT107), .Z(new_n846));
  AOI21_X1  g645(.A(new_n599), .B1(new_n822), .B2(KEYINPUT110), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n837), .B1(new_n847), .B2(new_n828), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(new_n672), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n270), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n731), .A2(new_n493), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n477), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n566), .A2(new_n371), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  AOI21_X1  g657(.A(G120gat), .B1(new_n844), .B2(new_n645), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n675), .A2(new_n372), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n856), .B2(new_n860), .ZN(G1341gat));
  INV_X1    g660(.A(new_n856), .ZN(new_n862));
  OAI21_X1  g661(.A(G127gat), .B1(new_n862), .B2(new_n673), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n383), .A3(new_n619), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1342gat));
  OAI21_X1  g664(.A(G134gat), .B1(new_n862), .B2(new_n600), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n600), .A2(new_n368), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n843), .A2(G134gat), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT56), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n870), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n492), .A2(new_n271), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT113), .Z(new_n873));
  AND3_X1   g672(.A1(new_n841), .A2(new_n732), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n566), .A2(G141gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n492), .A2(new_n854), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n849), .B2(new_n271), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n270), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n619), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n599), .B1(new_n826), .B2(new_n810), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT112), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n833), .B(new_n836), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n822), .A2(new_n600), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(KEYINPUT112), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n883), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n882), .B1(new_n889), .B2(new_n846), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n674), .B(new_n878), .C1(new_n879), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G141gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n876), .B2(new_n892), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT114), .B1(new_n891), .B2(G141gat), .ZN(new_n897));
  OAI22_X1  g696(.A1(new_n895), .A2(new_n896), .B1(KEYINPUT58), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n896), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n897), .A2(KEYINPUT58), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n894), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(G1344gat));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n645), .B(new_n878), .C1(new_n879), .C2(new_n890), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n905));
  INV_X1    g704(.A(G148gat), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(KEYINPUT59), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n905), .B1(new_n904), .B2(new_n907), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n672), .B1(new_n829), .B2(new_n838), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n881), .B1(new_n911), .B2(new_n801), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n831), .A2(new_n832), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n887), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT118), .B1(new_n884), .B2(new_n914), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n917), .A3(new_n883), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n270), .B1(new_n918), .B2(new_n800), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n912), .B1(new_n919), .B2(KEYINPUT57), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n877), .A2(new_n799), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n910), .B1(new_n922), .B2(G148gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n908), .A2(new_n909), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n799), .A2(G148gat), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n841), .A2(new_n732), .A3(new_n873), .A4(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT116), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n903), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n921), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n918), .A2(new_n800), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n271), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n880), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n912), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT59), .B1(new_n934), .B2(new_n906), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n904), .A2(new_n907), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n905), .ZN(new_n937));
  OAI211_X1 g736(.A(KEYINPUT119), .B(new_n927), .C1(new_n937), .C2(new_n908), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n929), .A2(new_n938), .ZN(G1345gat));
  NAND3_X1  g738(.A1(new_n874), .A2(new_n216), .A3(new_n619), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n880), .B1(new_n840), .B2(new_n270), .ZN(new_n941));
  INV_X1    g740(.A(new_n890), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n877), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(new_n672), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n944), .B2(new_n216), .ZN(G1346gat));
  AOI21_X1  g744(.A(new_n217), .B1(new_n943), .B2(new_n599), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n841), .A2(new_n873), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n868), .A2(G162gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n949), .B(new_n950), .ZN(G1347gat));
  NOR2_X1   g750(.A1(new_n840), .A2(new_n648), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n842), .A2(new_n731), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G169gat), .B1(new_n955), .B2(new_n674), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n648), .A2(new_n367), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n477), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n958), .B1(new_n851), .B2(new_n852), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n566), .A2(new_n273), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1348gat));
  OAI21_X1  g760(.A(new_n274), .B1(new_n954), .B2(new_n799), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT121), .Z(new_n963));
  NOR2_X1   g762(.A1(new_n675), .A2(new_n274), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n959), .B2(new_n964), .ZN(G1349gat));
  AOI21_X1  g764(.A(new_n315), .B1(new_n959), .B2(new_n672), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n955), .A2(new_n312), .A3(new_n619), .ZN(new_n967));
  OR3_X1    g766(.A1(new_n966), .A2(KEYINPUT60), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(KEYINPUT60), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1350gat));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n313), .A3(new_n599), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n959), .A2(new_n599), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(G190gat), .ZN(new_n974));
  AOI211_X1 g773(.A(KEYINPUT61), .B(new_n313), .C1(new_n959), .C2(new_n599), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(G1351gat));
  NOR2_X1   g775(.A1(new_n872), .A2(new_n732), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n952), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g777(.A1(new_n566), .A2(G197gat), .ZN(new_n979));
  OR3_X1    g778(.A1(new_n978), .A2(KEYINPUT122), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(KEYINPUT122), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n492), .A2(new_n957), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n983), .B1(new_n933), .B2(new_n912), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(new_n674), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(G197gat), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT123), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n987), .B(new_n988), .ZN(G1352gat));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n991));
  INV_X1    g790(.A(G204gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n992), .B1(new_n990), .B2(KEYINPUT124), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n799), .A2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  OR3_X1    g794(.A1(new_n978), .A2(new_n991), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n991), .B1(new_n978), .B2(new_n995), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n992), .B1(new_n984), .B2(new_n766), .ZN(new_n999));
  OR3_X1    g798(.A1(new_n998), .A2(KEYINPUT125), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g799(.A(KEYINPUT125), .B1(new_n998), .B2(new_n999), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1353gat));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n619), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1003), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(KEYINPUT63), .B1(new_n1003), .B2(G211gat), .ZN(new_n1005));
  OR2_X1    g804(.A1(new_n883), .A2(G211gat), .ZN(new_n1006));
  OAI22_X1  g805(.A1(new_n1004), .A2(new_n1005), .B1(new_n978), .B2(new_n1006), .ZN(G1354gat));
  INV_X1    g806(.A(G218gat), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1008), .B1(new_n978), .B2(new_n600), .ZN(new_n1009));
  OR2_X1    g808(.A1(new_n1009), .A2(KEYINPUT126), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n984), .A2(G218gat), .A3(new_n599), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(KEYINPUT126), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(KEYINPUT127), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1015));
  NAND4_X1  g814(.A1(new_n1010), .A2(new_n1015), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1014), .A2(new_n1016), .ZN(G1355gat));
endmodule


