//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n192), .B(KEYINPUT64), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n188), .A2(new_n190), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(new_n191), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n196), .A2(new_n197), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT65), .A2(G134), .ZN(new_n206));
  AOI21_X1  g020(.A(G137), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT66), .B1(new_n207), .B2(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT65), .A2(G134), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT65), .A2(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n205), .A2(new_n206), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(new_n209), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n202), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  AOI211_X1 g035(.A(G131), .B(new_n219), .C1(new_n208), .C2(new_n215), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n201), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n207), .A2(KEYINPUT66), .A3(KEYINPUT11), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n213), .B1(new_n212), .B2(new_n214), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n220), .B(new_n202), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n209), .A2(G134), .ZN(new_n227));
  OAI21_X1  g041(.A(G131), .B1(new_n207), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT68), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G128), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n188), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n231), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n196), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n193), .A2(new_n240), .A3(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n226), .A2(new_n228), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n223), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G119), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  INV_X1    g061(.A(G119), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G116), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n245), .A2(KEYINPUT70), .A3(G119), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT2), .B(G113), .Z(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n244), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n255));
  INV_X1    g069(.A(new_n242), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n226), .A2(new_n228), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(KEYINPUT72), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n226), .A2(new_n259), .A3(new_n228), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n220), .B1(new_n224), .B2(new_n225), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n226), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n201), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n195), .A2(KEYINPUT71), .A3(new_n200), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n258), .A2(new_n260), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n253), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n255), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n260), .A3(new_n242), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n263), .A2(new_n267), .ZN(new_n273));
  AND4_X1   g087(.A1(new_n255), .A2(new_n272), .A3(new_n269), .A4(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n254), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G237), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G210), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(KEYINPUT27), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G101), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n281), .B(KEYINPUT73), .Z(new_n282));
  NOR3_X1   g096(.A1(new_n275), .A2(KEYINPUT29), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n272), .A2(new_n273), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n253), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n270), .B2(new_n274), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT29), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n281), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n268), .A2(new_n269), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT30), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n195), .A2(new_n200), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n262), .B2(new_n226), .ZN(new_n293));
  INV_X1    g107(.A(new_n243), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n244), .A2(new_n297), .A3(new_n291), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n296), .A2(new_n298), .B1(KEYINPUT30), .B2(new_n268), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n290), .B1(new_n299), .B2(new_n253), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n283), .B1(new_n288), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G472), .B1(new_n303), .B2(G902), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n272), .A2(KEYINPUT30), .A3(new_n273), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n297), .B1(new_n244), .B2(new_n291), .ZN(new_n306));
  AOI211_X1 g120(.A(KEYINPUT69), .B(KEYINPUT30), .C1(new_n223), .C2(new_n243), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n253), .B(new_n305), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n281), .A3(new_n289), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT31), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n275), .A2(new_n282), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT31), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n308), .A2(new_n312), .A3(new_n281), .A4(new_n289), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT32), .ZN(new_n315));
  NOR2_X1   g129(.A1(G472), .A2(G902), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n304), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G122), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G116), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT92), .ZN(new_n322));
  INV_X1    g136(.A(G107), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n245), .A2(G122), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n325), .A2(KEYINPUT94), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(KEYINPUT94), .ZN(new_n327));
  INV_X1    g141(.A(new_n322), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n324), .B(KEYINPUT14), .ZN(new_n329));
  OAI21_X1  g143(.A(G107), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT68), .B(G128), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G143), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n333), .A2(KEYINPUT93), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(KEYINPUT93), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n218), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n189), .A2(G128), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n337), .B1(new_n336), .B2(new_n338), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n326), .B(new_n331), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(new_n324), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G107), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n325), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n338), .B(KEYINPUT13), .Z(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n334), .B2(new_n335), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n342), .B(new_n345), .C1(new_n204), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT9), .B(G234), .ZN(new_n350));
  INV_X1    g164(.A(G217), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n350), .A2(new_n351), .A3(G953), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n348), .A3(new_n352), .ZN(new_n355));
  AOI21_X1  g169(.A(G902), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G478), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n357), .A2(KEYINPUT15), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n356), .B(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G902), .ZN(new_n360));
  INV_X1    g174(.A(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G125), .ZN(new_n362));
  INV_X1    g176(.A(G125), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G140), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n362), .A2(new_n364), .A3(KEYINPUT75), .A4(KEYINPUT16), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n362), .A2(new_n364), .A3(KEYINPUT16), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT16), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n361), .A3(G125), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT75), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n187), .B(new_n365), .C1(new_n366), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n362), .A2(new_n364), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n369), .B(new_n368), .C1(new_n373), .C2(new_n367), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n187), .B1(new_n374), .B2(new_n365), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n276), .A2(new_n277), .A3(G214), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(G143), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT17), .A3(G131), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n378), .B(new_n202), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n376), .B(new_n380), .C1(new_n381), .C2(KEYINPUT17), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(KEYINPUT18), .A3(G131), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n373), .B(G146), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT18), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n378), .B1(new_n385), .B2(new_n202), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT91), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n382), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n390), .B1(new_n382), .B2(new_n387), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n360), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G475), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n365), .B1(new_n366), .B2(new_n370), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G146), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n373), .B1(new_n399), .B2(KEYINPUT19), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n373), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n381), .B(new_n398), .C1(G146), .C2(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n403), .A2(new_n387), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n392), .B1(new_n404), .B2(new_n390), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT20), .ZN(new_n406));
  NOR2_X1   g220(.A1(G475), .A2(G902), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n396), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G952), .ZN(new_n412));
  AOI211_X1 g226(.A(G953), .B(new_n412), .C1(G234), .C2(G237), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(G898), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G234), .ZN(new_n417));
  OAI211_X1 g231(.A(G902), .B(G953), .C1(new_n417), .C2(new_n276), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n419), .B(KEYINPUT95), .Z(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n359), .A2(new_n411), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G214), .B1(G237), .B2(G902), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n239), .A2(new_n363), .A3(new_n241), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n201), .A2(new_n363), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT86), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G224), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(G953), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n292), .A2(G125), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n426), .A2(KEYINPUT7), .A3(new_n429), .A4(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n430), .B1(G125), .B2(new_n242), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n429), .A2(KEYINPUT7), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT8), .ZN(new_n438));
  INV_X1    g252(.A(G101), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n323), .A2(G104), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n389), .A2(G107), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n389), .A2(KEYINPUT3), .A3(G107), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n323), .A2(G104), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT3), .B1(new_n389), .B2(G107), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n445), .A2(KEYINPUT82), .A3(new_n439), .A4(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT3), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n323), .A3(G104), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n446), .A2(new_n449), .A3(new_n439), .A4(new_n441), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n442), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n454));
  INV_X1    g268(.A(G113), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT5), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n246), .B2(new_n456), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n454), .A2(new_n457), .B1(new_n251), .B2(new_n252), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n453), .A2(new_n458), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n438), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n433), .A2(KEYINPUT88), .A3(new_n436), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n446), .A2(new_n449), .A3(new_n441), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT81), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT4), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n446), .A2(new_n449), .A3(KEYINPUT81), .A4(new_n441), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(new_n467), .A3(G101), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n253), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n447), .A2(new_n452), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(G101), .A3(new_n468), .ZN(new_n474));
  AND4_X1   g288(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT4), .A4(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n467), .B1(new_n447), .B2(new_n452), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(new_n476), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n471), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n437), .A3(new_n459), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n463), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n453), .B(new_n458), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n481), .A2(new_n438), .B1(new_n434), .B2(new_n435), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT88), .B1(new_n482), .B2(new_n433), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n360), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n437), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n473), .A2(KEYINPUT4), .A3(new_n474), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n476), .A2(new_n472), .A3(new_n474), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n470), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n485), .B1(new_n489), .B2(new_n460), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(KEYINPUT6), .A3(new_n479), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n426), .A2(new_n432), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n428), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n494), .B(new_n485), .C1(new_n489), .C2(new_n460), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT87), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT87), .A4(new_n495), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n484), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT89), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n501), .ZN(new_n505));
  AOI211_X1 g319(.A(new_n505), .B(new_n484), .C1(new_n498), .C2(new_n499), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n422), .B(new_n423), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT23), .B1(new_n232), .B2(G119), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n232), .A2(G119), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT23), .A4(G119), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR3_X1    g327(.A1(new_n513), .A2(KEYINPUT77), .A3(G110), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n510), .B1(new_n332), .B2(G119), .ZN(new_n515));
  XOR2_X1   g329(.A(KEYINPUT24), .B(G110), .Z(new_n516));
  OR3_X1    g330(.A1(new_n515), .A2(KEYINPUT78), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT77), .B1(new_n513), .B2(G110), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT78), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n514), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n373), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n375), .B1(new_n187), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n515), .A2(new_n516), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n372), .B2(new_n375), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT74), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n513), .B2(G110), .ZN(new_n527));
  INV_X1    g341(.A(G110), .ZN(new_n528));
  AOI211_X1 g342(.A(KEYINPUT74), .B(new_n528), .C1(new_n511), .C2(new_n512), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT76), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n525), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n398), .A2(new_n371), .B1(new_n515), .B2(new_n516), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n528), .B1(new_n511), .B2(new_n512), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(new_n526), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT76), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n523), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT22), .B(G137), .ZN(new_n538));
  INV_X1    g352(.A(G221), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n539), .A2(new_n417), .A3(G953), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n538), .B(new_n540), .Z(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n523), .B(new_n541), .C1(new_n532), .C2(new_n536), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n360), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT79), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n351), .B1(G234), .B2(new_n360), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n545), .A2(new_n547), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n543), .A2(KEYINPUT25), .A3(new_n360), .A4(new_n544), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(KEYINPUT79), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n549), .A2(G902), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n554), .B(KEYINPUT80), .Z(new_n555));
  NAND2_X1  g369(.A1(new_n543), .A2(new_n544), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n550), .A2(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G469), .ZN(new_n559));
  INV_X1    g373(.A(new_n442), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n232), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n241), .B1(new_n193), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n450), .A2(new_n451), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n450), .A2(new_n451), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n560), .B(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n242), .B2(new_n453), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n263), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n263), .A2(new_n566), .A3(KEYINPUT12), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(KEYINPUT84), .A3(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n265), .A2(new_n266), .A3(new_n469), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n475), .B2(new_n477), .ZN(new_n573));
  INV_X1    g387(.A(new_n263), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n453), .A2(new_n242), .A3(KEYINPUT10), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT84), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n567), .A2(new_n580), .A3(new_n568), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G110), .B(G140), .ZN(new_n583));
  INV_X1    g397(.A(G227), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G953), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n583), .B(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n265), .A2(new_n266), .A3(new_n469), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n487), .B2(new_n488), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n576), .A2(new_n577), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n263), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n587), .B1(new_n591), .B2(new_n579), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT85), .ZN(new_n593));
  OAI22_X1  g407(.A1(new_n582), .A2(new_n586), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n559), .B(new_n360), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n559), .A2(new_n360), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n579), .A2(new_n581), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n570), .A2(KEYINPUT84), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT12), .B1(new_n263), .B2(new_n566), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n586), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n591), .A2(new_n579), .A3(new_n587), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n596), .B(new_n598), .C1(new_n605), .C2(new_n559), .ZN(new_n606));
  INV_X1    g420(.A(new_n350), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n539), .B1(new_n607), .B2(new_n360), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n319), .A2(new_n508), .A3(new_n558), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  AND3_X1   g426(.A1(new_n606), .A2(new_n558), .A3(new_n609), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n312), .B1(new_n300), .B2(new_n281), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n311), .A2(new_n313), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n316), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n314), .B2(new_n360), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n410), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n622), .A2(new_n408), .B1(G475), .B2(new_n395), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n349), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n354), .A2(new_n625), .A3(KEYINPUT33), .A4(new_n355), .ZN(new_n626));
  INV_X1    g440(.A(new_n355), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n352), .B1(new_n341), .B2(new_n348), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT96), .B1(new_n341), .B2(new_n348), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  OAI22_X1  g444(.A1(new_n627), .A2(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n357), .B1(new_n626), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n357), .A2(new_n360), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n360), .B1(new_n627), .B2(new_n628), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(G478), .ZN(new_n636));
  NOR4_X1   g450(.A1(new_n623), .A2(new_n632), .A3(new_n636), .A4(new_n421), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n498), .A2(new_n499), .ZN(new_n638));
  INV_X1    g452(.A(new_n484), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n501), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n637), .B(new_n423), .C1(new_n506), .C2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n621), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G104), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NAND2_X1  g460(.A1(new_n359), .A2(new_n623), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n421), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n648), .B(new_n423), .C1(new_n506), .C2(new_n640), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n621), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NAND2_X1  g467(.A1(new_n550), .A2(new_n553), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n537), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n537), .A2(new_n656), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n658), .A2(new_n555), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT98), .B1(new_n654), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n663));
  AOI211_X1 g477(.A(new_n663), .B(new_n660), .C1(new_n550), .C2(new_n553), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n508), .A2(new_n620), .A3(new_n665), .A4(new_n610), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  OAI21_X1  g482(.A(new_n423), .B1(new_n640), .B2(new_n506), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n669), .A2(new_n662), .A3(new_n664), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n414), .B1(new_n418), .B2(G900), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT99), .Z(new_n672));
  NOR2_X1   g486(.A1(new_n647), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n670), .A2(new_n319), .A3(new_n610), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  NOR2_X1   g489(.A1(new_n504), .A2(new_n506), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT38), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n285), .A2(new_n289), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n618), .B1(new_n679), .B2(new_n282), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n309), .A2(new_n680), .B1(G472), .B2(G902), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n683), .B1(new_n317), .B2(new_n318), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n654), .A2(new_n661), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n359), .A2(new_n411), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n686), .A2(new_n687), .A3(new_n423), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n678), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n672), .B(KEYINPUT39), .Z(new_n690));
  NAND2_X1  g504(.A1(new_n610), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT40), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n189), .ZN(G45));
  NOR2_X1   g508(.A1(new_n632), .A2(new_n636), .ZN(new_n695));
  INV_X1    g509(.A(new_n672), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n411), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n670), .A2(new_n319), .A3(new_n610), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  OAI21_X1  g514(.A(new_n360), .B1(new_n594), .B2(new_n595), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n609), .A3(new_n596), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n642), .A2(new_n319), .A3(new_n558), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND4_X1  g521(.A1(new_n650), .A2(new_n319), .A3(new_n558), .A4(new_n704), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NOR2_X1   g523(.A1(new_n669), .A2(new_n703), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n319), .A2(new_n710), .A3(new_n422), .A4(new_n665), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  INV_X1    g526(.A(new_n313), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n309), .A2(KEYINPUT31), .B1(new_n282), .B2(new_n286), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n713), .B1(new_n714), .B2(KEYINPUT102), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n286), .A2(new_n282), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n716), .B1(new_n614), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n316), .B(KEYINPUT101), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n619), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n687), .B(new_n423), .C1(new_n640), .C2(new_n506), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n703), .A2(new_n421), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n721), .A2(new_n723), .A3(new_n558), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NAND4_X1  g540(.A1(new_n721), .A2(new_n710), .A3(new_n685), .A4(new_n698), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  NAND2_X1  g542(.A1(new_n604), .A2(KEYINPUT103), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n591), .A2(new_n579), .A3(new_n730), .A4(new_n587), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n603), .A2(new_n729), .A3(G469), .A4(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n596), .A2(new_n598), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT105), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n604), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n737), .A2(new_n730), .B1(new_n582), .B2(new_n586), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n733), .A3(G469), .A4(new_n729), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n732), .A2(KEYINPUT104), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n596), .A4(new_n598), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n500), .A2(new_n503), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n638), .A2(new_n501), .A3(new_n639), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n746), .A3(new_n423), .A4(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n747), .B(new_n423), .C1(new_n503), .C2(new_n500), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n609), .A2(new_n744), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n558), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n616), .A2(KEYINPUT32), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n752), .B1(new_n755), .B2(new_n304), .ZN(new_n756));
  NOR2_X1   g570(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n751), .A2(new_n756), .A3(new_n698), .A4(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n750), .A2(new_n748), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n608), .B1(new_n736), .B2(new_n743), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n756), .A3(new_n698), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n757), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND4_X1  g579(.A1(new_n760), .A2(new_n756), .A3(new_n673), .A4(new_n761), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  OR2_X1    g581(.A1(new_n617), .A2(new_n619), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n411), .A2(new_n632), .A3(new_n636), .A4(KEYINPUT43), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n623), .A2(KEYINPUT108), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n411), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n695), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n769), .B1(new_n773), .B2(KEYINPUT43), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n768), .A2(new_n685), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT109), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n774), .A2(new_n685), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n779), .A3(KEYINPUT44), .A4(new_n768), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n750), .A2(new_n748), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n775), .B2(new_n776), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n738), .A2(KEYINPUT45), .A3(new_n729), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n559), .B1(new_n605), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n598), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n596), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n609), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n690), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n781), .A2(KEYINPUT110), .A3(new_n783), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n786), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT111), .B(G137), .Z(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(G39));
  NOR2_X1   g617(.A1(new_n697), .A2(new_n558), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n760), .A2(new_n755), .A3(new_n304), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n797), .A2(KEYINPUT47), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n796), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n361), .ZN(G42));
  INV_X1    g624(.A(new_n423), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n773), .A2(new_n608), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n702), .A2(new_n596), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n558), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT112), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n817));
  OR4_X1    g631(.A1(new_n678), .A2(new_n816), .A3(new_n684), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n760), .A2(new_n413), .A3(new_n704), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n752), .A3(new_n684), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n820), .B(new_n623), .C1(new_n632), .C2(new_n636), .ZN(new_n821));
  INV_X1    g635(.A(new_n774), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n685), .A3(new_n721), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n677), .A2(new_n811), .A3(new_n704), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n721), .A2(new_n558), .A3(new_n413), .A4(new_n774), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(KEYINPUT50), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n827), .A2(KEYINPUT50), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n821), .B(new_n824), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n806), .B(new_n808), .C1(new_n609), .C2(new_n813), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n826), .A2(new_n782), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n832), .B2(new_n833), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n831), .B(KEYINPUT51), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n838));
  AND2_X1   g652(.A1(new_n832), .A2(new_n835), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n830), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n710), .ZN(new_n841));
  OAI211_X1 g655(.A(G952), .B(new_n277), .C1(new_n826), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n695), .A2(new_n411), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n820), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT120), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n823), .A2(new_n756), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT48), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n837), .A2(new_n840), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n676), .A2(new_n811), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n613), .A3(new_n620), .A4(new_n648), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n611), .A2(new_n666), .A3(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n637), .B(new_n423), .C1(new_n504), .C2(new_n506), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n745), .A2(new_n747), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT113), .A3(new_n423), .A4(new_n637), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n856), .A2(new_n858), .A3(new_n620), .A4(new_n613), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n606), .A2(new_n609), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n755), .B2(new_n304), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n359), .A2(new_n411), .A3(new_n672), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n760), .A2(new_n861), .A3(new_n665), .A4(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n853), .A2(new_n766), .A3(new_n859), .A4(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n744), .A2(new_n609), .A3(new_n748), .A4(new_n750), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n721), .A2(new_n685), .A3(new_n698), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT114), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n720), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n715), .B2(new_n718), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n869), .A2(new_n686), .A3(new_n619), .A4(new_n697), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n760), .A3(new_n871), .A4(new_n761), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n685), .A2(new_n608), .A3(new_n672), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n744), .A2(new_n684), .A3(new_n723), .A4(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n674), .A2(new_n699), .A3(new_n727), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n861), .B(new_n670), .C1(new_n673), .C2(new_n698), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .A3(new_n727), .A4(new_n877), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n875), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n708), .A2(new_n705), .A3(new_n711), .A4(new_n725), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n759), .B2(new_n763), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n874), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n880), .A2(new_n882), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n867), .A2(new_n872), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n766), .A2(new_n863), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n859), .A2(new_n611), .A3(new_n666), .A4(new_n852), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n888), .A2(new_n885), .A3(new_n889), .A4(new_n892), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n886), .A2(new_n887), .B1(new_n893), .B2(new_n875), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n874), .A2(new_n883), .A3(KEYINPUT115), .A4(new_n885), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n850), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n875), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n864), .B2(new_n873), .ZN(new_n899));
  INV_X1    g713(.A(new_n890), .ZN(new_n900));
  INV_X1    g714(.A(new_n891), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT116), .A4(new_n889), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n899), .A2(new_n885), .A3(new_n883), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n897), .A2(new_n903), .A3(new_n850), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT117), .B1(new_n896), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n888), .A2(new_n885), .A3(KEYINPUT53), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n892), .A2(new_n889), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n887), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n895), .A3(new_n897), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n912), .A3(new_n904), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n849), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(G952), .A2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n818), .B1(new_n914), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n277), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n360), .B1(new_n897), .B2(new_n903), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n491), .A2(new_n495), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n493), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n918), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT56), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n897), .A2(new_n903), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(G902), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n925), .B(new_n923), .C1(new_n927), .C2(new_n503), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(G51));
  XNOR2_X1  g746(.A(new_n926), .B(new_n850), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n597), .B(KEYINPUT57), .Z(new_n934));
  OAI22_X1  g748(.A1(new_n933), .A2(new_n934), .B1(new_n595), .B2(new_n594), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n919), .A2(new_n787), .A3(new_n789), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n917), .B1(new_n935), .B2(new_n936), .ZN(G54));
  AND3_X1   g751(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n918), .B1(new_n938), .B2(new_n405), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n405), .B2(new_n938), .ZN(G60));
  XOR2_X1   g754(.A(new_n633), .B(KEYINPUT59), .Z(new_n941));
  NAND3_X1  g755(.A1(new_n626), .A2(new_n631), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n918), .B1(new_n933), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n906), .A2(new_n913), .A3(new_n941), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n626), .A2(new_n631), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(G63));
  NAND2_X1  g760(.A1(new_n658), .A2(new_n659), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n926), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n897), .B2(new_n903), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n952), .B(new_n918), .C1(new_n557), .C2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT61), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT61), .B1(new_n954), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  OAI21_X1  g772(.A(G953), .B1(new_n415), .B2(new_n427), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT123), .Z(new_n960));
  NOR2_X1   g774(.A1(new_n891), .A2(new_n884), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n921), .B1(G898), .B2(new_n277), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  XOR2_X1   g778(.A(new_n299), .B(KEYINPUT124), .Z(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(new_n402), .Z(new_n966));
  INV_X1    g780(.A(new_n756), .ZN(new_n967));
  AOI211_X1 g781(.A(new_n691), .B(new_n967), .C1(new_n843), .C2(new_n647), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n809), .B1(new_n760), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n881), .A2(new_n727), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n971), .B(new_n972), .C1(new_n689), .C2(new_n692), .ZN(new_n973));
  OAI21_X1  g787(.A(KEYINPUT62), .B1(new_n693), .B2(new_n970), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n969), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n801), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n966), .B1(new_n977), .B2(G953), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n756), .A2(new_n723), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n766), .B1(new_n798), .B2(new_n979), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n980), .A2(new_n809), .A3(new_n970), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n801), .A2(new_n981), .A3(new_n277), .A4(new_n764), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n966), .B1(G900), .B2(G953), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(G900), .ZN(new_n986));
  OAI21_X1  g800(.A(G953), .B1(new_n584), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n985), .B(new_n987), .ZN(G72));
  INV_X1    g802(.A(new_n300), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n989), .A2(new_n281), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n801), .A2(new_n981), .A3(new_n764), .A4(new_n961), .ZN(new_n991));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT125), .Z(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n995), .A2(new_n917), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n989), .A2(new_n281), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n910), .A2(new_n997), .A3(new_n990), .A4(new_n993), .ZN(new_n998));
  INV_X1    g812(.A(new_n994), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n977), .B2(new_n961), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n996), .B(new_n998), .C1(new_n997), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(KEYINPUT126), .ZN(new_n1002));
  INV_X1    g816(.A(new_n997), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n977), .A2(new_n961), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n999), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1005), .A2(new_n1006), .A3(new_n998), .A4(new_n996), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1002), .A2(new_n1007), .ZN(G57));
endmodule


