//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT68), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT69), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  OR4_X1    g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n458), .B1(new_n465), .B2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AOI211_X1 g042(.A(KEYINPUT70), .B(new_n467), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n460), .A2(new_n462), .A3(G137), .A4(new_n467), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n459), .A2(G2105), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G101), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  NOR4_X1   g049(.A1(new_n474), .A2(new_n459), .A3(KEYINPUT71), .A4(G2105), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n469), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n460), .A2(new_n462), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n467), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(G2105), .ZN(new_n481));
  AOI22_X1  g056(.A1(G124), .A2(new_n480), .B1(new_n481), .B2(G136), .ZN(new_n482));
  NOR3_X1   g057(.A1(KEYINPUT72), .A2(G100), .A3(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT72), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT73), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n467), .ZN(new_n491));
  OAI211_X1 g066(.A(KEYINPUT75), .B(new_n490), .C1(new_n491), .C2(KEYINPUT76), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT74), .B1(new_n467), .B2(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n460), .A2(new_n462), .A3(G126), .A4(G2105), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT75), .ZN(new_n502));
  AND4_X1   g077(.A1(G138), .A2(new_n460), .A3(new_n462), .A4(new_n467), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n491), .B2(KEYINPUT75), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n492), .B(new_n501), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n516), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XOR2_X1   g100(.A(new_n525), .B(KEYINPUT7), .Z(new_n526));
  INV_X1    g101(.A(new_n518), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n520), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n533));
  INV_X1    g108(.A(new_n520), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n535), .B2(new_n529), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n528), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n515), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n518), .A2(new_n541), .B1(new_n520), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n515), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n518), .A2(new_n547), .B1(new_n520), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT78), .B1(new_n546), .B2(new_n549), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT79), .Z(G188));
  NAND2_X1  g136(.A1(new_n527), .A2(G91), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT80), .B(G65), .Z(new_n563));
  AOI22_X1  g138(.A1(new_n513), .A2(new_n563), .B1(G78), .B2(G543), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n534), .B2(G53), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  NOR3_X1   g142(.A1(new_n520), .A2(KEYINPUT9), .A3(new_n567), .ZN(new_n568));
  OAI221_X1 g143(.A(new_n562), .B1(new_n515), .B2(new_n564), .C1(new_n566), .C2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  XNOR2_X1  g145(.A(new_n531), .B(KEYINPUT77), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT81), .B1(new_n571), .B2(new_n528), .ZN(new_n572));
  OAI211_X1 g147(.A(KEYINPUT81), .B(new_n528), .C1(new_n532), .C2(new_n536), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G286));
  NAND2_X1  g151(.A1(new_n527), .A2(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n534), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT82), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n527), .A2(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n510), .A2(new_n512), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n585), .A2(new_n590), .A3(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n515), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n518), .A2(new_n595), .B1(new_n520), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n527), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n518), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n601), .A2(new_n604), .B1(G54), .B2(new_n534), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n587), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n515), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(new_n608), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G321));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(G299), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n575), .B2(new_n616), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(new_n575), .B2(new_n616), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  INV_X1    g196(.A(new_n554), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n616), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n612), .A2(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n616), .B2(new_n624), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g201(.A(new_n479), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n472), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT84), .B(G2100), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n629), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n480), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n481), .A2(G135), .ZN(new_n634));
  OR2_X1    g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n635), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G2096), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n632), .A2(new_n639), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT16), .B(G1341), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(G14), .B1(new_n646), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n646), .A2(new_n652), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT17), .ZN(new_n657));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT85), .ZN(new_n661));
  INV_X1    g236(.A(new_n659), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n662), .A2(new_n656), .A3(new_n658), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n659), .B1(new_n656), .B2(new_n658), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n657), .B2(new_n658), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT88), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n672), .A2(new_n673), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT20), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n675), .A2(new_n677), .A3(new_n680), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n687), .B(new_n690), .Z(G229));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G22), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(G1971), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(G6), .ZN(new_n697));
  INV_X1    g272(.A(G305), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n692), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G16), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(new_n580), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n696), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT90), .B(G29), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n480), .A2(G119), .ZN(new_n715));
  OR2_X1    g290(.A1(G95), .A2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT91), .Z(new_n718));
  AOI211_X1 g293(.A(new_n715), .B(new_n718), .C1(G131), .C2(new_n481), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n714), .B1(new_n719), .B2(new_n713), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT35), .B(G1991), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT92), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n692), .A2(G24), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n598), .B2(new_n692), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1986), .Z(new_n726));
  NAND4_X1  g301(.A1(new_n710), .A2(new_n711), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT36), .Z(new_n728));
  AOI22_X1  g303(.A1(G129), .A2(new_n480), .B1(new_n481), .B2(G141), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT26), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G105), .B2(new_n472), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  MUX2_X1   g308(.A(G32), .B(new_n733), .S(G29), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT100), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT27), .B(G1996), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n713), .A2(G26), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  INV_X1    g314(.A(new_n481), .ZN(new_n740));
  INV_X1    g315(.A(G140), .ZN(new_n741));
  OR3_X1    g316(.A1(new_n740), .A2(KEYINPUT95), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(KEYINPUT95), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n480), .A2(G128), .ZN(new_n744));
  OR2_X1    g319(.A1(G104), .A2(G2105), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n745), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n746));
  AND4_X1   g321(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n739), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G2067), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n692), .A2(G5), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G171), .B2(new_n692), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT102), .ZN(new_n754));
  INV_X1    g329(.A(G1961), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n737), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n748), .A2(G33), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n481), .A2(G139), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n472), .A2(G103), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT96), .B(KEYINPUT25), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n759), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n627), .A2(G127), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n467), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT97), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n758), .B1(new_n770), .B2(new_n748), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n771), .A2(G2072), .B1(new_n755), .B2(new_n754), .ZN(new_n772));
  NAND2_X1  g347(.A1(G168), .A2(G16), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G16), .B2(G21), .ZN(new_n774));
  INV_X1    g349(.A(G1966), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n772), .B(new_n776), .C1(G2072), .C2(new_n771), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n637), .A2(new_n713), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT101), .B(KEYINPUT31), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G11), .ZN(new_n780));
  OR2_X1    g355(.A1(KEYINPUT30), .A2(G28), .ZN(new_n781));
  NAND2_X1  g356(.A1(KEYINPUT30), .A2(G28), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n778), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n713), .A2(G27), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n713), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n784), .B1(G2078), .B2(new_n786), .C1(new_n774), .C2(new_n775), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n613), .A2(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G4), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT24), .B(G34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n713), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT98), .Z(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n477), .B2(new_n748), .ZN(new_n794));
  INV_X1    g369(.A(G2084), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n789), .A2(new_n790), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n790), .B2(new_n789), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n757), .A2(new_n777), .A3(new_n787), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT99), .B1(new_n794), .B2(new_n795), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT23), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n692), .A2(G20), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n800), .B(new_n801), .C1(G299), .C2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n800), .B2(new_n801), .ZN(new_n803));
  INV_X1    g378(.A(G1956), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n794), .A2(KEYINPUT99), .A3(new_n795), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G2078), .B2(new_n786), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n798), .A2(new_n799), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n713), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n713), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT29), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G2090), .Z(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G19), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n554), .B2(G16), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT94), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1341), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT103), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(KEYINPUT103), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n728), .B1(new_n819), .B2(new_n820), .ZN(G311));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  INV_X1    g397(.A(new_n728), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(G150));
  AOI22_X1  g399(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n515), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  INV_X1    g402(.A(G55), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n518), .A2(new_n827), .B1(new_n520), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n552), .B2(new_n553), .ZN(new_n831));
  INV_X1    g406(.A(new_n830), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(new_n550), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n612), .A2(new_n620), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n832), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XOR2_X1   g419(.A(new_n719), .B(new_n629), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n488), .B(G160), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n637), .ZN(new_n847));
  INV_X1    g422(.A(new_n480), .ZN(new_n848));
  INV_X1    g423(.A(G130), .ZN(new_n849));
  OR3_X1    g424(.A1(new_n848), .A2(KEYINPUT105), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT105), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n481), .A2(G142), .ZN(new_n852));
  OR2_X1    g427(.A1(G106), .A2(G2105), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n847), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n847), .A2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n845), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  INV_X1    g436(.A(new_n845), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n857), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n507), .B(new_n733), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n747), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(new_n768), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n770), .B2(new_n866), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n860), .A2(new_n863), .A3(new_n868), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g449(.A1(new_n832), .A2(new_n616), .ZN(new_n875));
  XNOR2_X1  g450(.A(G303), .B(new_n580), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n598), .B(KEYINPUT106), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n698), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n878), .A2(new_n698), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n878), .A2(new_n698), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n876), .A3(new_n879), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT42), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT108), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n882), .A2(KEYINPUT107), .A3(new_n884), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT107), .B1(new_n882), .B2(new_n884), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT42), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n612), .B(G299), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n613), .A2(G299), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n613), .A2(G299), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n834), .B(new_n624), .ZN(new_n900));
  MUX2_X1   g475(.A(new_n893), .B(new_n899), .S(new_n900), .Z(new_n901));
  XNOR2_X1  g476(.A(new_n891), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n875), .B1(new_n902), .B2(new_n616), .ZN(G295));
  OAI21_X1  g478(.A(new_n875), .B1(new_n902), .B2(new_n616), .ZN(G331));
  INV_X1    g479(.A(KEYINPUT111), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT81), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n537), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G301), .B1(new_n908), .B2(new_n573), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n537), .A2(G171), .ZN(new_n910));
  OAI22_X1  g485(.A1(new_n909), .A2(new_n910), .B1(new_n831), .B2(new_n833), .ZN(new_n911));
  OAI21_X1  g486(.A(G171), .B1(new_n572), .B2(new_n574), .ZN(new_n912));
  INV_X1    g487(.A(new_n910), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n834), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n906), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(new_n834), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT109), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n905), .B1(new_n919), .B2(new_n893), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n911), .A2(new_n914), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n899), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT110), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n899), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR4_X1   g501(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT111), .A4(new_n892), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n920), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(new_n889), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n899), .B1(new_n915), .B2(new_n918), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n911), .A2(new_n914), .A3(new_n893), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n889), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n872), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n889), .B1(new_n930), .B2(new_n931), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n934), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n932), .A2(new_n872), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n938), .B(new_n939), .C1(new_n928), .C2(new_n889), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n933), .B2(new_n935), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT112), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n945), .B(KEYINPUT44), .C1(new_n940), .C2(new_n941), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n937), .B1(new_n944), .B2(new_n946), .ZN(G397));
  INV_X1    g522(.A(new_n469), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n501), .A2(new_n492), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT75), .B1(new_n491), .B2(KEYINPUT76), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n950), .B(KEYINPUT4), .C1(KEYINPUT75), .C2(new_n491), .ZN(new_n951));
  AOI21_X1  g526(.A(G1384), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n948), .B1(new_n952), .B2(KEYINPUT45), .ZN(new_n953));
  OAI211_X1 g528(.A(G40), .B(new_n470), .C1(new_n473), .C2(new_n475), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n503), .A2(new_n504), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n506), .B1(new_n956), .B2(KEYINPUT75), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n501), .A2(new_n492), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n954), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G2078), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n953), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(KEYINPUT50), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n466), .A2(new_n468), .A3(new_n954), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n507), .A2(new_n967), .A3(new_n955), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n963), .A2(new_n964), .B1(new_n755), .B2(new_n969), .ZN(new_n970));
  AOI211_X1 g545(.A(new_n964), .B(G2078), .C1(new_n465), .C2(G2105), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n961), .B(new_n971), .C1(new_n960), .C2(new_n959), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(G171), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n953), .A2(new_n961), .A3(KEYINPUT53), .A4(new_n962), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(G301), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n977), .A2(KEYINPUT54), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT126), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n973), .A2(new_n979), .A3(G171), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n973), .A2(G171), .ZN(new_n983));
  AOI21_X1  g558(.A(G301), .B1(new_n970), .B2(new_n976), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n969), .A2(G2090), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n953), .A2(new_n961), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n695), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(G303), .A2(G8), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(KEYINPUT115), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n989), .A2(new_n998), .A3(G8), .ZN(new_n999));
  XOR2_X1   g574(.A(KEYINPUT117), .B(KEYINPUT49), .Z(new_n1000));
  INV_X1    g575(.A(new_n590), .ZN(new_n1001));
  INV_X1    g576(.A(G86), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n591), .B1(new_n518), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(G1981), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n585), .A2(new_n1005), .A3(new_n590), .A4(new_n591), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1000), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(KEYINPUT118), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n952), .B2(new_n966), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(KEYINPUT118), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1004), .A2(new_n1006), .A3(KEYINPUT49), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT116), .B(G1976), .Z(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n703), .A2(G1976), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n966), .A2(new_n955), .A3(new_n507), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(G8), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT52), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1013), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n999), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1009), .B1(new_n986), .B2(new_n988), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(new_n994), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n987), .A2(new_n775), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n507), .A2(new_n967), .A3(new_n955), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n967), .B1(new_n507), .B2(new_n955), .ZN(new_n1029));
  OR3_X1    g604(.A1(new_n466), .A2(new_n468), .A3(new_n954), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n795), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1009), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n537), .A2(G8), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1026), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n969), .A2(G2084), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1966), .B1(new_n953), .B2(new_n961), .ZN(new_n1038));
  OAI21_X1  g613(.A(G8), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(KEYINPUT51), .A3(new_n1034), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT125), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(new_n1035), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT125), .B(new_n1034), .C1(new_n1027), .C2(new_n1032), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1036), .B(new_n1040), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n981), .A2(new_n985), .A3(new_n1025), .A4(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(G299), .B(KEYINPUT57), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n953), .A2(new_n961), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1030), .B1(KEYINPUT50), .B2(new_n959), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1956), .B1(new_n1050), .B2(new_n968), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1047), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  XOR2_X1   g628(.A(G299), .B(KEYINPUT57), .Z(new_n1054));
  NAND2_X1  g629(.A1(new_n969), .A2(new_n804), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n953), .A2(new_n961), .A3(new_n1048), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1052), .A2(new_n1053), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1053), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1061));
  XOR2_X1   g636(.A(new_n1061), .B(KEYINPUT122), .Z(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT58), .B(G1341), .Z(new_n1065));
  AND3_X1   g640(.A1(new_n1018), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1018), .B2(new_n1065), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1996), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n953), .A2(new_n961), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n622), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1063), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1067), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1018), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n554), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1072), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n1062), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1073), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1060), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  AND4_X1   g657(.A1(new_n955), .A2(new_n966), .A3(new_n750), .A4(new_n507), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n969), .B2(new_n790), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1084), .A2(KEYINPUT60), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1083), .ZN(new_n1086));
  OAI211_X1 g661(.A(KEYINPUT60), .B(new_n1086), .C1(new_n1031), .C2(G1348), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n613), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(KEYINPUT60), .A3(new_n612), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1088), .B1(new_n1087), .B2(new_n613), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1082), .B(new_n1085), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n1095), .B(new_n1083), .C1(new_n969), .C2(new_n790), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT123), .B1(new_n1096), .B2(new_n612), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(new_n1090), .A3(new_n1089), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1082), .B1(new_n1098), .B2(new_n1085), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1081), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1052), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1084), .A2(new_n612), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1057), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1046), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1021), .A2(new_n1023), .A3(new_n998), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G288), .A2(G1976), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1013), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1006), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1010), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  OR3_X1    g686(.A1(new_n1039), .A2(KEYINPUT119), .A3(G286), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT119), .B1(new_n1039), .B2(G286), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1025), .A2(KEYINPUT63), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT63), .B1(new_n1025), .B2(new_n1114), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1111), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT127), .B1(new_n1104), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n999), .B(new_n1021), .C1(new_n1023), .C2(new_n994), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1025), .A2(new_n1114), .A3(KEYINPUT63), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1110), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT127), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1103), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1085), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1093), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1129), .B2(new_n1081), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1124), .B(new_n1125), .C1(new_n1130), .C2(new_n1046), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1045), .A2(KEYINPUT62), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1045), .A2(KEYINPUT62), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(new_n984), .A3(new_n1025), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1118), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n952), .A2(KEYINPUT45), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n966), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n719), .B(new_n721), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT114), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n747), .B(G2067), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n733), .B(new_n1069), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1137), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1137), .A2(G1986), .A3(G290), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1137), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(G1986), .A3(G290), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1145), .B1(new_n1151), .B2(KEYINPUT113), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(KEYINPUT113), .B2(new_n1151), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1135), .A2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1146), .A2(KEYINPUT48), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1146), .A2(KEYINPUT48), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1144), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1140), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1148), .B1(new_n1158), .B2(new_n733), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1148), .A2(KEYINPUT46), .A3(new_n1069), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT46), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1137), .B2(G1996), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT47), .Z(new_n1164));
  NAND2_X1  g739(.A1(new_n747), .A2(new_n750), .ZN(new_n1165));
  INV_X1    g740(.A(new_n721), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n719), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1142), .B2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n1157), .B(new_n1164), .C1(new_n1148), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1154), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g745(.A(G319), .B1(new_n653), .B2(new_n654), .ZN(new_n1172));
  NOR3_X1   g746(.A1(G229), .A2(G227), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n873), .A3(new_n1173), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


