//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT70), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT70), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AOI21_X1  g006(.A(G143), .B1(KEYINPUT65), .B2(KEYINPUT85), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n191), .A2(G214), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G214), .ZN(new_n195));
  AOI211_X1 g009(.A(new_n195), .B(G953), .C1(new_n188), .C2(new_n190), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT65), .B(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT85), .ZN(new_n198));
  OAI211_X1 g012(.A(G131), .B(new_n194), .C1(new_n196), .C2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT86), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(G214), .A3(new_n192), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT65), .A2(G143), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT65), .A2(G143), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT85), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(G131), .B1(new_n207), .B2(new_n194), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n200), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n194), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT86), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT87), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n194), .ZN(new_n216));
  AOI21_X1  g030(.A(G953), .B1(new_n188), .B2(new_n190), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n217), .A2(G214), .B1(new_n204), .B2(new_n205), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n212), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT86), .A3(new_n199), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT87), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n213), .ZN(new_n222));
  XNOR2_X1  g036(.A(G125), .B(G140), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT16), .ZN(new_n224));
  INV_X1    g038(.A(G125), .ZN(new_n225));
  OR3_X1    g039(.A1(new_n225), .A2(KEYINPUT16), .A3(G140), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(G146), .A3(new_n226), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n227), .A2(KEYINPUT75), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(KEYINPUT75), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n223), .B(KEYINPUT19), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n215), .A2(new_n222), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n210), .B1(new_n235), .B2(new_n212), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n223), .B(new_n231), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n236), .B(new_n237), .C1(new_n235), .C2(new_n199), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G113), .B(G122), .ZN(new_n240));
  INV_X1    g054(.A(G104), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n224), .A2(new_n226), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n231), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n227), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n207), .A2(KEYINPUT17), .A3(G131), .A4(new_n194), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n249), .A2(KEYINPUT88), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(KEYINPUT88), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT17), .B1(new_n220), .B2(new_n213), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n238), .B(new_n242), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT89), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(new_n255), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n244), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n259));
  NOR2_X1   g073(.A1(G475), .A2(G902), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(new_n255), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT17), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n263), .B1(new_n209), .B2(new_n214), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n249), .A2(KEYINPUT88), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n249), .A2(KEYINPUT88), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n247), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n268), .A2(KEYINPUT89), .A3(new_n238), .A4(new_n242), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n262), .A2(new_n269), .B1(new_n239), .B2(new_n243), .ZN(new_n270));
  INV_X1    g084(.A(new_n260), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT20), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n238), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n243), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n256), .B2(new_n257), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G475), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n192), .A2(G952), .ZN(new_n280));
  INV_X1    g094(.A(G234), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(new_n187), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n282), .B(KEYINPUT93), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(KEYINPUT73), .B(G902), .Z(new_n285));
  AOI211_X1 g099(.A(new_n192), .B(new_n285), .C1(G234), .C2(G237), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT21), .B(G898), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT91), .ZN(new_n290));
  XNOR2_X1  g104(.A(G116), .B(G122), .ZN(new_n291));
  INV_X1    g105(.A(G107), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT14), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G122), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(G116), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n292), .B1(new_n297), .B2(KEYINPUT14), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n290), .A2(new_n293), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n291), .A2(KEYINPUT91), .A3(new_n292), .ZN(new_n300));
  INV_X1    g114(.A(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G143), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n197), .B2(new_n301), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(G134), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n204), .A2(G128), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(new_n302), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n299), .B(new_n300), .C1(new_n304), .C2(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n296), .A2(G116), .ZN(new_n309));
  OAI21_X1  g123(.A(G107), .B1(new_n309), .B2(new_n297), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n293), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(KEYINPUT90), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT13), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n303), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G134), .B1(new_n306), .B2(KEYINPUT13), .ZN(new_n315));
  OAI22_X1  g129(.A1(new_n314), .A2(new_n315), .B1(G134), .B2(new_n303), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n308), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT9), .B(G234), .ZN(new_n318));
  INV_X1    g132(.A(G217), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n318), .A2(new_n319), .A3(G953), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n308), .B(new_n320), .C1(new_n312), .C2(new_n316), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(KEYINPUT92), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT92), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n317), .A2(new_n325), .A3(new_n321), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n285), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G478), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT15), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n327), .B(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n273), .A2(new_n279), .A3(new_n289), .A4(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n319), .B1(new_n285), .B2(G234), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n337));
  INV_X1    g151(.A(G110), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n301), .A2(G119), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G128), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n301), .A2(KEYINPUT23), .A3(G119), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n339), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT24), .B(G110), .ZN(new_n347));
  OAI221_X1 g161(.A(new_n247), .B1(new_n338), .B2(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n338), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n349), .A2(new_n350), .B1(new_n231), .B2(new_n223), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n229), .A3(new_n228), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT76), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT22), .B(G137), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n348), .A2(new_n352), .A3(new_n357), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n285), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n337), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n361), .B(new_n285), .C1(KEYINPUT77), .C2(KEYINPUT25), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n336), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n335), .A2(G902), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G472), .A2(G902), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT11), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n305), .B2(G137), .ZN(new_n373));
  INV_X1    g187(.A(G137), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT11), .A3(G134), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n305), .A2(G137), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(G131), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n231), .B1(new_n202), .B2(new_n203), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n231), .A2(G143), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(KEYINPUT0), .A2(G128), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT0), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n301), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n385), .B2(KEYINPUT64), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n382), .B(new_n386), .C1(KEYINPUT64), .C2(new_n385), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT65), .ZN(new_n388));
  INV_X1    g202(.A(G143), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT65), .A2(G143), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(G146), .A3(new_n391), .ZN(new_n392));
  OR3_X1    g206(.A1(new_n389), .A2(KEYINPUT66), .A3(G146), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n231), .A2(G143), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT66), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n392), .A2(new_n393), .A3(new_n395), .A4(new_n385), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n378), .A2(new_n387), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n301), .A2(KEYINPUT1), .ZN(new_n398));
  AND4_X1   g212(.A1(new_n392), .A2(new_n393), .A3(new_n395), .A4(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT67), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n380), .B1(new_n197), .B2(new_n231), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT1), .B1(new_n389), .B2(G146), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G128), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n400), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n382), .A2(KEYINPUT67), .A3(new_n403), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n399), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n377), .A2(G131), .ZN(new_n408));
  INV_X1    g222(.A(new_n376), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n305), .A2(G137), .ZN(new_n410));
  OAI21_X1  g224(.A(G131), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n397), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n414), .A2(KEYINPUT68), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(KEYINPUT68), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n392), .A2(new_n393), .A3(new_n395), .A4(new_n398), .ZN(new_n418));
  AOI221_X4 g232(.A(new_n400), .B1(new_n402), .B2(G128), .C1(new_n379), .C2(new_n381), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT67), .B1(new_n382), .B2(new_n403), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n412), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n423), .A2(KEYINPUT68), .A3(new_n414), .A4(new_n397), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT2), .ZN(new_n426));
  INV_X1    g240(.A(G113), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT69), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT69), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT2), .A3(G113), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n428), .A2(new_n430), .B1(new_n426), .B2(new_n427), .ZN(new_n431));
  XNOR2_X1  g245(.A(G116), .B(G119), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT31), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n217), .A2(G210), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT27), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT26), .B(G101), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n431), .B(new_n432), .Z(new_n440));
  OAI211_X1 g254(.A(new_n397), .B(new_n440), .C1(new_n407), .C2(new_n412), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n434), .A2(new_n435), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT72), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n413), .A2(new_n433), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT28), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT28), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n439), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n440), .B1(new_n417), .B2(new_n424), .ZN(new_n451));
  INV_X1    g265(.A(new_n441), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT72), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n435), .A4(new_n439), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n443), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n439), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n451), .A2(new_n457), .A3(new_n452), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT71), .B1(new_n458), .B2(new_n435), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n434), .A2(new_n439), .A3(new_n441), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT71), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT31), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n371), .B1(new_n456), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n465));
  NOR4_X1   g279(.A1(new_n451), .A2(KEYINPUT31), .A3(new_n457), .A4(new_n452), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n449), .B1(new_n466), .B2(new_n454), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n467), .A2(new_n443), .A3(new_n459), .A4(new_n462), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT32), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n371), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT74), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n446), .A2(KEYINPUT29), .A3(new_n439), .A4(new_n448), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n285), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n457), .B1(new_n451), .B2(new_n452), .ZN(new_n475));
  INV_X1    g289(.A(new_n448), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(KEYINPUT28), .B2(new_n445), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT29), .B1(new_n477), .B2(new_n439), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G472), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n478), .A2(new_n475), .ZN(new_n482));
  OAI211_X1 g296(.A(KEYINPUT74), .B(G472), .C1(new_n482), .C2(new_n474), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n370), .B1(new_n471), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G214), .B1(G237), .B2(G902), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT80), .ZN(new_n487));
  INV_X1    g301(.A(new_n378), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n387), .A2(new_n396), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT3), .B1(new_n241), .B2(G107), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT3), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n292), .A3(G104), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n241), .A2(G107), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G101), .ZN(new_n496));
  INV_X1    g310(.A(G101), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n491), .A2(new_n493), .A3(new_n497), .A4(new_n494), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n500), .A3(G101), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n392), .A2(new_n395), .A3(new_n393), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n301), .B1(new_n379), .B2(KEYINPUT1), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n418), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n292), .A2(G104), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n241), .A2(G107), .ZN(new_n507));
  OAI21_X1  g321(.A(G101), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n498), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT10), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n490), .A2(new_n502), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n509), .A2(KEYINPUT78), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n498), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n421), .A2(KEYINPUT10), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n488), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n511), .A2(new_n512), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n499), .A2(new_n387), .A3(new_n396), .A4(new_n501), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n518), .A2(new_n520), .A3(new_n488), .A4(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT79), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n513), .A2(KEYINPUT79), .A3(new_n488), .A4(new_n518), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G140), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n192), .A2(G227), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n527), .B(new_n528), .Z(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n487), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(new_n525), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n511), .B1(new_n421), .B2(new_n517), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n533), .A2(new_n534), .A3(new_n378), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n533), .B2(new_n378), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n537), .A3(new_n530), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n532), .A2(new_n537), .A3(new_n487), .A4(new_n530), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G469), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n285), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n532), .A2(new_n537), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n529), .ZN(new_n545));
  INV_X1    g359(.A(new_n519), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n532), .A2(new_n530), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n542), .B1(new_n548), .B2(new_n277), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT82), .B(G224), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(G953), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n489), .A2(G125), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n225), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(KEYINPUT81), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT81), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n407), .B2(new_n225), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n553), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(KEYINPUT81), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n407), .A2(new_n557), .A3(new_n225), .ZN(new_n561));
  INV_X1    g375(.A(new_n553), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n554), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n433), .A2(new_n501), .A3(new_n499), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n432), .A2(KEYINPUT5), .ZN(new_n566));
  INV_X1    g380(.A(G116), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n567), .A2(KEYINPUT5), .A3(G119), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(new_n427), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n431), .A2(new_n432), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n517), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G122), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n565), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT6), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n565), .A2(new_n571), .ZN(new_n575));
  INV_X1    g389(.A(new_n572), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(KEYINPUT6), .A3(new_n573), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n564), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI211_X1 g394(.A(G125), .B(new_n399), .C1(new_n405), .C2(new_n406), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n581), .A2(new_n557), .B1(G125), .B2(new_n489), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n582), .A2(KEYINPUT7), .A3(new_n562), .A4(new_n560), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n572), .B(new_n584), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n570), .A2(new_n510), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n571), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n565), .A2(new_n571), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n587), .B1(new_n588), .B2(new_n572), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n556), .B2(new_n558), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n583), .A2(new_n589), .A3(new_n591), .A4(new_n559), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n580), .A2(new_n592), .A3(new_n277), .ZN(new_n593));
  OAI21_X1  g407(.A(G210), .B1(G237), .B2(G902), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT84), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n580), .A2(new_n592), .A3(new_n277), .A4(new_n594), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G221), .B1(new_n318), .B2(G902), .ZN(new_n599));
  AND4_X1   g413(.A1(new_n486), .A2(new_n551), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n334), .A2(new_n485), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  AOI21_X1  g416(.A(new_n480), .B1(new_n468), .B2(new_n285), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n464), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI211_X1 g419(.A(KEYINPUT95), .B(new_n480), .C1(new_n468), .C2(new_n285), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI211_X1 g422(.A(G469), .B(new_n363), .C1(new_n539), .C2(new_n540), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n369), .B(new_n599), .C1(new_n609), .C2(new_n549), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n273), .A2(new_n279), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n324), .A2(new_n613), .A3(new_n326), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n322), .A2(KEYINPUT33), .A3(new_n323), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n363), .A2(new_n328), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n614), .A2(KEYINPUT96), .A3(new_n615), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n327), .A2(new_n328), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT97), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n617), .A2(new_n618), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n621), .A4(new_n620), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n486), .ZN(new_n628));
  INV_X1    g442(.A(new_n594), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n593), .A2(new_n629), .ZN(new_n630));
  AOI211_X1 g444(.A(new_n288), .B(new_n628), .C1(new_n630), .C2(new_n597), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n612), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n611), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NAND3_X1  g449(.A1(new_n261), .A2(new_n272), .A3(KEYINPUT98), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n258), .A2(new_n637), .A3(new_n259), .A4(new_n260), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n636), .A2(new_n279), .A3(new_n330), .A4(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n631), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n611), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT35), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR2_X1   g459(.A1(new_n358), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n353), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n367), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n366), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n334), .A2(new_n607), .A3(new_n600), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  AOI21_X1  g468(.A(new_n628), .B1(new_n630), .B2(new_n597), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n551), .A2(new_n599), .A3(new_n655), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n468), .A2(new_n469), .A3(new_n371), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n469), .B1(new_n468), .B2(new_n371), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n484), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n286), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(G900), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT100), .Z(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(new_n283), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n639), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n656), .A2(new_n659), .A3(new_n664), .A4(new_n651), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT101), .B(G128), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G30));
  AOI21_X1  g481(.A(new_n331), .B1(new_n273), .B2(new_n279), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n598), .B(KEYINPUT38), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n486), .A3(new_n650), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n663), .B(new_n672), .Z(new_n673));
  NAND3_X1  g487(.A1(new_n551), .A2(new_n599), .A3(new_n673), .ZN(new_n674));
  AOI211_X1 g488(.A(new_n669), .B(new_n671), .C1(KEYINPUT40), .C2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n445), .A2(new_n439), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(G902), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n439), .B1(new_n451), .B2(new_n452), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n480), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n471), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n675), .B(new_n681), .C1(KEYINPUT40), .C2(new_n674), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n197), .ZN(G45));
  INV_X1    g497(.A(new_n663), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n612), .A2(new_n627), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n656), .A2(new_n659), .A3(new_n686), .A4(new_n651), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  NAND2_X1  g502(.A1(KEYINPUT103), .A2(G469), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n540), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n538), .B2(new_n531), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n690), .B1(new_n692), .B2(new_n363), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n541), .A2(new_n285), .A3(new_n689), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n693), .A2(new_n694), .A3(new_n599), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n659), .A2(new_n632), .A3(new_n369), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND4_X1  g512(.A1(new_n659), .A2(new_n641), .A3(new_n369), .A4(new_n695), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  AOI21_X1  g514(.A(new_n650), .B1(new_n471), .B2(new_n484), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n693), .A2(new_n694), .A3(new_n599), .A4(new_n655), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n334), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  OAI21_X1  g519(.A(new_n285), .B1(new_n456), .B2(new_n463), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n467), .B(new_n443), .C1(new_n435), .C2(new_n458), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n706), .A2(G472), .B1(new_n371), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n695), .A2(new_n369), .A3(new_n708), .A4(new_n289), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n655), .B1(new_n668), .B2(new_n710), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n261), .A2(new_n272), .B1(new_n278), .B2(G475), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n712), .A2(KEYINPUT104), .A3(new_n331), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT105), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n668), .A2(new_n710), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT104), .B1(new_n712), .B2(new_n331), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n655), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n709), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n296), .ZN(G24));
  NAND3_X1  g534(.A1(new_n686), .A2(new_n651), .A3(new_n708), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT106), .B1(new_n721), .B2(new_n702), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n706), .A2(G472), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n707), .A2(new_n371), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n651), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n685), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n703), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  NAND2_X1  g544(.A1(new_n599), .A2(new_n486), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n598), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n547), .A2(KEYINPUT107), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n526), .A2(new_n734), .A3(new_n530), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n545), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n542), .B1(new_n736), .B2(new_n277), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n732), .B1(new_n609), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g554(.A(KEYINPUT108), .B(new_n732), .C1(new_n609), .C2(new_n737), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n485), .A3(new_n686), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n485), .A3(KEYINPUT42), .A4(new_n686), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  AND3_X1   g562(.A1(new_n742), .A2(new_n485), .A3(new_n664), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n305), .ZN(G36));
  NOR2_X1   g564(.A1(new_n598), .A2(new_n628), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT43), .B1(new_n712), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n627), .A2(new_n712), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n608), .A3(new_n651), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n752), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n542), .B1(new_n548), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n761), .B2(new_n736), .ZN(new_n763));
  NAND2_X1  g577(.A1(G469), .A2(G902), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n543), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n767), .A2(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n766), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(KEYINPUT109), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n599), .A3(new_n673), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n760), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n599), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n599), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n659), .A2(new_n685), .A3(new_n369), .A4(new_n752), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NOR3_X1   g596(.A1(new_n755), .A2(new_n370), .A3(new_n731), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT111), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n693), .A2(new_n694), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT49), .Z(new_n786));
  NOR4_X1   g600(.A1(new_n784), .A2(new_n786), .A3(new_n670), .A4(new_n681), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT112), .ZN(new_n788));
  INV_X1    g602(.A(new_n695), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n789), .A2(new_n283), .A3(new_n752), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n756), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n725), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n369), .A2(new_n790), .A3(new_n471), .A4(new_n680), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n612), .A2(new_n627), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n789), .A2(new_n486), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n670), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n369), .A2(new_n756), .A3(new_n284), .A4(new_n708), .ZN(new_n800));
  OR2_X1    g614(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(new_n799), .B2(new_n800), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n795), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(KEYINPUT119), .ZN(new_n805));
  INV_X1    g619(.A(new_n599), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n785), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n777), .A2(new_n778), .A3(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n800), .A2(new_n751), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n804), .A2(KEYINPUT119), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n805), .A2(KEYINPUT51), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n793), .A2(new_n612), .A3(new_n627), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n280), .ZN(new_n814));
  INV_X1    g628(.A(new_n485), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n791), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT48), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n814), .B(new_n817), .C1(new_n703), .C2(new_n800), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n810), .A2(KEYINPUT116), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n810), .A2(KEYINPUT116), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n819), .A2(new_n820), .A3(new_n804), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n812), .B(new_n818), .C1(new_n821), .C2(KEYINPUT51), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n749), .B1(new_n745), .B2(new_n746), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n699), .A2(new_n696), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n712), .A2(new_n331), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n288), .B(new_n628), .C1(new_n596), .C2(new_n597), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n825), .B(new_n826), .C1(new_n712), .C2(new_n627), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n827), .A2(new_n605), .A3(new_n610), .A4(new_n606), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n719), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n652), .A2(new_n601), .A3(new_n704), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n551), .A2(new_n599), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n598), .A2(new_n330), .A3(new_n628), .A4(new_n663), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n279), .A2(new_n638), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n636), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n838), .A2(new_n701), .B1(new_n726), .B2(new_n742), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n823), .A2(new_n829), .A3(new_n830), .A4(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n701), .B(new_n656), .C1(new_n664), .C2(new_n686), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n727), .B1(new_n726), .B2(new_n703), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n725), .A2(new_n685), .A3(new_n702), .A4(KEYINPUT106), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n609), .A2(new_n737), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n845), .A2(new_n651), .A3(new_n806), .A4(new_n663), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n681), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n718), .B2(new_n714), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT114), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n714), .A2(new_n718), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n681), .A3(new_n846), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n729), .A2(new_n851), .A3(new_n852), .A4(new_n841), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n840), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n849), .A2(new_n853), .A3(KEYINPUT52), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(new_n849), .B2(new_n853), .ZN(new_n859));
  INV_X1    g673(.A(new_n844), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n855), .B1(new_n860), .B2(new_n851), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n859), .A2(new_n840), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n858), .B1(new_n862), .B2(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  INV_X1    g678(.A(new_n859), .ZN(new_n865));
  INV_X1    g679(.A(new_n840), .ZN(new_n866));
  INV_X1    g680(.A(new_n861), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT53), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  INV_X1    g683(.A(new_n857), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n859), .A3(new_n840), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n868), .B(new_n869), .C1(new_n871), .C2(KEYINPUT53), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n864), .A2(KEYINPUT115), .A3(new_n872), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n872), .A2(KEYINPUT115), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n822), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(G952), .A2(G953), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n788), .B1(new_n875), .B2(new_n876), .ZN(G75));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n856), .B2(new_n857), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n859), .A2(new_n840), .A3(new_n861), .A4(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n363), .B(new_n595), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n577), .A2(new_n579), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n564), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT55), .Z(new_n884));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n192), .A2(G952), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT120), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n363), .B(new_n629), .C1(new_n878), .C2(new_n880), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n884), .B1(new_n891), .B2(new_n885), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n890), .A2(KEYINPUT121), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT121), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(G51));
  OAI21_X1  g709(.A(new_n363), .B1(new_n878), .B2(new_n880), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n763), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT54), .B1(new_n878), .B2(new_n880), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n872), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n764), .B(KEYINPUT57), .Z(new_n900));
  AOI21_X1  g714(.A(new_n692), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n900), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n898), .B2(new_n872), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT122), .B1(new_n905), .B2(new_n692), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n888), .B1(new_n903), .B2(new_n906), .ZN(G54));
  NAND2_X1  g721(.A1(KEYINPUT58), .A2(G475), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n270), .B1(new_n896), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n888), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n896), .A2(new_n270), .A3(new_n908), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(G60));
  NAND2_X1  g727(.A1(G478), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT59), .Z(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n899), .A2(new_n614), .A3(new_n615), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n889), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n873), .A2(new_n874), .A3(new_n916), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n614), .A2(new_n615), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT123), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n878), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n868), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n647), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n928), .B(new_n889), .C1(new_n361), .C2(new_n927), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n927), .A2(new_n361), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n933), .A2(new_n889), .A3(new_n928), .A4(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(G66));
  OAI21_X1  g749(.A(G953), .B1(new_n287), .B2(new_n552), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n829), .A2(new_n830), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n938), .B2(G953), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT125), .Z(new_n940));
  INV_X1    g754(.A(G898), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n882), .B1(new_n941), .B2(G953), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n940), .B(new_n942), .ZN(G69));
  XNOR2_X1  g757(.A(new_n425), .B(new_n232), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n825), .B1(new_n712), .B2(new_n627), .ZN(new_n945));
  OR4_X1    g759(.A1(new_n815), .A2(new_n945), .A3(new_n674), .A4(new_n752), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n773), .A2(new_n781), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n860), .A2(new_n682), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT62), .ZN(new_n949));
  OR3_X1    g763(.A1(new_n947), .A2(KEYINPUT126), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT126), .B1(new_n947), .B2(new_n949), .ZN(new_n951));
  AOI211_X1 g765(.A(G953), .B(new_n944), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n944), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n773), .A2(new_n781), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n850), .A2(new_n485), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n860), .B(new_n823), .C1(new_n772), .C2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n192), .ZN(new_n958));
  NAND2_X1  g772(.A1(G900), .A2(G953), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n952), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n959), .ZN(new_n963));
  NAND2_X1  g777(.A1(G227), .A2(G900), .ZN(new_n964));
  AND4_X1   g778(.A1(G953), .A2(new_n963), .A3(new_n964), .A4(new_n944), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n962), .A2(new_n965), .ZN(G72));
  NAND3_X1  g780(.A1(new_n950), .A2(new_n938), .A3(new_n951), .ZN(new_n967));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT127), .Z(new_n970));
  AOI21_X1  g784(.A(new_n678), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n970), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n957), .B2(new_n938), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n453), .A2(new_n457), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n910), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n460), .A2(new_n475), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n863), .A2(new_n969), .A3(new_n976), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n971), .A2(new_n975), .A3(new_n977), .ZN(G57));
endmodule


