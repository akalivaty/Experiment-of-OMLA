

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  INV_X1 U322 ( .A(n557), .ZN(n458) );
  INV_X1 U323 ( .A(n523), .ZN(n535) );
  NOR2_X1 U324 ( .A1(n467), .A2(n526), .ZN(n533) );
  XNOR2_X1 U325 ( .A(n454), .B(KEYINPUT124), .ZN(n567) );
  AND2_X1 U326 ( .A1(n523), .A2(n453), .ZN(n454) );
  XOR2_X2 U327 ( .A(n575), .B(KEYINPUT41), .Z(n503) );
  XOR2_X1 U328 ( .A(n339), .B(n338), .Z(n290) );
  XNOR2_X1 U329 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n418) );
  XNOR2_X1 U330 ( .A(n419), .B(n418), .ZN(n531) );
  XNOR2_X1 U331 ( .A(n340), .B(n290), .ZN(n341) );
  XNOR2_X1 U332 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U333 ( .A(n348), .B(n404), .Z(n578) );
  XOR2_X1 U334 ( .A(n309), .B(n308), .Z(n523) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n455) );
  XNOR2_X1 U336 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(G183GAT), .B(KEYINPUT86), .Z(n292) );
  XNOR2_X1 U338 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n291) );
  XNOR2_X1 U339 ( .A(n292), .B(n291), .ZN(n304) );
  XOR2_X1 U340 ( .A(G15GAT), .B(G127GAT), .Z(n334) );
  XOR2_X1 U341 ( .A(KEYINPUT20), .B(G190GAT), .Z(n294) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(G99GAT), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U344 ( .A(n334), .B(n295), .Z(n297) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U347 ( .A(n298), .B(G71GAT), .Z(n302) );
  XOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n300) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n420) );
  XNOR2_X1 U351 ( .A(n420), .B(G176GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U354 ( .A(KEYINPUT85), .B(G134GAT), .Z(n306) );
  XNOR2_X1 U355 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(n307), .ZN(n437) );
  INV_X1 U358 ( .A(n437), .ZN(n308) );
  XOR2_X1 U359 ( .A(KEYINPUT93), .B(KEYINPUT90), .Z(n311) );
  XNOR2_X1 U360 ( .A(KEYINPUT22), .B(KEYINPUT95), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U362 ( .A(G211GAT), .B(KEYINPUT94), .Z(n313) );
  XNOR2_X1 U363 ( .A(KEYINPUT24), .B(KEYINPUT89), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U365 ( .A(n315), .B(n314), .Z(n325) );
  XNOR2_X1 U366 ( .A(G204GAT), .B(KEYINPUT21), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n316), .B(KEYINPUT92), .ZN(n317) );
  XOR2_X1 U368 ( .A(n317), .B(KEYINPUT91), .Z(n319) );
  XNOR2_X1 U369 ( .A(G197GAT), .B(G218GAT), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n429) );
  XNOR2_X1 U371 ( .A(G106GAT), .B(G78GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n320), .B(G148GAT), .ZN(n394) );
  XOR2_X1 U373 ( .A(n394), .B(KEYINPUT23), .Z(n322) );
  NAND2_X1 U374 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n429), .B(n323), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U378 ( .A(G22GAT), .B(G155GAT), .Z(n337) );
  XOR2_X1 U379 ( .A(n326), .B(n337), .Z(n329) );
  XOR2_X1 U380 ( .A(G50GAT), .B(G162GAT), .Z(n362) );
  XNOR2_X1 U381 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n327), .B(KEYINPUT2), .ZN(n436) );
  XNOR2_X1 U383 ( .A(n362), .B(n436), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n465) );
  XOR2_X1 U385 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n331) );
  XNOR2_X1 U386 ( .A(KEYINPUT14), .B(KEYINPUT83), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n344) );
  XOR2_X1 U388 ( .A(KEYINPUT81), .B(G211GAT), .Z(n333) );
  XNOR2_X1 U389 ( .A(G8GAT), .B(G183GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n427) );
  XOR2_X1 U391 ( .A(n334), .B(n427), .Z(n336) );
  NAND2_X1 U392 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n342) );
  XOR2_X1 U394 ( .A(KEYINPUT71), .B(G1GAT), .Z(n376) );
  XNOR2_X1 U395 ( .A(n376), .B(n337), .ZN(n340) );
  XOR2_X1 U396 ( .A(KEYINPUT12), .B(KEYINPUT84), .Z(n339) );
  XNOR2_X1 U397 ( .A(G78GAT), .B(G64GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U399 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n346) );
  XNOR2_X1 U400 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U402 ( .A(G57GAT), .B(n347), .Z(n404) );
  XNOR2_X1 U403 ( .A(KEYINPUT114), .B(n578), .ZN(n566) );
  XOR2_X1 U404 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n350) );
  XNOR2_X1 U405 ( .A(G134GAT), .B(KEYINPUT65), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n366) );
  XOR2_X1 U407 ( .A(G36GAT), .B(G190GAT), .Z(n423) );
  XOR2_X1 U408 ( .A(n423), .B(G92GAT), .Z(n352) );
  XOR2_X1 U409 ( .A(G99GAT), .B(G85GAT), .Z(n386) );
  XNOR2_X1 U410 ( .A(G218GAT), .B(n386), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n358) );
  XOR2_X1 U412 ( .A(G29GAT), .B(G43GAT), .Z(n354) );
  XNOR2_X1 U413 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n380) );
  XOR2_X1 U415 ( .A(KEYINPUT9), .B(n380), .Z(n356) );
  NAND2_X1 U416 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U418 ( .A(n358), .B(n357), .Z(n364) );
  XOR2_X1 U419 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n360) );
  XNOR2_X1 U420 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U424 ( .A(n366), .B(n365), .Z(n557) );
  NOR2_X1 U425 ( .A1(n566), .A2(n557), .ZN(n410) );
  XOR2_X1 U426 ( .A(G22GAT), .B(G197GAT), .Z(n368) );
  XNOR2_X1 U427 ( .A(G15GAT), .B(G141GAT), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U429 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n370) );
  XNOR2_X1 U430 ( .A(G8GAT), .B(KEYINPUT70), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n384) );
  XOR2_X1 U433 ( .A(G113GAT), .B(G36GAT), .Z(n374) );
  XNOR2_X1 U434 ( .A(G169GAT), .B(G50GAT), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U436 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U437 ( .A1(G229GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U439 ( .A(n379), .B(KEYINPUT29), .Z(n382) );
  XNOR2_X1 U440 ( .A(n380), .B(KEYINPUT68), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U442 ( .A(n384), .B(n383), .Z(n504) );
  INV_X1 U443 ( .A(n504), .ZN(n571) );
  XNOR2_X1 U444 ( .A(G176GAT), .B(G92GAT), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n385), .B(G64GAT), .ZN(n428) );
  XNOR2_X1 U446 ( .A(n428), .B(n386), .ZN(n390) );
  INV_X1 U447 ( .A(n390), .ZN(n388) );
  AND2_X1 U448 ( .A1(G230GAT), .A2(G233GAT), .ZN(n389) );
  INV_X1 U449 ( .A(n389), .ZN(n387) );
  NAND2_X1 U450 ( .A1(n388), .A2(n387), .ZN(n392) );
  NAND2_X1 U451 ( .A1(n390), .A2(n389), .ZN(n391) );
  NAND2_X1 U452 ( .A1(n392), .A2(n391), .ZN(n393) );
  XOR2_X1 U453 ( .A(n393), .B(KEYINPUT75), .Z(n396) );
  XNOR2_X1 U454 ( .A(n394), .B(KEYINPUT32), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U456 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n398) );
  XNOR2_X1 U457 ( .A(G120GAT), .B(G204GAT), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U459 ( .A(n400), .B(n399), .Z(n406) );
  XOR2_X1 U460 ( .A(KEYINPUT77), .B(KEYINPUT33), .Z(n402) );
  XNOR2_X1 U461 ( .A(KEYINPUT76), .B(KEYINPUT78), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U464 ( .A(n406), .B(n405), .Z(n575) );
  NAND2_X1 U465 ( .A1(n571), .A2(n503), .ZN(n408) );
  XOR2_X1 U466 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n409) );
  NAND2_X1 U468 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n411), .B(KEYINPUT47), .ZN(n417) );
  XOR2_X1 U470 ( .A(KEYINPUT67), .B(KEYINPUT45), .Z(n413) );
  XOR2_X1 U471 ( .A(KEYINPUT36), .B(n458), .Z(n581) );
  NAND2_X1 U472 ( .A1(n578), .A2(n581), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n415) );
  INV_X1 U474 ( .A(n575), .ZN(n457) );
  NAND2_X1 U475 ( .A1(n457), .A2(n504), .ZN(n414) );
  NOR2_X1 U476 ( .A1(n415), .A2(n414), .ZN(n416) );
  NOR2_X1 U477 ( .A1(n417), .A2(n416), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(KEYINPUT96), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n421), .B(KEYINPUT97), .ZN(n422) );
  XOR2_X1 U480 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U481 ( .A1(G226GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U483 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U485 ( .A(n431), .B(n430), .Z(n521) );
  XOR2_X1 U486 ( .A(n521), .B(KEYINPUT122), .Z(n432) );
  NOR2_X1 U487 ( .A1(n531), .A2(n432), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n433), .B(KEYINPUT54), .ZN(n450) );
  XOR2_X1 U489 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n435) );
  XNOR2_X1 U490 ( .A(G1GAT), .B(G57GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U492 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n439) );
  XOR2_X1 U493 ( .A(n437), .B(n436), .Z(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n449) );
  NAND2_X1 U496 ( .A1(G225GAT), .A2(G233GAT), .ZN(n447) );
  XOR2_X1 U497 ( .A(G155GAT), .B(G148GAT), .Z(n443) );
  XNOR2_X1 U498 ( .A(G29GAT), .B(G127GAT), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U500 ( .A(G162GAT), .B(G85GAT), .Z(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n518) );
  INV_X1 U504 ( .A(n518), .ZN(n532) );
  NAND2_X1 U505 ( .A1(n450), .A2(n532), .ZN(n569) );
  NOR2_X1 U506 ( .A1(n465), .A2(n569), .ZN(n452) );
  XNOR2_X1 U507 ( .A(KEYINPUT55), .B(KEYINPUT123), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U509 ( .A1(n567), .A2(n557), .ZN(n456) );
  XOR2_X1 U510 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n475) );
  NAND2_X1 U511 ( .A1(n571), .A2(n457), .ZN(n488) );
  NAND2_X1 U512 ( .A1(n458), .A2(n578), .ZN(n459) );
  XOR2_X1 U513 ( .A(KEYINPUT16), .B(n459), .Z(n473) );
  XOR2_X1 U514 ( .A(n521), .B(KEYINPUT98), .Z(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT27), .ZN(n467) );
  XOR2_X1 U516 ( .A(n465), .B(KEYINPUT28), .Z(n501) );
  INV_X1 U517 ( .A(n501), .ZN(n526) );
  NAND2_X1 U518 ( .A1(n535), .A2(n533), .ZN(n461) );
  NOR2_X1 U519 ( .A1(n532), .A2(n461), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT99), .ZN(n472) );
  INV_X1 U521 ( .A(n521), .ZN(n494) );
  NOR2_X1 U522 ( .A1(n535), .A2(n494), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n465), .A2(n463), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n464), .B(KEYINPUT25), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n465), .A2(n535), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n466), .B(KEYINPUT26), .ZN(n570) );
  NOR2_X1 U527 ( .A1(n570), .A2(n467), .ZN(n547) );
  INV_X1 U528 ( .A(n547), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n532), .A2(n470), .ZN(n471) );
  NAND2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n484) );
  NAND2_X1 U532 ( .A1(n473), .A2(n484), .ZN(n506) );
  NOR2_X1 U533 ( .A1(n488), .A2(n506), .ZN(n482) );
  NAND2_X1 U534 ( .A1(n482), .A2(n518), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U536 ( .A(G1GAT), .B(n476), .Z(G1324GAT) );
  NAND2_X1 U537 ( .A1(n521), .A2(n482), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n477), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n479) );
  NAND2_X1 U540 ( .A1(n482), .A2(n523), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n481) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT101), .Z(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U544 ( .A1(n526), .A2(n482), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U546 ( .A1(n581), .A2(n484), .ZN(n485) );
  NOR2_X1 U547 ( .A1(n578), .A2(n485), .ZN(n487) );
  XNOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(n517) );
  NOR2_X1 U550 ( .A1(n517), .A2(n488), .ZN(n490) );
  XNOR2_X1 U551 ( .A(KEYINPUT105), .B(KEYINPUT38), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n500) );
  NOR2_X1 U553 ( .A1(n500), .A2(n532), .ZN(n492) );
  XNOR2_X1 U554 ( .A(KEYINPUT103), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U556 ( .A(G29GAT), .B(n493), .Z(G1328GAT) );
  NOR2_X1 U557 ( .A1(n494), .A2(n500), .ZN(n495) );
  XOR2_X1 U558 ( .A(KEYINPUT106), .B(n495), .Z(n496) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  XNOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n498) );
  NOR2_X1 U561 ( .A1(n535), .A2(n500), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NOR2_X1 U564 ( .A1(n501), .A2(n500), .ZN(n502) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n508) );
  NAND2_X1 U567 ( .A1(n503), .A2(n504), .ZN(n505) );
  XOR2_X1 U568 ( .A(KEYINPUT109), .B(n505), .Z(n516) );
  NOR2_X1 U569 ( .A1(n516), .A2(n506), .ZN(n512) );
  NAND2_X1 U570 ( .A1(n512), .A2(n518), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n509), .Z(G1332GAT) );
  NAND2_X1 U573 ( .A1(n521), .A2(n512), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n523), .A2(n512), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n514) );
  NAND2_X1 U578 ( .A1(n512), .A2(n526), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n515), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT111), .Z(n520) );
  NOR2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n527), .A2(n518), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n527), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n527), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(KEYINPUT112), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n529) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n531), .A2(n532), .ZN(n548) );
  NAND2_X1 U595 ( .A1(n548), .A2(n533), .ZN(n534) );
  NOR2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n543), .A2(n571), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U600 ( .A1(n543), .A2(n503), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n542) );
  XOR2_X1 U603 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n540) );
  NAND2_X1 U604 ( .A1(n543), .A2(n566), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U608 ( .A1(n543), .A2(n557), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n549), .B(KEYINPUT119), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n571), .A2(n558), .ZN(n550) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n552) );
  NAND2_X1 U617 ( .A1(n558), .A2(n503), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  XOR2_X1 U620 ( .A(G155GAT), .B(KEYINPUT121), .Z(n556) );
  NAND2_X1 U621 ( .A1(n558), .A2(n578), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n567), .A2(n571), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT57), .B(KEYINPUT126), .Z(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT125), .B(n563), .Z(n565) );
  NAND2_X1 U631 ( .A1(n567), .A2(n503), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n580) );
  NAND2_X1 U636 ( .A1(n580), .A2(n571), .ZN(n574) );
  XOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .Z(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT59), .B(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n580), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n580), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

