//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202));
  XOR2_X1   g001(.A(G211gat), .B(G218gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT72), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n204), .A2(KEYINPUT72), .A3(new_n206), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n203), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G141gat), .B(G148gat), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  AND2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n217), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n219), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI211_X1 g026(.A(KEYINPUT75), .B(new_n217), .C1(new_n223), .C2(new_n224), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n218), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n222), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n215), .A2(new_n216), .A3(new_n226), .A4(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT3), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n214), .B1(new_n232), .B2(KEYINPUT29), .ZN(new_n233));
  NAND2_X1  g032(.A1(G228gat), .A2(G233gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n231), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n225), .A2(new_n226), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT75), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n225), .A2(new_n219), .A3(new_n226), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n236), .B1(new_n240), .B2(new_n218), .ZN(new_n241));
  INV_X1    g040(.A(new_n203), .ZN(new_n242));
  NAND2_X1  g041(.A1(G211gat), .A2(G218gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT22), .ZN(new_n244));
  OR2_X1    g043(.A1(G197gat), .A2(G204gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(G197gat), .A2(G204gat), .ZN(new_n246));
  AOI221_X4 g045(.A(new_n208), .B1(new_n243), .B2(new_n244), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT72), .B1(new_n204), .B2(new_n206), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n242), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT29), .B1(new_n249), .B2(new_n212), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n241), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n233), .A2(new_n235), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(new_n250), .B2(KEYINPUT79), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT79), .B(new_n255), .C1(new_n211), .C2(new_n213), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n241), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT80), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n233), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT80), .B(new_n214), .C1(new_n232), .C2(KEYINPUT29), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n252), .B1(new_n262), .B2(new_n234), .ZN(new_n263));
  INV_X1    g062(.A(G22gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n202), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT31), .B(G50gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n234), .ZN(new_n270));
  INV_X1    g069(.A(new_n252), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n264), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI211_X1 g071(.A(G22gat), .B(new_n252), .C1(new_n262), .C2(new_n234), .ZN(new_n273));
  OAI22_X1  g072(.A1(new_n265), .A2(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G22gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n263), .A2(new_n264), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(new_n202), .A3(new_n277), .A4(new_n268), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G134gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(KEYINPUT70), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G120gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(KEYINPUT1), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(G120gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(G113gat), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n284), .B(new_n280), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G127gat), .ZN(new_n291));
  INV_X1    g090(.A(G127gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n283), .A2(new_n292), .A3(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT24), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n303), .B(new_n304), .C1(G183gat), .C2(G190gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT25), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n299), .A4(new_n297), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n308), .A2(KEYINPUT64), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n304), .A2(KEYINPUT65), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n315), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n311), .A2(new_n313), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n307), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n314), .A2(new_n316), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n320), .A2(KEYINPUT66), .A3(new_n311), .A4(new_n313), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n306), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT27), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT27), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G183gat), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n324), .B1(new_n326), .B2(G183gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n310), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n323), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT28), .A4(new_n310), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT26), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n297), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n334), .B(new_n301), .C1(new_n336), .C2(new_n295), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT69), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT69), .ZN(new_n340));
  AOI211_X1 g139(.A(new_n340), .B(new_n337), .C1(new_n331), .C2(new_n332), .ZN(new_n341));
  OAI22_X1  g140(.A1(new_n322), .A2(KEYINPUT67), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n314), .B(new_n316), .C1(KEYINPUT64), .C2(new_n308), .ZN(new_n343));
  OAI22_X1  g142(.A1(new_n303), .A2(new_n312), .B1(G183gat), .B2(G190gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n318), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n307), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n321), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n306), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT67), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n294), .B1(new_n342), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G227gat), .ZN(new_n353));
  INV_X1    g152(.A(G233gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n339), .A2(new_n341), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n349), .A2(new_n350), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n322), .A2(KEYINPUT67), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n283), .A2(new_n292), .A3(new_n289), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n292), .B1(new_n283), .B2(new_n289), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n356), .A2(new_n357), .A3(new_n358), .A4(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n355), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT32), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT33), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G71gat), .B(G99gat), .Z(new_n367));
  XNOR2_X1  g166(.A(G15gat), .B(G43gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT71), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n364), .B1(new_n369), .B2(KEYINPUT33), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n363), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n371), .B1(new_n363), .B2(new_n372), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT34), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n352), .A2(new_n362), .ZN(new_n377));
  INV_X1    g176(.A(new_n355), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI211_X1 g178(.A(KEYINPUT34), .B(new_n355), .C1(new_n352), .C2(new_n362), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n383), .B(new_n370), .C1(new_n374), .C2(new_n373), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT84), .B1(new_n279), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n274), .A2(new_n278), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n382), .A4(new_n384), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n241), .B2(new_n361), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n229), .A2(new_n231), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n294), .A3(KEYINPUT76), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n241), .A2(new_n361), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n391), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n393), .A2(new_n401), .A3(new_n395), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n253), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n229), .A2(KEYINPUT3), .A3(new_n231), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n361), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n394), .A2(new_n294), .A3(KEYINPUT4), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n402), .A2(new_n398), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT4), .B1(new_n394), .B2(new_n294), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n395), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(KEYINPUT4), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n405), .A2(new_n391), .A3(new_n398), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n400), .A2(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G57gat), .B(G85gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT78), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT6), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n407), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n410), .A2(new_n411), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(KEYINPUT6), .A3(new_n423), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n342), .B2(new_n351), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n337), .B1(new_n331), .B2(new_n332), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n347), .B2(new_n348), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n428), .B1(new_n432), .B2(KEYINPUT29), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT73), .ZN(new_n434));
  INV_X1    g233(.A(new_n214), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT73), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n436), .B(new_n428), .C1(new_n432), .C2(KEYINPUT29), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n430), .A2(new_n434), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n255), .B(new_n428), .C1(new_n342), .C2(new_n351), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n429), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n214), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n438), .A2(new_n441), .A3(new_n445), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT30), .A3(new_n448), .ZN(new_n449));
  OR3_X1    g248(.A1(new_n442), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n427), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT35), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n390), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n279), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT36), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n385), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n382), .A2(new_n384), .A3(KEYINPUT36), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n394), .A2(new_n294), .A3(KEYINPUT76), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT76), .B1(new_n394), .B2(new_n294), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT4), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n408), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n405), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT39), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n399), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n418), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT39), .B1(new_n397), .B2(new_n399), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n470), .B1(new_n399), .B2(new_n466), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n461), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT40), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT40), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n461), .B(new_n474), .C1(new_n469), .C2(new_n471), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n424), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n387), .B1(new_n476), .B2(new_n451), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n425), .A2(new_n426), .A3(new_n448), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n214), .B1(new_n439), .B2(new_n440), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n430), .A2(new_n434), .A3(new_n437), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n214), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(KEYINPUT83), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n485), .A3(new_n214), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n480), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n446), .B1(new_n442), .B2(KEYINPUT37), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n479), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n479), .B1(new_n442), .B2(KEYINPUT37), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(new_n446), .C1(KEYINPUT37), .C2(new_n442), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n478), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n456), .B(new_n460), .C1(new_n477), .C2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n385), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n494), .A2(new_n427), .A3(new_n387), .A4(new_n451), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n453), .ZN(new_n496));
  AND4_X1   g295(.A1(KEYINPUT85), .A2(new_n455), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n390), .A2(new_n454), .B1(new_n453), .B2(new_n495), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT85), .B1(new_n498), .B2(new_n493), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G36gat), .ZN(new_n501));
  AND2_X1   g300(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G29gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n509));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n509), .B2(new_n510), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n513));
  OR3_X1    g312(.A1(new_n512), .A2(KEYINPUT87), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT87), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(G1gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(G1gat), .B2(new_n519), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G8gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n512), .A2(new_n523), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n512), .B(new_n523), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n526), .B(KEYINPUT13), .Z(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT88), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G197gat), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT11), .B(G169gat), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n541), .B(KEYINPUT12), .Z(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n516), .A2(new_n524), .B1(new_n523), .B2(new_n512), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(KEYINPUT18), .A3(new_n526), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n530), .A2(new_n537), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n528), .A2(new_n529), .B1(new_n534), .B2(new_n536), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n543), .B1(new_n548), .B2(new_n545), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n500), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(new_n221), .ZN(new_n553));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G71gat), .B(G78gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G127gat), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n523), .B1(KEYINPUT21), .B2(new_n561), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n564), .B(new_n292), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(new_n566), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n556), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n566), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n567), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n555), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT92), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT91), .B(G92gat), .Z(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(KEYINPUT89), .A2(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n579), .A2(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT8), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(KEYINPUT90), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(KEYINPUT90), .B2(new_n585), .ZN(new_n587));
  AND2_X1   g386(.A1(KEYINPUT89), .A2(KEYINPUT7), .ZN(new_n588));
  OR3_X1    g387(.A1(new_n588), .A2(new_n581), .A3(new_n582), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G99gat), .B(G106gat), .Z(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n518), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n516), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n595), .A2(new_n512), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n578), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  NAND3_X1  g404(.A1(new_n597), .A2(new_n578), .A3(new_n599), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n601), .A2(new_n602), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(KEYINPUT93), .ZN(new_n608));
  INV_X1    g407(.A(new_n606), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(new_n600), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n561), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n592), .A2(new_n561), .A3(new_n593), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n615), .A2(new_n614), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT94), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n617), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n619), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n619), .B1(new_n613), .B2(new_n615), .ZN(new_n625));
  XOR2_X1   g424(.A(G120gat), .B(G148gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT95), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  NOR2_X1   g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n621), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n618), .A2(new_n620), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n629), .B1(new_n632), .B2(new_n625), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n575), .A2(new_n611), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n551), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n427), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(G1gat), .Z(G1324gat));
  INV_X1    g439(.A(new_n451), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  NAND4_X1  g441(.A1(new_n551), .A2(new_n641), .A3(new_n637), .A4(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n643), .A2(KEYINPUT96), .A3(KEYINPUT42), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT42), .B1(new_n643), .B2(KEYINPUT96), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n551), .A2(new_n641), .A3(new_n637), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n646), .A2(KEYINPUT97), .A3(G8gat), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT97), .B1(new_n646), .B2(G8gat), .ZN(new_n648));
  OAI22_X1  g447(.A1(new_n644), .A2(new_n645), .B1(new_n647), .B2(new_n648), .ZN(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n638), .B2(new_n460), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n385), .A2(G15gat), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n638), .B2(new_n651), .ZN(G1326gat));
  NOR2_X1   g451(.A1(new_n638), .A2(new_n387), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT43), .B(G22gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NOR2_X1   g454(.A1(new_n575), .A2(new_n634), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n611), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n500), .A2(new_n550), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n660), .A2(G29gat), .A3(new_n427), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT98), .B(KEYINPUT45), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n611), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n497), .B2(new_n499), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n455), .A2(new_n493), .A3(new_n496), .ZN(new_n668));
  INV_X1    g467(.A(new_n611), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n665), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n547), .A2(new_n549), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675), .B2(new_n427), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n663), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n664), .A2(new_n676), .A3(new_n677), .ZN(G1328gat));
  NOR3_X1   g477(.A1(new_n660), .A2(G36gat), .A3(new_n451), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT46), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G36gat), .B1(new_n675), .B2(new_n451), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(G1329gat));
  INV_X1    g483(.A(new_n460), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n672), .A2(new_n685), .A3(new_n674), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(G43gat), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT47), .B1(new_n687), .B2(KEYINPUT99), .ZN(new_n688));
  INV_X1    g487(.A(G43gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n659), .A2(new_n689), .A3(new_n494), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n687), .B(new_n690), .C1(KEYINPUT99), .C2(KEYINPUT47), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(G1330gat));
  NOR2_X1   g493(.A1(new_n387), .A2(G50gat), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n667), .A2(new_n279), .A3(new_n671), .A4(new_n674), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n659), .A2(new_n695), .B1(new_n696), .B2(G50gat), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(KEYINPUT100), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1331gat));
  NAND4_X1  g499(.A1(new_n673), .A2(new_n575), .A3(new_n611), .A4(new_n634), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n498), .B2(new_n493), .ZN(new_n702));
  INV_X1    g501(.A(new_n427), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT101), .B(G57gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1332gat));
  AOI21_X1  g505(.A(new_n451), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT102), .ZN(new_n709));
  NOR2_X1   g508(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1333gat));
  NAND2_X1  g510(.A1(new_n702), .A2(new_n685), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n385), .A2(G71gat), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n712), .A2(G71gat), .B1(new_n702), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g514(.A1(new_n702), .A2(new_n279), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT103), .B(G78gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1335gat));
  NOR3_X1   g517(.A1(new_n550), .A2(new_n575), .A3(new_n635), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n672), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G85gat), .B1(new_n720), .B2(new_n427), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n550), .A2(new_n575), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n668), .A2(new_n669), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n668), .A2(KEYINPUT51), .A3(new_n669), .A4(new_n722), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n723), .A2(KEYINPUT104), .A3(new_n724), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(new_n634), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n703), .A2(new_n580), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n721), .B1(new_n730), .B2(new_n731), .ZN(G1336gat));
  NOR3_X1   g531(.A1(new_n635), .A2(new_n451), .A3(G92gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n728), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n728), .A2(new_n736), .A3(new_n729), .A4(new_n733), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n667), .A2(new_n641), .A3(new_n671), .A4(new_n719), .ZN(new_n738));
  INV_X1    g537(.A(new_n579), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n735), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n735), .A2(new_n740), .A3(KEYINPUT106), .A4(new_n737), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n738), .A2(new_n739), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n725), .A2(new_n727), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(new_n733), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT52), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n749), .ZN(G1337gat));
  OAI21_X1  g549(.A(G99gat), .B1(new_n720), .B2(new_n460), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n385), .A2(G99gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n730), .B2(new_n752), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n672), .A2(new_n279), .A3(new_n719), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT107), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n672), .A2(new_n756), .A3(new_n279), .A4(new_n719), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n755), .A2(G106gat), .A3(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n387), .A2(new_n635), .A3(G106gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n728), .A2(new_n729), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n754), .A2(G106gat), .B1(new_n747), .B2(new_n759), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n758), .A2(new_n762), .B1(new_n761), .B2(new_n763), .ZN(G1339gat));
  NOR2_X1   g563(.A1(new_n636), .A2(new_n550), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT108), .B1(new_n636), .B2(new_n550), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n616), .A2(new_n617), .A3(new_n772), .A4(new_n620), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n774), .A2(new_n621), .A3(KEYINPUT54), .A4(new_n624), .ZN(new_n775));
  INV_X1    g574(.A(new_n629), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n632), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(KEYINPUT55), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n631), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n544), .A2(new_n526), .B1(new_n531), .B2(new_n532), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n541), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n546), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT55), .B1(new_n775), .B2(new_n778), .ZN(new_n784));
  NOR4_X1   g583(.A1(new_n780), .A2(new_n611), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n634), .A2(new_n546), .A3(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT110), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n634), .A2(new_n546), .A3(new_n788), .A4(new_n782), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n631), .B(new_n779), .C1(new_n547), .C2(new_n549), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n787), .B(new_n789), .C1(new_n790), .C2(new_n784), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n785), .B1(new_n791), .B2(new_n611), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n769), .B1(new_n792), .B2(new_n575), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n387), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n794), .A2(KEYINPUT111), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n385), .B1(new_n794), .B2(KEYINPUT111), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n703), .A2(new_n451), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(G113gat), .A3(new_n550), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n793), .A2(new_n703), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n390), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n451), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n285), .B1(new_n804), .B2(new_n673), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n801), .A2(new_n805), .ZN(G1340gat));
  NAND3_X1  g605(.A1(new_n800), .A2(G120gat), .A3(new_n634), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n287), .B1(new_n804), .B2(new_n635), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(G1341gat));
  NAND2_X1  g608(.A1(new_n797), .A2(new_n799), .ZN(new_n810));
  INV_X1    g609(.A(new_n575), .ZN(new_n811));
  XNOR2_X1  g610(.A(KEYINPUT70), .B(G127gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n803), .A2(new_n451), .A3(new_n575), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n812), .ZN(G1342gat));
  NOR2_X1   g614(.A1(new_n641), .A2(new_n611), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n803), .A2(new_n280), .A3(new_n816), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(KEYINPUT56), .Z(new_n818));
  OAI21_X1  g617(.A(G134gat), .B1(new_n810), .B2(new_n611), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1343gat));
  INV_X1    g619(.A(new_n785), .ZN(new_n821));
  INV_X1    g620(.A(new_n786), .ZN(new_n822));
  INV_X1    g621(.A(new_n790), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n775), .B2(new_n778), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT55), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n775), .A2(new_n824), .A3(new_n778), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n822), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n821), .B1(new_n830), .B2(new_n669), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n831), .A2(new_n811), .B1(new_n768), .B2(new_n767), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT57), .B1(new_n832), .B2(new_n387), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n799), .A2(new_n460), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT112), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n793), .A2(new_n279), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n833), .B(new_n835), .C1(KEYINPUT57), .C2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G141gat), .B1(new_n837), .B2(new_n673), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n793), .A2(new_n703), .A3(new_n279), .A4(new_n460), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n641), .ZN(new_n840));
  INV_X1    g639(.A(G141gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n550), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(G1344gat));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n846), .B(G148gat), .C1(new_n837), .C2(new_n635), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n836), .A2(KEYINPUT57), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n835), .A2(new_n634), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n575), .B1(new_n831), .B2(KEYINPUT115), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n827), .A2(new_n825), .A3(KEYINPUT55), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n786), .B1(new_n852), .B2(new_n790), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n785), .B1(new_n853), .B2(new_n611), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n765), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n387), .A2(KEYINPUT57), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n849), .B(new_n850), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G148gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n848), .B1(new_n861), .B2(KEYINPUT59), .ZN(new_n862));
  AOI211_X1 g661(.A(KEYINPUT116), .B(new_n846), .C1(new_n860), .C2(G148gat), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n847), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(G148gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n840), .A2(new_n865), .A3(new_n634), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(G1345gat));
  OAI21_X1  g666(.A(G155gat), .B1(new_n837), .B2(new_n811), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n840), .A2(new_n221), .A3(new_n575), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1346gat));
  OAI21_X1  g669(.A(G162gat), .B1(new_n837), .B2(new_n611), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n816), .A2(new_n222), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n839), .B2(new_n872), .ZN(G1347gat));
  NOR2_X1   g672(.A1(new_n703), .A2(new_n451), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n797), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(G169gat), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(new_n673), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n793), .A2(new_n427), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n451), .B1(new_n386), .B2(new_n389), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(G169gat), .B1(new_n880), .B2(new_n550), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n877), .A2(new_n881), .ZN(G1348gat));
  OAI21_X1  g681(.A(G176gat), .B1(new_n875), .B2(new_n635), .ZN(new_n883));
  INV_X1    g682(.A(G176gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n884), .A3(new_n634), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1349gat));
  AND3_X1   g685(.A1(new_n575), .A2(new_n325), .A3(new_n327), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n878), .A2(new_n879), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n878), .A2(KEYINPUT117), .A3(new_n879), .A4(new_n887), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n890), .A2(new_n891), .B1(new_n892), .B2(KEYINPUT60), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(KEYINPUT60), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n795), .A2(new_n796), .A3(new_n575), .A4(new_n874), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G183gat), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n894), .B1(new_n893), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n797), .A2(new_n669), .A3(new_n874), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G190gat), .ZN(new_n901));
  XNOR2_X1  g700(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(G190gat), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n880), .A2(new_n310), .A3(new_n669), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n903), .A2(new_n905), .A3(new_n908), .ZN(G1351gat));
  NOR3_X1   g708(.A1(new_n685), .A2(new_n387), .A3(new_n451), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n878), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912), .B2(new_n550), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n849), .B1(new_n857), .B2(new_n859), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT121), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n793), .B2(new_n279), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n831), .A2(KEYINPUT115), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n811), .B1(new_n854), .B2(new_n855), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n918), .A2(new_n919), .B1(new_n550), .B2(new_n636), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n917), .B1(new_n920), .B2(new_n858), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n460), .A2(new_n874), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT122), .ZN(new_n926));
  INV_X1    g725(.A(G197gat), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n926), .A2(new_n927), .A3(new_n673), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n913), .B1(new_n924), .B2(new_n928), .ZN(G1352gat));
  AND2_X1   g728(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n930));
  NOR2_X1   g729(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g731(.A(KEYINPUT123), .B(G204gat), .Z(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n911), .A2(new_n635), .A3(new_n934), .ZN(new_n935));
  MUX2_X1   g734(.A(new_n932), .B(new_n930), .S(new_n935), .Z(new_n936));
  AOI211_X1 g735(.A(new_n635), .B(new_n926), .C1(new_n915), .C2(new_n923), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n933), .ZN(G1353gat));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  INV_X1    g738(.A(G211gat), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n811), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n921), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n942), .B2(KEYINPUT63), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n849), .B(new_n941), .C1(new_n857), .C2(new_n859), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G211gat), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(KEYINPUT126), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT125), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n944), .A2(new_n950), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n943), .A2(new_n947), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n912), .A2(new_n940), .A3(new_n575), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1354gat));
  AOI21_X1  g753(.A(G218gat), .B1(new_n912), .B2(new_n669), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n669), .A2(G218gat), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT127), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n926), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n955), .B1(new_n924), .B2(new_n958), .ZN(G1355gat));
endmodule


