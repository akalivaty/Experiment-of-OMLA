//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(KEYINPUT22), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n202), .B1(new_n209), .B2(KEYINPUT29), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G141gat), .ZN(new_n216));
  INV_X1    g015(.A(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT79), .A3(new_n212), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n215), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n222), .B1(new_n220), .B2(new_n223), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT80), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n230));
  INV_X1    g029(.A(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT2), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n229), .B(new_n230), .C1(new_n234), .C2(new_n222), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n225), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n210), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n225), .A2(new_n202), .A3(new_n228), .A4(new_n235), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n209), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G78gat), .B(G106gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G228gat), .A2(G233gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(G22gat), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT31), .B(G50gat), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n244), .B(new_n248), .Z(new_n249));
  INV_X1    g048(.A(KEYINPUT32), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n251));
  INV_X1    g050(.A(G183gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT27), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT27), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G183gat), .ZN(new_n255));
  INV_X1    g054(.A(G190gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n257), .A2(new_n259), .B1(G183gat), .B2(G190gat), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT26), .B1(new_n263), .B2(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n261), .A4(new_n262), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT27), .B(G183gat), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(KEYINPUT66), .A3(new_n258), .A4(new_n256), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n260), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT65), .B(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT23), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(G176gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n265), .A2(KEYINPUT23), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n273), .A2(new_n275), .B1(new_n263), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n281), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT64), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT25), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n280), .A2(new_n283), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n276), .A2(new_n263), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n289), .B1(new_n275), .B2(new_n261), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n272), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G120gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G113gat), .ZN(new_n294));
  INV_X1    g093(.A(G113gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G120gat), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT1), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n298));
  XNOR2_X1  g097(.A(G127gat), .B(G134gat), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n297), .ZN(new_n301));
  INV_X1    g100(.A(G134gat), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n304));
  INV_X1    g103(.A(G127gat), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT69), .B1(new_n302), .B2(G127gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n305), .A3(G134gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n301), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n298), .B1(new_n297), .B2(new_n299), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n300), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n251), .B1(new_n292), .B2(new_n313), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n261), .A2(KEYINPUT65), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G169gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n275), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n288), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n289), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n307), .A2(new_n309), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT68), .B(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G127gat), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n297), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n294), .A2(new_n296), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n299), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT70), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n324), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n323), .A2(new_n333), .A3(KEYINPUT71), .A4(new_n272), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n292), .A2(new_n313), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n314), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n250), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT33), .B1(new_n336), .B2(new_n338), .ZN(new_n340));
  XOR2_X1   g139(.A(G15gat), .B(G43gat), .Z(new_n341));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n339), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  AOI221_X4 g144(.A(new_n250), .B1(KEYINPUT33), .B2(new_n343), .C1(new_n336), .C2(new_n338), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n314), .A2(new_n337), .A3(new_n334), .A4(new_n335), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT34), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n337), .B2(KEYINPUT73), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n349), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n314), .A2(new_n335), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n337), .A4(new_n334), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n352), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n347), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n338), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT32), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT33), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n366), .A3(new_n343), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n353), .B1(new_n349), .B2(new_n350), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n339), .B1(new_n340), .B2(new_n344), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n357), .A2(new_n352), .A3(new_n358), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n249), .B1(new_n362), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(new_n292), .B2(new_n239), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n323), .B2(new_n272), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n209), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n292), .A2(new_n375), .ZN(new_n379));
  INV_X1    g178(.A(new_n209), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n323), .B2(new_n272), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n379), .B(new_n380), .C1(new_n381), .C2(new_n375), .ZN(new_n382));
  XOR2_X1   g181(.A(G8gat), .B(G36gat), .Z(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT30), .A4(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT77), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n378), .B2(new_n382), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n378), .A2(new_n382), .A3(new_n385), .ZN(new_n389));
  XOR2_X1   g188(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n228), .A2(new_n235), .ZN(new_n393));
  INV_X1    g192(.A(new_n224), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT2), .B1(new_n227), .B2(new_n211), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n219), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n333), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n313), .A2(new_n236), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT81), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(KEYINPUT5), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT3), .B1(new_n393), .B2(new_n396), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(new_n238), .A3(new_n313), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n313), .B2(new_n236), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n397), .A2(KEYINPUT4), .A3(new_n333), .ZN(new_n408));
  INV_X1    g207(.A(new_n402), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n405), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT82), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n410), .A2(new_n412), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n403), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT0), .ZN(new_n417));
  XNOR2_X1  g216(.A(G57gat), .B(G85gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421));
  INV_X1    g220(.A(new_n419), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(new_n403), .C1(new_n413), .C2(new_n414), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  OR3_X1    g223(.A1(new_n415), .A2(new_n421), .A3(new_n419), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n392), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n367), .A2(new_n369), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n427), .A2(KEYINPUT72), .B1(new_n370), .B2(new_n368), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT72), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n367), .A2(new_n429), .A3(new_n369), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT75), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT72), .B1(new_n345), .B2(new_n346), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n368), .A2(new_n370), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n432), .A2(KEYINPUT75), .A3(new_n430), .A4(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n373), .B(new_n426), .C1(new_n431), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT35), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n427), .A2(new_n433), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI211_X1 g238(.A(new_n249), .B(new_n439), .C1(new_n372), .C2(new_n362), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n441), .A2(KEYINPUT35), .A3(new_n392), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n445), .B1(new_n362), .B2(new_n372), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n431), .B2(new_n435), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n361), .B1(new_n347), .B2(new_n360), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n438), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n445), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n244), .B(new_n248), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n424), .A2(new_n425), .ZN(new_n454));
  INV_X1    g253(.A(new_n392), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT37), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n378), .A2(new_n382), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT85), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n378), .A2(new_n382), .A3(new_n460), .A4(new_n457), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT38), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n378), .A2(new_n382), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n385), .B1(new_n464), .B2(KEYINPUT37), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n462), .A2(KEYINPUT86), .A3(new_n463), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n462), .A2(new_n465), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT38), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n441), .A2(new_n470), .A3(new_n389), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT39), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n402), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n476), .A2(new_n419), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n474), .B2(new_n402), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n398), .A2(new_n399), .A3(new_n409), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT83), .A4(new_n409), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n477), .A2(KEYINPUT40), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n423), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n476), .A2(new_n419), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n483), .B2(new_n478), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n489), .B2(KEYINPUT40), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n477), .A2(new_n484), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(KEYINPUT84), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n486), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n249), .B1(new_n494), .B2(new_n392), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n456), .B1(new_n473), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n452), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n444), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G36gat), .ZN(new_n499));
  AND2_X1   g298(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G29gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n505), .A2(KEYINPUT15), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(KEYINPUT15), .ZN(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(KEYINPUT17), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n509), .B2(new_n510), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(G1gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  MUX2_X1   g317(.A(G1gat), .B(new_n517), .S(new_n518), .Z(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT89), .B(G8gat), .Z(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n519), .B2(new_n523), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n515), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT91), .B1(new_n525), .B2(new_n526), .ZN(new_n530));
  INV_X1    g329(.A(new_n526), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n531), .A2(new_n521), .A3(new_n532), .A4(new_n524), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n533), .A3(new_n511), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n528), .A2(KEYINPUT18), .A3(new_n529), .A4(new_n534), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(new_n529), .ZN(new_n540));
  INV_X1    g339(.A(new_n534), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n511), .B1(new_n530), .B2(new_n533), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT88), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G113gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(new_n216), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n547), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT12), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n543), .A4(new_n551), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n498), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT93), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G57gat), .B(G64gat), .Z(new_n559));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  INV_X1    g360(.A(G71gat), .ZN(new_n562));
  INV_X1    g361(.A(G78gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G71gat), .B(G78gat), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n565), .B(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(KEYINPUT21), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT95), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G183gat), .B(G211gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n530), .A2(new_n533), .B1(KEYINPUT21), .B2(new_n568), .ZN(new_n575));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n575), .B(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT7), .ZN(new_n584));
  XNOR2_X1  g383(.A(G99gat), .B(G106gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n584), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n585), .B1(new_n584), .B2(new_n589), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT97), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(new_n512), .B2(new_n514), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n593), .B(KEYINPUT98), .C1(new_n512), .C2(new_n514), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n590), .A2(new_n591), .ZN(new_n599));
  AND2_X1   g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n511), .A2(new_n599), .B1(KEYINPUT41), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n598), .A2(new_n601), .A3(new_n603), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n600), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT96), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n609), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n603), .B1(new_n598), .B2(new_n601), .ZN(new_n613));
  INV_X1    g412(.A(new_n601), .ZN(new_n614));
  AOI211_X1 g413(.A(new_n614), .B(new_n604), .C1(new_n596), .C2(new_n597), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n612), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n611), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n605), .A2(KEYINPUT99), .A3(new_n606), .A4(new_n610), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n582), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n568), .A2(new_n599), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n565), .A2(new_n566), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n565), .A2(new_n566), .ZN(new_n625));
  OAI22_X1  g424(.A1(new_n624), .A2(new_n625), .B1(new_n590), .B2(new_n591), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n592), .B(KEYINPUT100), .C1(new_n624), .C2(new_n625), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT10), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n622), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n622), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n628), .A2(new_n634), .A3(new_n629), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n635), .A3(new_n639), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n621), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n558), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n441), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g446(.A(new_n520), .B1(new_n645), .B2(new_n392), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n558), .A2(new_n644), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n649), .A2(new_n455), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT42), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n652), .A2(KEYINPUT42), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n649), .B2(new_n452), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n450), .A2(G15gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n649), .B2(new_n657), .ZN(G1326gat));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n645), .B2(new_n249), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n649), .A2(KEYINPUT101), .A3(new_n453), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n645), .A2(new_n661), .A3(new_n249), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT101), .B1(new_n649), .B2(new_n453), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n659), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(G1327gat));
  INV_X1    g467(.A(new_n582), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n618), .A2(new_n619), .ZN(new_n670));
  INV_X1    g469(.A(new_n643), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT102), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n558), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n454), .A2(G29gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n675), .A2(new_n680), .A3(new_n676), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n620), .B1(new_n444), .B2(new_n497), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT104), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n437), .A2(new_n443), .B1(new_n452), .B2(new_n496), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n685), .B(KEYINPUT44), .C1(new_n686), .C2(new_n620), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n456), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n468), .A2(new_n469), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n472), .A2(new_n424), .A3(new_n425), .A4(new_n389), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n485), .A2(new_n423), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT84), .B1(new_n491), .B2(new_n492), .ZN(new_n694));
  AOI211_X1 g493(.A(new_n487), .B(KEYINPUT40), .C1(new_n477), .C2(new_n484), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n453), .B1(new_n696), .B2(new_n455), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n689), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n432), .A2(new_n433), .A3(new_n430), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT75), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n434), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n702), .A2(new_n446), .B1(new_n450), .B2(new_n445), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  AOI22_X1  g503(.A1(new_n436), .A2(KEYINPUT35), .B1(new_n440), .B2(new_n442), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT105), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n444), .A2(new_n497), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n620), .A2(KEYINPUT44), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT106), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n706), .A2(new_n712), .A3(new_n708), .A4(new_n709), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n688), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n555), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n582), .A2(new_n715), .A3(new_n643), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n714), .A2(new_n441), .A3(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n679), .B(new_n681), .C1(new_n503), .C2(new_n717), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n714), .A2(new_n392), .A3(new_n716), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n714), .A2(KEYINPUT107), .A3(new_n392), .A4(new_n716), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(G36gat), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n455), .A2(G36gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n675), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n675), .A2(new_n727), .A3(new_n724), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n723), .A2(new_n726), .A3(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(G43gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n674), .B2(new_n450), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n714), .A2(G43gat), .A3(new_n703), .A4(new_n716), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT47), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(new_n735), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1330gat));
  INV_X1    g536(.A(G50gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n674), .B2(new_n453), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n714), .A2(G50gat), .A3(new_n249), .A4(new_n716), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT48), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n739), .A2(new_n743), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1331gat));
  AND2_X1   g544(.A1(new_n706), .A2(new_n708), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n621), .A2(new_n555), .A3(new_n671), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n441), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g550(.A1(new_n455), .A2(KEYINPUT108), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n455), .A2(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n748), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  AND2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n756), .B2(new_n757), .ZN(G1333gat));
  NOR2_X1   g559(.A1(new_n452), .A2(new_n562), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n747), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT109), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n562), .B1(new_n748), .B2(new_n450), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n748), .A2(new_n453), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n563), .ZN(G1335gat));
  NOR3_X1   g569(.A1(new_n582), .A2(new_n555), .A3(new_n671), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n714), .A2(new_n441), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n582), .A2(new_n555), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n682), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n682), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n775), .A2(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n441), .A2(new_n587), .A3(new_n643), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n772), .A2(new_n587), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  NAND3_X1  g583(.A1(new_n714), .A2(new_n754), .A3(new_n771), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n754), .A2(new_n588), .A3(new_n643), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT112), .Z(new_n788));
  NAND2_X1  g587(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n714), .A2(new_n392), .A3(new_n771), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G92gat), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n780), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n775), .A2(KEYINPUT114), .A3(new_n776), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n788), .B(KEYINPUT113), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n791), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n790), .A2(new_n791), .B1(new_n793), .B2(new_n799), .ZN(G1337gat));
  NAND3_X1  g599(.A1(new_n714), .A2(new_n703), .A3(new_n771), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G99gat), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n450), .A2(G99gat), .A3(new_n671), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n782), .B2(new_n803), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n714), .A2(new_n249), .A3(new_n771), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G106gat), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n671), .A2(G106gat), .A3(new_n453), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n781), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n805), .A2(G106gat), .B1(new_n797), .B2(new_n808), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(G1339gat));
  NOR3_X1   g612(.A1(new_n541), .A2(new_n542), .A3(new_n540), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n529), .B1(new_n528), .B2(new_n534), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n550), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n554), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n618), .A2(new_n619), .A3(new_n817), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n630), .A2(new_n622), .A3(new_n632), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n633), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n622), .C1(new_n630), .C2(new_n632), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n640), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT116), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n820), .A2(new_n823), .A3(KEYINPUT55), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(new_n642), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n824), .A2(new_n830), .A3(new_n825), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n818), .A2(new_n832), .A3(KEYINPUT117), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n643), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n832), .B2(new_n715), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n620), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT117), .B1(new_n818), .B2(new_n832), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n838), .A2(new_n669), .B1(new_n715), .B2(new_n644), .ZN(new_n839));
  INV_X1    g638(.A(new_n440), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n754), .A2(new_n454), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(new_n295), .A3(new_n715), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n839), .A2(new_n454), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n702), .A2(new_n373), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(new_n755), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n555), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n844), .B1(new_n849), .B2(new_n295), .ZN(G1340gat));
  NOR3_X1   g649(.A1(new_n843), .A2(new_n293), .A3(new_n671), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n643), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n293), .ZN(G1341gat));
  NOR2_X1   g652(.A1(new_n669), .A2(G127gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n755), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n843), .A2(new_n669), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n305), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n855), .B(KEYINPUT118), .C1(new_n305), .C2(new_n856), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1342gat));
  NOR2_X1   g660(.A1(new_n620), .A2(new_n392), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n326), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n843), .B2(new_n620), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  NAND2_X1  g666(.A1(new_n842), .A2(new_n452), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n839), .B2(new_n453), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n833), .A2(new_n837), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n828), .A2(new_n642), .ZN(new_n872));
  XNOR2_X1  g671(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(new_n820), .B2(new_n823), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT120), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n824), .A2(new_n873), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n877), .A2(new_n878), .A3(new_n642), .A4(new_n828), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n555), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n670), .B1(new_n880), .B2(new_n834), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n669), .B1(new_n871), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n644), .A2(new_n715), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n453), .A2(new_n869), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n868), .B1(new_n870), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n216), .B1(new_n887), .B2(new_n555), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n838), .A2(new_n669), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n883), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n703), .A2(new_n453), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n441), .A3(new_n891), .ZN(new_n892));
  NOR4_X1   g691(.A1(new_n892), .A2(G141gat), .A3(new_n715), .A4(new_n754), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT58), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n845), .A2(KEYINPUT121), .A3(new_n891), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n715), .A2(G141gat), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n896), .A2(new_n897), .A3(new_n755), .A4(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  AOI211_X1 g699(.A(new_n715), .B(new_n868), .C1(new_n870), .C2(new_n886), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n899), .B(new_n900), .C1(new_n901), .C2(new_n216), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n894), .A2(new_n902), .ZN(G1344gat));
  NAND2_X1  g702(.A1(new_n890), .A2(new_n885), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n818), .A2(new_n832), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n880), .A2(new_n834), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n905), .B(new_n907), .C1(new_n908), .C2(new_n670), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT122), .B1(new_n881), .B2(new_n906), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(new_n669), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n453), .B1(new_n911), .B2(new_n883), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n904), .B1(new_n912), .B2(KEYINPUT57), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n913), .A2(new_n452), .A3(new_n643), .A4(new_n842), .ZN(new_n914));
  AND2_X1   g713(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n671), .A2(KEYINPUT59), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n914), .A2(new_n915), .B1(new_n887), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n896), .A2(new_n897), .A3(new_n643), .A4(new_n755), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(KEYINPUT59), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n919), .B2(G148gat), .ZN(G1345gat));
  NAND4_X1  g719(.A1(new_n896), .A2(new_n897), .A3(new_n582), .A4(new_n755), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n582), .A2(G155gat), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT123), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n921), .A2(new_n231), .B1(new_n887), .B2(new_n923), .ZN(G1346gat));
  NAND4_X1  g723(.A1(new_n896), .A2(new_n897), .A3(new_n232), .A4(new_n862), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n887), .A2(new_n670), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n232), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n441), .A2(new_n455), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n841), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n715), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n846), .A2(new_n754), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n839), .A2(new_n441), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n273), .A3(new_n555), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(new_n933), .ZN(G1348gat));
  OAI21_X1  g733(.A(G176gat), .B1(new_n929), .B2(new_n671), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(new_n262), .A3(new_n643), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1349gat));
  NAND4_X1  g736(.A1(new_n890), .A2(new_n440), .A3(new_n582), .A4(new_n928), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n841), .A2(KEYINPUT124), .A3(new_n582), .A4(new_n928), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n941), .A3(G183gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n932), .A2(new_n270), .A3(new_n582), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT60), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n256), .A3(new_n670), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT125), .ZN(new_n950));
  OAI21_X1  g749(.A(G190gat), .B1(new_n929), .B2(new_n620), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(G1351gat));
  NAND2_X1  g754(.A1(new_n891), .A2(new_n754), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n839), .A2(new_n441), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(G197gat), .B1(new_n957), .B2(new_n555), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n452), .A2(new_n928), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n913), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n555), .A2(G197gat), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(G1352gat));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  AOI21_X1  g763(.A(G204gat), .B1(new_n964), .B2(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n957), .A2(new_n643), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n961), .A2(new_n643), .ZN(new_n969));
  INV_X1    g768(.A(G204gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n957), .A2(new_n204), .A3(new_n582), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n913), .A2(new_n582), .A3(new_n960), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  NAND3_X1  g775(.A1(new_n957), .A2(new_n205), .A3(new_n670), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n961), .A2(new_n670), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n205), .ZN(G1355gat));
endmodule


