//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND3_X1  g0008(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n202), .A2(G50), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G116), .ZN(new_n214));
  INV_X1    g0014(.A(G270), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G250), .B(G257), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n229), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G50), .B(G68), .Z(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(G107), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G97), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n220), .A2(G107), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n237), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G1), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G13), .A3(G20), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n248), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  INV_X1    g0053(.A(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n247), .A2(new_n259), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n245), .A2(G20), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G68), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n250), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT11), .B1(new_n256), .B2(new_n259), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT14), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  OAI211_X1 g0070(.A(G1), .B(G13), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G274), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n258), .B1(G33), .B2(G41), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(new_n273), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G238), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT65), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n280), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT65), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G226), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G97), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n279), .B1(new_n293), .B2(new_n275), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI211_X1 g0096(.A(KEYINPUT13), .B(new_n279), .C1(new_n293), .C2(new_n275), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n268), .B(G169), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n295), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n289), .B1(new_n283), .B2(new_n287), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n300), .A2(G232), .B1(G33), .B2(G97), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n271), .B1(new_n301), .B2(new_n290), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT13), .B1(new_n302), .B2(new_n279), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(new_n303), .A3(G179), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n299), .A2(new_n303), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n268), .B1(new_n306), .B2(G169), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n267), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n259), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n246), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n262), .A2(G50), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n310), .A2(new_n311), .B1(G50), .B2(new_n246), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT67), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n312), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  INV_X1    g0115(.A(G150), .ZN(new_n316));
  INV_X1    g0116(.A(new_n251), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n315), .A2(new_n255), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n254), .B1(new_n201), .B2(new_n212), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n259), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT9), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n314), .A2(KEYINPUT9), .A3(new_n320), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n274), .B1(new_n277), .B2(new_n213), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n288), .A2(G222), .A3(new_n289), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n288), .A2(G1698), .ZN(new_n328));
  XOR2_X1   g0128(.A(KEYINPUT66), .B(G223), .Z(new_n329));
  OAI221_X1 g0129(.A(new_n327), .B1(new_n253), .B2(new_n288), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n330), .B2(new_n275), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(G190), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT10), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n323), .A2(new_n324), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT10), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n331), .A2(new_n325), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n333), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G244), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n274), .B1(new_n277), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n288), .A2(G232), .A3(new_n289), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n343), .B1(new_n238), .B2(new_n288), .C1(new_n328), .C2(new_n278), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n344), .B2(new_n275), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n261), .A2(G77), .A3(new_n262), .ZN(new_n348));
  XOR2_X1   g0148(.A(new_n348), .B(KEYINPUT68), .Z(new_n349));
  NAND2_X1  g0149(.A1(new_n247), .A2(new_n253), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n315), .A2(new_n317), .B1(new_n254), .B2(new_n253), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT15), .B(G87), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n255), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n259), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n347), .B(new_n355), .C1(G169), .C2(new_n345), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n345), .A2(G190), .ZN(new_n357));
  INV_X1    g0157(.A(new_n355), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n357), .B(new_n358), .C1(new_n325), .C2(new_n345), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n331), .A2(new_n346), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(new_n321), .C1(G169), .C2(new_n331), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n356), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(G200), .B1(new_n296), .B2(new_n297), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n299), .A2(new_n303), .A3(G190), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n266), .A3(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n308), .A2(new_n340), .A3(new_n362), .A4(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n274), .B1(new_n277), .B2(new_n219), .ZN(new_n367));
  NOR2_X1   g0167(.A1(G223), .A2(G1698), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n213), .B2(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT69), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n280), .ZN(new_n371));
  NAND2_X1  g0171(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(G33), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(new_n373), .A3(new_n284), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT71), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n271), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(KEYINPUT71), .A3(new_n375), .ZN(new_n379));
  AOI211_X1 g0179(.A(G179), .B(new_n367), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(new_n377), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(new_n379), .A3(new_n275), .ZN(new_n382));
  INV_X1    g0182(.A(new_n367), .ZN(new_n383));
  AOI21_X1  g0183(.A(G169), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT72), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G169), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n374), .A2(KEYINPUT71), .A3(new_n375), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT71), .B1(new_n374), .B2(new_n375), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n387), .A2(new_n388), .A3(new_n271), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n386), .B1(new_n389), .B2(new_n367), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT72), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n382), .A2(new_n346), .A3(new_n383), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n385), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n315), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n262), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n396), .A2(new_n310), .B1(new_n246), .B2(new_n395), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n283), .A2(new_n254), .A3(new_n287), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT70), .ZN(new_n402));
  AND2_X1   g0202(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n403));
  NOR2_X1   g0203(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n269), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n285), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n254), .A2(KEYINPUT7), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n402), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  AOI211_X1 g0209(.A(KEYINPUT70), .B(new_n407), .C1(new_n405), .C2(new_n285), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n401), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G68), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n218), .A2(new_n248), .ZN(new_n413));
  OAI21_X1  g0213(.A(G20), .B1(new_n413), .B2(new_n201), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n251), .A2(G159), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT16), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n403), .A2(new_n404), .A3(new_n269), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n400), .B(new_n254), .C1(new_n419), .C2(new_n281), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(G20), .B1(new_n373), .B2(new_n284), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n400), .ZN(new_n423));
  OAI211_X1 g0223(.A(KEYINPUT16), .B(new_n417), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n259), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n398), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n394), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT18), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n380), .A2(new_n384), .A3(KEYINPUT72), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n391), .B1(new_n390), .B2(new_n392), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n429), .B(new_n426), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n371), .A2(new_n372), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n282), .B1(new_n433), .B2(new_n269), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT70), .B1(new_n434), .B2(new_n407), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n406), .A2(new_n402), .A3(new_n408), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n435), .A2(new_n436), .B1(new_n400), .B2(new_n399), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n417), .B1(new_n437), .B2(new_n248), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT16), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n248), .B1(new_n422), .B2(new_n400), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n403), .A2(new_n404), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n281), .B1(new_n442), .B2(G33), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT7), .B1(new_n443), .B2(G20), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n416), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n309), .B1(new_n445), .B2(KEYINPUT16), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n397), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G200), .B1(new_n389), .B2(new_n367), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n382), .A2(G190), .A3(new_n383), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(KEYINPUT73), .A2(KEYINPUT17), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT73), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n447), .A2(new_n450), .A3(new_n451), .A4(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n416), .B1(new_n411), .B2(G68), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n446), .B1(new_n456), .B2(KEYINPUT16), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(new_n398), .A3(new_n449), .A4(new_n448), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(new_n452), .A3(new_n453), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n428), .A2(new_n432), .A3(new_n455), .A4(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n366), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n272), .A2(G1), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT5), .B(G41), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n275), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G264), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n464), .A2(new_n271), .A3(G274), .A4(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n373), .A2(new_n284), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n289), .A2(G250), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT87), .B(G294), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n468), .A2(new_n469), .B1(new_n269), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n221), .A2(new_n289), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n373), .A2(new_n284), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT86), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n443), .A2(KEYINPUT86), .A3(new_n472), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n466), .B(new_n467), .C1(new_n477), .C2(new_n271), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n325), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n476), .A2(new_n475), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n275), .B1(new_n480), .B2(new_n471), .ZN(new_n481));
  INV_X1    g0281(.A(G190), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(new_n466), .A4(new_n467), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT25), .B1(new_n247), .B2(new_n238), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT85), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n238), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT84), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n245), .A2(G33), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT74), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n261), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n486), .A2(new_n488), .B1(new_n238), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT83), .ZN(new_n494));
  INV_X1    g0294(.A(G87), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n495), .A2(KEYINPUT22), .A3(G20), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n288), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n373), .A2(new_n254), .A3(G87), .A4(new_n284), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT22), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT23), .B1(new_n254), .B2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT23), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(new_n238), .A3(G20), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n501), .B(new_n503), .C1(new_n214), .C2(new_n255), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT82), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n494), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT24), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n309), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n288), .A2(new_n496), .B1(new_n498), .B2(KEYINPUT22), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n504), .B(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT83), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n500), .A2(new_n494), .A3(new_n505), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(KEYINPUT24), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n493), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n484), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n478), .A2(new_n386), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n481), .A2(new_n346), .A3(new_n466), .A4(new_n467), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n515), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT88), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n484), .A2(new_n515), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT88), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n522), .B(new_n523), .C1(new_n515), .C2(new_n519), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n443), .A2(new_n254), .A3(G68), .ZN(new_n526));
  OR2_X1    g0326(.A1(KEYINPUT79), .A2(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(KEYINPUT79), .A2(G87), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n527), .A2(new_n220), .A3(new_n238), .A4(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n292), .B2(new_n254), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n254), .A2(G33), .A3(G97), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n529), .A2(new_n531), .B1(new_n532), .B2(new_n530), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n259), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n352), .A2(new_n247), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n489), .B(KEYINPUT74), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n310), .ZN(new_n539));
  INV_X1    g0339(.A(new_n352), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n541), .B(KEYINPUT80), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n271), .B(G250), .C1(G1), .C2(new_n272), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n271), .A2(G274), .A3(new_n463), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT77), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT77), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n289), .A2(G238), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n468), .A2(new_n550), .B1(new_n269), .B2(new_n214), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT78), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n443), .A2(new_n552), .A3(G244), .A4(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n373), .A2(G244), .A3(G1698), .A4(new_n284), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT78), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n549), .B1(new_n556), .B2(new_n271), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n537), .A2(new_n542), .B1(new_n557), .B2(new_n386), .ZN(new_n558));
  INV_X1    g0358(.A(new_n557), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n346), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n539), .A2(G87), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n535), .A2(new_n536), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n557), .B2(G200), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT81), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n557), .B2(new_n482), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n553), .A2(new_n555), .ZN(new_n567));
  INV_X1    g0367(.A(new_n551), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n275), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n570), .A2(KEYINPUT81), .A3(G190), .A4(new_n549), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n564), .A2(new_n566), .A3(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n247), .A2(new_n214), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n492), .B2(new_n214), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G283), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n577), .B(new_n254), .C1(G33), .C2(new_n220), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n214), .A2(G20), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n259), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n580), .B(KEYINPUT20), .ZN(new_n581));
  OAI21_X1  g0381(.A(G169), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  MUX2_X1   g0382(.A(G257), .B(G264), .S(G1698), .Z(new_n583));
  NAND2_X1  g0383(.A1(new_n443), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n283), .A2(G303), .A3(new_n287), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n271), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n465), .A2(G270), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n467), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n574), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(G190), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n576), .A2(new_n581), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(new_n325), .C2(new_n589), .ZN(new_n593));
  INV_X1    g0393(.A(new_n589), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n576), .A2(new_n581), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT21), .A4(G169), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n589), .A3(G179), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n590), .A2(new_n593), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n437), .A2(new_n238), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n239), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g0401(.A(G97), .B(G107), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n603), .A2(new_n254), .B1(new_n253), .B2(new_n317), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n259), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n246), .A2(G97), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n539), .B2(G97), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT75), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n464), .A2(new_n463), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(G257), .A3(new_n271), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n608), .B1(new_n610), .B2(new_n467), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n610), .A2(new_n608), .A3(new_n467), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT4), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(new_n341), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n288), .A2(new_n289), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n287), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n286), .B1(new_n284), .B2(new_n285), .ZN(new_n617));
  OAI211_X1 g0417(.A(G250), .B(G1698), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n373), .A2(G244), .A3(new_n289), .A4(new_n284), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n613), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n615), .A2(new_n618), .A3(new_n620), .A4(new_n577), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n611), .B(new_n612), .C1(new_n621), .C2(new_n275), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n605), .A2(new_n607), .B1(new_n622), .B2(new_n346), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n275), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT76), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n612), .A2(new_n611), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n624), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n386), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n604), .B1(new_n411), .B2(G107), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n607), .B1(new_n631), .B2(new_n309), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n624), .A2(new_n626), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n632), .B1(G200), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT76), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(G190), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n573), .A2(new_n598), .A3(new_n630), .A4(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n462), .A2(new_n525), .A3(new_n639), .ZN(G372));
  INV_X1    g0440(.A(new_n361), .ZN(new_n641));
  INV_X1    g0441(.A(new_n432), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n429), .B1(new_n394), .B2(new_n426), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n459), .A2(new_n455), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n365), .ZN(new_n646));
  INV_X1    g0446(.A(new_n356), .ZN(new_n647));
  OAI21_X1  g0447(.A(G169), .B1(new_n296), .B2(new_n297), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n304), .A3(new_n298), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n647), .B1(new_n650), .B2(new_n267), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n644), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n340), .B(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n641), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n596), .A2(new_n590), .A3(new_n597), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n515), .B2(new_n519), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n559), .A2(G190), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n484), .A2(new_n515), .B1(new_n658), .B2(new_n564), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n657), .A2(new_n638), .A3(new_n659), .A4(new_n630), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(new_n561), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n561), .A2(new_n572), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n630), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n658), .A2(new_n564), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n561), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n665), .B1(new_n667), .B2(new_n630), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n461), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n655), .A2(new_n671), .ZN(G369));
  NAND3_X1  g0472(.A1(new_n245), .A2(new_n254), .A3(G13), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  INV_X1    g0475(.A(G213), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G343), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT90), .Z(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n595), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n598), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n656), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n679), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n521), .B(new_n524), .C1(new_n515), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n520), .A2(new_n679), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n520), .A2(new_n685), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n656), .A2(new_n679), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n521), .A2(new_n524), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n206), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n529), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n210), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n663), .A2(new_n665), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT26), .B1(new_n667), .B2(new_n630), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n561), .A3(new_n660), .A4(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .A3(new_n685), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n679), .B1(new_n661), .B2(new_n669), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n466), .B1(new_n477), .B2(new_n271), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n584), .A2(new_n585), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n275), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(G179), .A3(new_n467), .A4(new_n587), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n635), .A2(new_n712), .A3(new_n559), .A4(new_n636), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n708), .A2(new_n557), .A3(new_n711), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(KEYINPUT30), .A3(new_n635), .A4(new_n636), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n589), .A2(G179), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n633), .A2(new_n718), .A3(new_n478), .A4(new_n557), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT31), .B1(new_n720), .B2(new_n679), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n638), .A2(new_n598), .A3(new_n630), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n662), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n521), .A3(new_n524), .A4(new_n685), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n707), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n706), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT91), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n706), .A2(new_n728), .A3(KEYINPUT91), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n700), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(G13), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n245), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n695), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n684), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G330), .B2(new_n682), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n258), .B1(G20), .B2(new_n386), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n346), .A2(new_n325), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(new_n254), .A3(G190), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT93), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(KEYINPUT93), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(G159), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(G20), .B1(new_n743), .B2(new_n482), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT95), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G97), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n750), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n254), .A2(G179), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n527), .B2(new_n528), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n254), .A2(new_n346), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n482), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n761), .B1(G50), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n762), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n766), .A2(new_n482), .A3(G200), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G58), .A2(new_n767), .B1(new_n768), .B2(G77), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n763), .A2(G190), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n759), .A2(new_n482), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n770), .A2(G68), .B1(new_n772), .B2(G107), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n765), .A2(new_n769), .A3(new_n288), .A4(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n749), .B1(new_n748), .B2(G159), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n758), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n764), .B(KEYINPUT96), .Z(new_n777));
  INV_X1    g0577(.A(G326), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n777), .A2(new_n778), .B1(new_n470), .B2(new_n755), .ZN(new_n779));
  INV_X1    g0579(.A(G317), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n770), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  INV_X1    g0584(.A(G303), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n783), .B1(new_n784), .B2(new_n771), .C1(new_n785), .C2(new_n760), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G311), .A2(new_n768), .B1(new_n767), .B2(G322), .ZN(new_n787));
  INV_X1    g0587(.A(new_n288), .ZN(new_n788));
  INV_X1    g0588(.A(G329), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(new_n747), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n779), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n742), .B1(new_n776), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n742), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n237), .A2(new_n272), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n210), .A2(G45), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n468), .A2(new_n206), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n288), .A2(new_n206), .ZN(new_n801));
  XOR2_X1   g0601(.A(G355), .B(KEYINPUT92), .Z(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n802), .B1(G116), .B2(new_n206), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n796), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n792), .A2(new_n804), .A3(new_n739), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT97), .ZN(new_n806));
  INV_X1    g0606(.A(new_n795), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n682), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n741), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  OAI21_X1  g0610(.A(new_n359), .B1(new_n358), .B2(new_n685), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n356), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n647), .A2(new_n685), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n705), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n662), .A2(new_n630), .A3(new_n665), .ZN(new_n817));
  AOI21_X1  g0617(.A(G169), .B1(new_n635), .B2(new_n636), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n632), .B1(G179), .B2(new_n633), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n560), .A2(new_n558), .B1(new_n658), .B2(new_n564), .ZN(new_n821));
  AOI21_X1  g0621(.A(KEYINPUT26), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n660), .A2(new_n561), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n815), .B(new_n685), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n728), .B1(new_n816), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(KEYINPUT100), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(KEYINPUT100), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n816), .A2(new_n826), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n739), .B1(new_n830), .B2(new_n727), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n739), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n742), .A2(new_n793), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n253), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n742), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n495), .A2(new_n771), .B1(new_n760), .B2(new_n238), .ZN(new_n837));
  INV_X1    g0637(.A(G294), .ZN(new_n838));
  INV_X1    g0638(.A(new_n767), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n788), .B1(new_n838), .B2(new_n839), .C1(new_n747), .C2(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n837), .B(new_n841), .C1(G303), .C2(new_n764), .ZN(new_n842));
  INV_X1    g0642(.A(new_n768), .ZN(new_n843));
  INV_X1    g0643(.A(new_n770), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n843), .A2(new_n214), .B1(new_n844), .B2(new_n784), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n757), .B1(KEYINPUT98), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(KEYINPUT98), .B2(new_n845), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G143), .A2(new_n767), .B1(new_n768), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  INV_X1    g0649(.A(new_n764), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n848), .B1(new_n849), .B2(new_n850), .C1(new_n316), .C2(new_n844), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT34), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n443), .B1(new_n747), .B2(new_n853), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n212), .A2(new_n760), .B1(new_n771), .B2(new_n248), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT99), .Z(new_n856));
  AOI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(G58), .C2(new_n756), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n842), .A2(new_n847), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n835), .B1(new_n836), .B2(new_n858), .C1(new_n815), .C2(new_n794), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n832), .A2(new_n859), .ZN(G384));
  NOR2_X1   g0660(.A1(new_n736), .A2(new_n245), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n704), .B(new_n461), .C1(new_n705), .C2(KEYINPUT29), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n655), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT107), .Z(new_n864));
  INV_X1    g0664(.A(new_n365), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n267), .B(new_n679), .C1(new_n650), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n267), .A2(new_n679), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n308), .A2(new_n365), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n825), .B2(new_n813), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n426), .A2(new_n677), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n458), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n385), .A2(new_n393), .B1(new_n457), .B2(new_n398), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n874), .A2(KEYINPUT37), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n417), .B1(new_n421), .B2(new_n423), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT16), .B1(new_n877), .B2(KEYINPUT103), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT103), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n445), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n425), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT104), .B1(new_n881), .B2(new_n397), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n439), .B1(new_n445), .B2(new_n879), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n877), .A2(KEYINPUT103), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n446), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n398), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n882), .A2(new_n677), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n882), .A2(new_n394), .A3(new_n887), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n458), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n876), .B1(KEYINPUT37), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n888), .B1(new_n644), .B2(new_n645), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n872), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(new_n876), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n888), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n460), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n893), .A2(new_n899), .A3(KEYINPUT105), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT105), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n872), .C1(new_n891), .C2(new_n892), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n871), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n644), .A2(new_n677), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n895), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n873), .B1(new_n644), .B2(new_n645), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT39), .B1(new_n910), .B2(new_n899), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n900), .A2(new_n902), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n911), .B1(new_n912), .B2(KEYINPUT39), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n650), .A2(new_n267), .A3(new_n685), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n905), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n864), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n869), .A2(new_n815), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n726), .B2(new_n723), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n900), .A2(new_n919), .A3(new_n902), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n910), .A2(new_n899), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n720), .A2(new_n679), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT31), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n525), .A2(new_n639), .A3(new_n679), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n929), .A2(new_n921), .A3(new_n918), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n920), .A2(new_n921), .B1(new_n922), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(new_n462), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n707), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n931), .B2(new_n932), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n861), .B1(new_n917), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n917), .B2(new_n934), .ZN(new_n936));
  INV_X1    g0736(.A(new_n603), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n214), .B(new_n209), .C1(new_n937), .C2(KEYINPUT35), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(KEYINPUT35), .B2(new_n937), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT36), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n210), .A2(new_n253), .A3(new_n413), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n941), .A2(KEYINPUT101), .B1(new_n212), .B2(G68), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(KEYINPUT101), .B2(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n735), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT102), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n936), .A2(new_n946), .ZN(G367));
  NAND2_X1  g0747(.A1(new_n632), .A2(new_n679), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n638), .A2(new_n630), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n820), .A2(new_n679), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(new_n692), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(KEYINPUT42), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n638), .A2(new_n520), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n679), .B1(new_n954), .B2(new_n630), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n952), .B2(KEYINPUT42), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n679), .A2(new_n563), .ZN(new_n958));
  MUX2_X1   g0758(.A(new_n561), .B(new_n667), .S(new_n958), .Z(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT108), .Z(new_n960));
  INV_X1    g0760(.A(KEYINPUT43), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n957), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n953), .A2(new_n956), .A3(new_n961), .A4(new_n960), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n689), .A2(new_n951), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n695), .B(KEYINPUT41), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n692), .A2(new_n690), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT109), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n970), .A2(new_n971), .A3(new_n951), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n971), .B1(new_n970), .B2(new_n951), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT44), .ZN(new_n975));
  INV_X1    g0775(.A(new_n951), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n690), .A3(new_n692), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n972), .B2(new_n973), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n975), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n689), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n692), .B1(new_n688), .B2(new_n691), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n987), .A2(new_n684), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n684), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n975), .A2(new_n981), .A3(new_n689), .A4(new_n983), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n986), .A2(new_n991), .A3(new_n733), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n969), .B1(new_n993), .B2(new_n733), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n968), .B1(new_n994), .B2(new_n738), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n960), .A2(new_n795), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n229), .A2(new_n799), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n796), .B1(new_n206), .B2(new_n352), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n739), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n777), .A2(new_n840), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n760), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT46), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n760), .B2(new_n214), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(new_n747), .C2(new_n780), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G283), .A2(new_n768), .B1(new_n767), .B2(G303), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n771), .A2(new_n220), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n470), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n770), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1006), .A2(new_n468), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n755), .A2(new_n238), .ZN(new_n1011));
  NOR4_X1   g0811(.A1(new_n1000), .A2(new_n1005), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(G143), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n777), .A2(new_n1013), .B1(new_n248), .B2(new_n755), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n771), .A2(new_n253), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G159), .B2(new_n770), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n218), .B2(new_n760), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G50), .A2(new_n768), .B1(new_n767), .B2(G150), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1018), .B(new_n288), .C1(new_n849), .C2(new_n747), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1014), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1012), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT110), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT47), .Z(new_n1023));
  AOI21_X1  g0823(.A(new_n999), .B1(new_n1023), .B2(new_n742), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n996), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT111), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n995), .A2(new_n1027), .ZN(G387));
  INV_X1    g0828(.A(KEYINPUT115), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n991), .A2(KEYINPUT112), .A3(new_n738), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT112), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n990), .B2(new_n737), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n686), .A2(new_n687), .A3(new_n795), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G303), .A2(new_n768), .B1(new_n767), .B2(G317), .ZN(new_n1034));
  INV_X1    g0834(.A(G322), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1034), .B1(new_n840), .B2(new_n844), .C1(new_n777), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n756), .A2(G283), .B1(new_n1008), .B2(new_n1001), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT49), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n468), .B1(new_n214), .B2(new_n771), .C1(new_n747), .C2(new_n778), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT114), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(G159), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1048), .A2(new_n850), .B1(new_n844), .B2(new_n315), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1007), .B(new_n1049), .C1(G77), .C2(new_n1001), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n443), .B1(new_n843), .B2(new_n248), .C1(new_n212), .C2(new_n839), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G150), .B2(new_n748), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n756), .A2(new_n540), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT113), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n836), .B1(new_n1047), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n233), .A2(new_n272), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1057), .A2(new_n799), .B1(new_n697), .B2(new_n801), .ZN(new_n1058));
  OR3_X1    g0858(.A1(new_n315), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT50), .B1(new_n315), .B2(G50), .ZN(new_n1060));
  AOI21_X1  g0860(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1059), .A2(new_n697), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(G107), .B2(new_n206), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n833), .B(new_n1056), .C1(new_n796), .C2(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1030), .A2(new_n1032), .B1(new_n1033), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n733), .A2(new_n991), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n731), .A2(new_n732), .A3(new_n990), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n695), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1029), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1066), .A2(new_n1069), .A3(new_n1029), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(G393));
  INV_X1    g0873(.A(KEYINPUT116), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n986), .B2(new_n992), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT116), .B1(new_n984), .B2(new_n985), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n951), .A2(new_n795), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n796), .B1(new_n220), .B2(new_n206), .C1(new_n243), .C2(new_n799), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n739), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n747), .A2(new_n1013), .B1(new_n248), .B2(new_n760), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT117), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n443), .B1(new_n495), .B2(new_n771), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT118), .Z(new_n1085));
  AOI22_X1  g0885(.A1(new_n767), .A2(G159), .B1(new_n764), .B2(G150), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT51), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n755), .A2(new_n253), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n843), .A2(new_n315), .B1(new_n844), .B2(new_n212), .ZN(new_n1089));
  OR3_X1    g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n767), .A2(G311), .B1(new_n764), .B2(G317), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT52), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n788), .B1(new_n843), .B2(new_n838), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n748), .B2(G322), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n844), .A2(new_n785), .B1(new_n771), .B2(new_n238), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G283), .B2(new_n1001), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(new_n214), .C2(new_n755), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1085), .A2(new_n1090), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1080), .B1(new_n1098), .B2(new_n742), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1077), .A2(new_n738), .B1(new_n1078), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1067), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n695), .A3(new_n993), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(G390));
  OAI211_X1 g0903(.A(new_n461), .B(G330), .C1(new_n927), .C2(new_n928), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n862), .A2(new_n655), .A3(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(G330), .B(new_n815), .C1(new_n927), .C2(new_n928), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n870), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n727), .A2(new_n815), .A3(new_n869), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n813), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n703), .A2(new_n685), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n812), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n705), .B2(new_n812), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1105), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n914), .B1(new_n1113), .B2(new_n870), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT39), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n900), .B2(new_n902), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1118), .B2(new_n911), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n914), .B(KEYINPUT119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n922), .B(new_n1120), .C1(new_n1111), .C2(new_n870), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1119), .A2(new_n1108), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1108), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1115), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1106), .A2(new_n870), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1119), .A2(new_n1108), .A3(new_n1121), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n862), .A2(new_n655), .A3(new_n1104), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1113), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n869), .B1(new_n727), .B2(new_n815), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1107), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1127), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1124), .A2(new_n1135), .A3(new_n695), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n738), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n913), .A2(new_n794), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n767), .A2(G132), .B1(new_n764), .B2(G128), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT120), .Z(new_n1141));
  OR3_X1    g0941(.A1(new_n760), .A2(KEYINPUT53), .A3(new_n316), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT53), .B1(new_n760), .B2(new_n316), .ZN(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1142), .B(new_n1143), .C1(new_n747), .C2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n788), .B1(new_n768), .B2(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n770), .A2(G137), .B1(new_n772), .B2(G50), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n1048), .C2(new_n755), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1141), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G97), .A2(new_n768), .B1(new_n767), .B2(G116), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1152), .B(new_n788), .C1(new_n838), .C2(new_n747), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n248), .A2(new_n771), .B1(new_n760), .B2(new_n495), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n238), .A2(new_n844), .B1(new_n850), .B2(new_n784), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1153), .A2(new_n1088), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n742), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n833), .B1(new_n315), .B2(new_n834), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1139), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1136), .A2(new_n1138), .A3(new_n1160), .ZN(G378));
  NAND2_X1  g0961(.A1(new_n913), .A2(new_n915), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n903), .A3(new_n904), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n654), .A2(new_n361), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n321), .A2(new_n677), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n654), .A2(new_n361), .A3(new_n1165), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1167), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n920), .A2(new_n921), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n707), .B1(new_n930), .B2(new_n922), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1163), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n916), .A3(new_n1177), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1182), .A2(new_n793), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n834), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n739), .B1(new_n1187), .B2(G50), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n468), .A2(new_n270), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n238), .A2(new_n839), .B1(new_n843), .B2(new_n352), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(G77), .C2(new_n1001), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n771), .A2(new_n218), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n220), .A2(new_n844), .B1(new_n850), .B2(new_n214), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n756), .C2(G68), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1191), .B(new_n1194), .C1(new_n784), .C2(new_n747), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT58), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G50), .B1(new_n269), .B2(new_n270), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1195), .A2(new_n1196), .B1(new_n1189), .B2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n767), .A2(G128), .B1(new_n764), .B2(G125), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n760), .B2(new_n1146), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G137), .A2(new_n768), .B1(new_n770), .B2(G132), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT121), .Z(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G150), .C2(new_n756), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n269), .B(new_n270), .C1(new_n771), .C2(new_n1048), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n748), .B2(G124), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT59), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1207), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1198), .B1(new_n1196), .B2(new_n1195), .C1(new_n1205), .C2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1188), .B1(new_n1210), .B2(new_n742), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1185), .A2(new_n738), .B1(new_n1186), .B2(new_n1211), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1183), .A2(new_n916), .A3(new_n1177), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n916), .B1(new_n1183), .B2(new_n1177), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1129), .B1(new_n1137), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n695), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1135), .A2(new_n1105), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT57), .B1(new_n1219), .B2(new_n1185), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1212), .B1(new_n1218), .B2(new_n1220), .ZN(G375));
  NAND3_X1  g1021(.A1(new_n1132), .A2(new_n1129), .A3(new_n1133), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n969), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1115), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n870), .A2(new_n793), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n739), .B1(new_n1187), .B2(G68), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n214), .A2(new_n844), .B1(new_n850), .B2(new_n838), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1015), .B(new_n1227), .C1(G97), .C2(new_n1001), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n748), .A2(G303), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n839), .A2(new_n784), .B1(new_n843), .B2(new_n238), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(new_n288), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1053), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n748), .A2(G128), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n756), .A2(G50), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n468), .B1(new_n768), .B2(G150), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1192), .B1(G159), .B2(new_n1001), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G137), .A2(new_n767), .B1(new_n770), .B2(new_n1147), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n853), .B2(new_n850), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT122), .Z(new_n1240));
  OAI21_X1  g1040(.A(new_n1232), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT123), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n836), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1226), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1216), .A2(new_n738), .B1(new_n1225), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1224), .A2(new_n1246), .ZN(G381));
  NAND3_X1  g1047(.A1(new_n1071), .A2(new_n809), .A3(new_n1072), .ZN(new_n1248));
  OR2_X1    g1048(.A1(G381), .A2(G384), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(G387), .A2(new_n1248), .A3(G390), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G378), .ZN(new_n1251));
  INV_X1    g1051(.A(G375), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(G407));
  NOR2_X1   g1053(.A1(new_n676), .A2(G343), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1251), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(G213), .A3(new_n1255), .ZN(G409));
  NAND2_X1  g1056(.A1(new_n1254), .A2(KEYINPUT125), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1216), .A2(new_n738), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1225), .A2(new_n1245), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1112), .A2(new_n1114), .A3(new_n1105), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT60), .B1(new_n1261), .B2(new_n1134), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n696), .B1(new_n1222), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1260), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT124), .B1(new_n832), .B2(new_n859), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n832), .A2(KEYINPUT124), .A3(new_n859), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1222), .A2(new_n1263), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n695), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1263), .B1(new_n1115), .B2(new_n1222), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1246), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1266), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1267), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1257), .B1(new_n1269), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1254), .A2(G2897), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1277), .B(new_n1257), .C1(new_n1269), .C2(new_n1275), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1212), .C1(new_n1218), .C2(new_n1220), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1219), .A2(new_n1185), .A3(new_n1223), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1212), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1251), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1254), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1072), .ZN(new_n1294));
  OAI21_X1  g1094(.A(G396), .B1(new_n1294), .B2(new_n1070), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1248), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(G387), .A2(new_n1102), .A3(new_n1100), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(G390), .A2(new_n1027), .A3(new_n995), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT126), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1298), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(G387), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT126), .B1(new_n1302), .B2(G390), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1297), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1302), .A2(G390), .B1(new_n1248), .B2(new_n1295), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n1298), .ZN(new_n1307));
  AND4_X1   g1107(.A1(new_n1305), .A2(new_n1298), .A3(new_n1299), .A4(new_n1296), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1304), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1254), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1292), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(KEYINPUT63), .A3(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1290), .A2(new_n1293), .A3(new_n1309), .A4(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1310), .A2(new_n1314), .A3(new_n1311), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1310), .B2(new_n1281), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1314), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1315), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1313), .B1(new_n1319), .B2(new_n1309), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1251), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1283), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1292), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(new_n1283), .A3(new_n1311), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(new_n1309), .ZN(G402));
endmodule


