//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n187));
  XNOR2_X1  g001(.A(G116), .B(G119), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G101), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n194), .A3(new_n198), .A4(new_n195), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT4), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n201), .A3(G101), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n189), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n195), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n190), .A2(G107), .ZN(new_n205));
  OAI21_X1  g019(.A(G101), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(new_n199), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n188), .A2(KEYINPUT5), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n210), .A2(KEYINPUT5), .A3(G119), .ZN(new_n211));
  INV_X1    g025(.A(G113), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n209), .A2(new_n213), .B1(new_n187), .B2(new_n188), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G110), .B(G122), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n203), .A2(new_n215), .A3(new_n217), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(KEYINPUT6), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT6), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(new_n222), .A3(new_n218), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT65), .A2(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(G143), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  INV_X1    g044(.A(G143), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT64), .A2(G143), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(G146), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n229), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT69), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n229), .A2(new_n234), .A3(new_n239), .A4(new_n236), .ZN(new_n240));
  INV_X1    g054(.A(new_n233), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT64), .A2(G143), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n226), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT65), .A2(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT65), .A2(G146), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n231), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n244), .A2(new_n245), .A3(new_n231), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n249));
  OAI21_X1  g063(.A(G128), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n238), .A2(new_n240), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G125), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G224), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n255), .B(KEYINPUT86), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT0), .B(G128), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(G146), .B1(new_n232), .B2(new_n233), .ZN(new_n259));
  AOI21_X1  g073(.A(G143), .B1(new_n227), .B2(new_n228), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n229), .A2(new_n234), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G125), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n253), .A2(new_n256), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n256), .B1(new_n253), .B2(new_n265), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n224), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n253), .A2(new_n265), .ZN(new_n270));
  OR2_X1    g084(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n256), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n217), .B(KEYINPUT8), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n208), .A2(KEYINPUT87), .A3(new_n214), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n208), .B2(new_n214), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT87), .B1(new_n208), .B2(new_n214), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n256), .A4(new_n265), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n274), .A2(new_n279), .A3(new_n220), .A4(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n269), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G210), .B1(G237), .B2(G902), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT89), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n283), .A2(new_n285), .A3(new_n269), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n269), .A2(new_n283), .A3(KEYINPUT89), .A4(new_n285), .ZN(new_n291));
  OAI21_X1  g105(.A(G214), .B1(G237), .B2(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(G234), .A2(G237), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(G952), .A3(new_n254), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(G902), .A3(G953), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT21), .B(G898), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  INV_X1    g116(.A(G217), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n302), .A2(new_n303), .A3(G953), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G122), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G116), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n210), .A2(G122), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n193), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n308), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G107), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n232), .A2(G128), .A3(new_n233), .ZN(new_n314));
  INV_X1    g128(.A(G134), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n235), .A2(G143), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT13), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n235), .B2(G143), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n241), .A2(new_n242), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(G128), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n314), .A2(new_n319), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT96), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n315), .B1(new_n323), .B2(KEYINPUT96), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n318), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n317), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n310), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT14), .ZN(new_n331));
  OAI21_X1  g145(.A(G107), .B1(new_n308), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT97), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n333), .B(new_n334), .C1(KEYINPUT14), .C2(new_n311), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n311), .A2(KEYINPUT14), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT97), .B1(new_n336), .B2(new_n332), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n330), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n305), .B1(new_n327), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n326), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n317), .B(new_n313), .C1(new_n340), .C2(new_n324), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(new_n337), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(new_n310), .C1(new_n328), .C2(new_n329), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n343), .A3(new_n304), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT98), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT98), .B(new_n305), .C1(new_n327), .C2(new_n338), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n282), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G478), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(KEYINPUT15), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n348), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G131), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(KEYINPUT70), .A2(G237), .ZN(new_n356));
  AOI21_X1  g170(.A(G953), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(G143), .A3(G214), .ZN(new_n358));
  INV_X1    g172(.A(new_n356), .ZN(new_n359));
  NOR2_X1   g173(.A1(KEYINPUT70), .A2(G237), .ZN(new_n360));
  OAI211_X1 g174(.A(G214), .B(new_n254), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n321), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n352), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT17), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT16), .ZN(new_n365));
  INV_X1    g179(.A(G140), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(G125), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n252), .A2(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n367), .B1(new_n370), .B2(new_n365), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(new_n226), .ZN(new_n372));
  XNOR2_X1  g186(.A(G125), .B(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT16), .ZN(new_n374));
  AOI21_X1  g188(.A(G146), .B1(new_n374), .B2(new_n367), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT92), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n226), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(G146), .A3(new_n367), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n364), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n358), .A2(new_n362), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G131), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n358), .A2(new_n362), .A3(new_n352), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT93), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n383), .A2(KEYINPUT93), .A3(new_n384), .A4(new_n385), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n381), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(new_n190), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n227), .A2(new_n228), .ZN(new_n393));
  MUX2_X1   g207(.A(new_n226), .B(new_n393), .S(new_n373), .Z(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n363), .B2(KEYINPUT18), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT18), .A2(G131), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT90), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n358), .A2(new_n362), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n390), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n383), .A2(new_n385), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n370), .B(KEYINPUT19), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n379), .B1(new_n405), .B2(new_n393), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n392), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G475), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n282), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT94), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT20), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n416), .A3(new_n413), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n403), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n392), .B1(new_n390), .B2(new_n402), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT95), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n390), .A2(new_n402), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT95), .A3(new_n408), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n282), .ZN(new_n424));
  OAI21_X1  g238(.A(G475), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n301), .A2(new_n351), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G221), .ZN(new_n428));
  INV_X1    g242(.A(new_n302), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(new_n282), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n238), .A2(new_n240), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n250), .A2(new_n247), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n208), .A2(KEYINPUT10), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n208), .A2(KEYINPUT10), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT82), .B1(new_n251), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G137), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT11), .A3(G134), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n315), .A2(G137), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT66), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(G134), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT11), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI211_X1 g262(.A(KEYINPUT66), .B(KEYINPUT11), .C1(new_n441), .C2(G134), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G131), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n444), .B(new_n352), .C1(new_n448), .C2(new_n449), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n229), .A2(new_n234), .A3(new_n262), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n257), .B1(new_n243), .B2(new_n246), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n202), .A3(new_n200), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n229), .A2(new_n234), .ZN(new_n460));
  OAI21_X1  g274(.A(G128), .B1(new_n259), .B2(new_n249), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n238), .A2(new_n240), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n459), .B1(new_n462), .B2(new_n207), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n440), .A2(new_n454), .A3(new_n458), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT83), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n463), .A2(new_n458), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT83), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n466), .A2(new_n467), .A3(new_n454), .A4(new_n440), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G140), .ZN(new_n470));
  INV_X1    g284(.A(G227), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G953), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n470), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n434), .A2(new_n208), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n462), .A2(new_n207), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n453), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT12), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT12), .B(new_n453), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n469), .A2(new_n474), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n469), .A2(KEYINPUT85), .A3(new_n474), .A4(new_n481), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n466), .A2(new_n440), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n453), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n469), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n473), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G469), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n282), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n282), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI221_X4 g308(.A(KEYINPUT84), .B1(new_n479), .B2(new_n480), .C1(new_n465), .C2(new_n468), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n469), .B2(new_n481), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n473), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n469), .A2(new_n474), .A3(new_n487), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(G469), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n494), .A3(new_n500), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n427), .A2(new_n431), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT80), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n357), .A2(G210), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT26), .B(G101), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT68), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n441), .B2(G134), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n446), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n443), .A2(new_n511), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n452), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n432), .B2(new_n433), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n264), .B1(new_n452), .B2(new_n451), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT73), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n189), .ZN(new_n520));
  INV_X1    g334(.A(new_n452), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n447), .B1(new_n315), .B2(G137), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT66), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n446), .A2(new_n445), .A3(new_n447), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n352), .B1(new_n525), .B2(new_n444), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n457), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT73), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n527), .B(new_n528), .C1(new_n251), .C2(new_n516), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n519), .A2(new_n520), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT28), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n530), .A2(KEYINPUT74), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT74), .B1(new_n530), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n517), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n520), .A3(new_n527), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT67), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n527), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n453), .A2(KEYINPUT67), .A3(new_n457), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n517), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n536), .B1(new_n540), .B2(new_n520), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT28), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n510), .B1(new_n534), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n535), .A2(KEYINPUT30), .A3(new_n527), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n189), .B(new_n544), .C1(new_n540), .C2(KEYINPUT30), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n536), .A3(new_n510), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT31), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n545), .A2(new_n536), .A3(new_n510), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n505), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n530), .A2(new_n531), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT74), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n530), .A2(KEYINPUT74), .A3(new_n531), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n542), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n510), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n558), .A2(KEYINPUT75), .A3(new_n547), .A4(new_n549), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G472), .A2(G902), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT32), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  INV_X1    g377(.A(new_n561), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n563), .B(new_n564), .C1(new_n551), .C2(new_n559), .ZN(new_n565));
  INV_X1    g379(.A(G472), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n189), .B1(new_n517), .B2(new_n518), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n536), .A2(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n533), .B(new_n532), .C1(KEYINPUT28), .C2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n510), .A2(KEYINPUT29), .ZN(new_n570));
  AOI21_X1  g384(.A(G902), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n545), .A2(new_n536), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT29), .B1(new_n572), .B2(new_n557), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n556), .B2(new_n557), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n566), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n562), .A2(new_n565), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT76), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT23), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n580));
  OAI211_X1 g394(.A(G119), .B(new_n235), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G119), .ZN(new_n582));
  OAI22_X1  g396(.A1(new_n577), .A2(new_n578), .B1(new_n582), .B2(G128), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n581), .B(new_n583), .C1(G119), .C2(new_n235), .ZN(new_n584));
  XNOR2_X1  g398(.A(G119), .B(G128), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT24), .B(G110), .Z(new_n586));
  AOI22_X1  g400(.A1(new_n584), .A2(G110), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n377), .A2(new_n379), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT77), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  OAI22_X1  g405(.A1(new_n584), .A2(G110), .B1(new_n585), .B2(new_n586), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n592), .B(new_n379), .C1(new_n393), .C2(new_n370), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT22), .B(G137), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n254), .A2(G221), .A3(G234), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n591), .A2(new_n593), .A3(new_n597), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n303), .B1(G234), .B2(new_n282), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT78), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n599), .A2(new_n600), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT25), .B1(new_n606), .B2(G902), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT25), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n599), .A2(new_n608), .A3(new_n282), .A4(new_n600), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n609), .A3(new_n601), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT79), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n605), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n605), .B2(new_n610), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n504), .B1(new_n576), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n560), .A2(new_n561), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n563), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n560), .A2(KEYINPUT32), .A3(new_n561), .ZN(new_n618));
  INV_X1    g432(.A(new_n575), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n612), .A2(new_n613), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(KEYINPUT80), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n503), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT99), .B(G101), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G3));
  AOI21_X1  g439(.A(G902), .B1(new_n551), .B2(new_n559), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n566), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n621), .A2(new_n431), .A3(new_n501), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT101), .Z(new_n635));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n292), .B1(new_n289), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n289), .A2(new_n636), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n287), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n346), .A2(new_n640), .A3(new_n347), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n339), .A2(new_n344), .A3(KEYINPUT33), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n349), .A2(G902), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n348), .A2(new_n349), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n418), .B2(new_n425), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n639), .A2(new_n300), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n635), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  INV_X1    g466(.A(new_n426), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(new_n351), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n300), .A3(new_n639), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n635), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR2_X1   g473(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n594), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n602), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n610), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n630), .A2(new_n631), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n502), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n501), .A2(new_n431), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n297), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n294), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n654), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n639), .A2(new_n663), .ZN(new_n675));
  OR4_X1    g489(.A1(new_n576), .A2(new_n668), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  INV_X1    g491(.A(new_n668), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n673), .B(KEYINPUT39), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT105), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n426), .A2(new_n351), .ZN(new_n684));
  INV_X1    g498(.A(new_n292), .ZN(new_n685));
  OR3_X1    g499(.A1(new_n684), .A2(new_n663), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n290), .A2(new_n291), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n562), .A2(new_n565), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n572), .A2(new_n510), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n282), .B1(new_n568), .B2(new_n510), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI211_X1 g508(.A(new_n686), .B(new_n689), .C1(new_n690), .C2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n682), .A2(new_n683), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT106), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n682), .A2(new_n698), .A3(new_n683), .A4(new_n695), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT107), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n321), .ZN(G45));
  NAND2_X1  g516(.A1(new_n647), .A2(new_n673), .ZN(new_n703));
  OR4_X1    g517(.A1(new_n576), .A2(new_n668), .A3(new_n675), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  AOI21_X1  g519(.A(new_n614), .B1(new_n690), .B2(new_n619), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n490), .A2(new_n282), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n492), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n709), .A2(new_n430), .A3(new_n648), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NOR3_X1   g527(.A1(new_n655), .A2(new_n709), .A3(new_n430), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n706), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  NOR2_X1   g530(.A1(new_n426), .A2(new_n351), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n663), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n690), .B2(new_n619), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n300), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n708), .A2(new_n431), .A3(new_n492), .A4(new_n639), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT108), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n582), .ZN(G21));
  NOR2_X1   g538(.A1(new_n709), .A2(new_n430), .ZN(new_n725));
  INV_X1    g539(.A(new_n639), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n299), .A3(new_n684), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n605), .A2(new_n610), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n561), .B(KEYINPUT109), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n569), .A2(new_n510), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n730), .B1(new_n731), .B2(new_n550), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n729), .B(new_n732), .C1(new_n626), .C2(new_n566), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n733), .A2(KEYINPUT110), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(KEYINPUT110), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n725), .B(new_n727), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n721), .B(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n663), .B(new_n732), .C1(new_n626), .C2(new_n566), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n703), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  INV_X1    g557(.A(new_n703), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n685), .B1(new_n290), .B2(new_n291), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n501), .A2(new_n431), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT42), .B1(new_n706), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n576), .A2(new_n746), .A3(new_n749), .A4(new_n728), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n352), .ZN(G33));
  INV_X1    g566(.A(new_n745), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n668), .A2(new_n674), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n706), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  OR2_X1    g570(.A1(new_n426), .A2(new_n646), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n632), .A2(new_n759), .A3(new_n663), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(new_n745), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(KEYINPUT112), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(KEYINPUT112), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n499), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n498), .B2(new_n499), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n768), .A2(new_n769), .A3(new_n491), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n493), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT46), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n772), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(KEYINPUT46), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n492), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n431), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n679), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n767), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n441), .ZN(G39));
  NOR4_X1   g594(.A1(new_n620), .A2(new_n621), .A3(new_n703), .A4(new_n753), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n776), .A2(KEYINPUT47), .A3(new_n431), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT47), .B1(new_n776), .B2(new_n431), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT113), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(KEYINPUT113), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NAND2_X1  g602(.A1(new_n759), .A2(new_n295), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT116), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n734), .A2(new_n735), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n685), .A3(new_n689), .A4(new_n725), .ZN(new_n793));
  NOR2_X1   g607(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n782), .A2(new_n783), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n708), .A2(KEYINPUT117), .A3(new_n492), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT117), .B1(new_n708), .B2(new_n492), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n797), .A2(new_n798), .A3(new_n431), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n745), .B(new_n792), .C1(new_n796), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n725), .A2(new_n745), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(new_n740), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n690), .A2(new_n694), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n801), .A2(new_n805), .A3(new_n614), .A4(new_n294), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n653), .A3(new_n646), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n795), .A2(new_n800), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n806), .A2(new_n647), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(G952), .A3(new_n254), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n576), .A2(new_n728), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n790), .A2(new_n813), .A3(new_n802), .ZN(new_n814));
  XOR2_X1   g628(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n812), .B(new_n816), .C1(new_n739), .C2(new_n792), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n808), .A2(new_n809), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n676), .A2(new_n742), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n639), .A2(new_n351), .A3(new_n426), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n663), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n805), .A2(new_n678), .A3(new_n673), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n821), .A2(new_n822), .A3(new_n704), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n676), .A2(new_n704), .A3(new_n742), .A4(new_n825), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n668), .A2(new_n614), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n626), .B(new_n628), .ZN(new_n833));
  INV_X1    g647(.A(new_n654), .ZN(new_n834));
  INV_X1    g648(.A(new_n647), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n301), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n665), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n831), .B1(new_n623), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n576), .A2(new_n504), .A3(new_n614), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT80), .B1(new_n620), .B2(new_n621), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n502), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n634), .A2(new_n836), .B1(new_n664), .B2(new_n502), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(KEYINPUT114), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n746), .A2(new_n740), .ZN(new_n846));
  INV_X1    g660(.A(new_n673), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n668), .A2(new_n753), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n719), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n849), .B(new_n755), .C1(new_n748), .C2(new_n750), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n706), .B1(new_n714), .B2(new_n710), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n851), .B(new_n736), .C1(new_n722), .C2(new_n720), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n845), .A2(new_n853), .A3(KEYINPUT115), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT115), .B1(new_n845), .B2(new_n853), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n830), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n676), .A2(new_n742), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n857), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n830), .B(new_n861), .C1(new_n854), .C2(new_n855), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n820), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n845), .A2(new_n853), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n860), .A2(KEYINPUT53), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n829), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI211_X1 g680(.A(KEYINPUT54), .B(new_n866), .C1(new_n856), .C2(new_n857), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n818), .A2(new_n819), .A3(new_n863), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(G952), .A2(G953), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n757), .A2(new_n728), .A3(new_n430), .A4(new_n685), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n689), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(KEYINPUT49), .B2(new_n709), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(KEYINPUT49), .B2(new_n709), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n868), .A2(new_n869), .B1(new_n805), .B2(new_n873), .ZN(G75));
  AOI21_X1  g688(.A(new_n866), .B1(new_n856), .B2(new_n857), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n282), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(G210), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n224), .B(new_n268), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT55), .Z(new_n880));
  AND3_X1   g694(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n877), .B2(new_n878), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n254), .A2(G952), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT120), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(G51));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n864), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n845), .A2(new_n853), .A3(KEYINPUT115), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n829), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(KEYINPUT53), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT54), .B1(new_n891), .B2(new_n866), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n875), .A2(new_n820), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n493), .B(KEYINPUT57), .Z(new_n896));
  OAI21_X1  g710(.A(new_n490), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n876), .A2(new_n770), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n885), .B1(new_n897), .B2(new_n898), .ZN(G54));
  NAND3_X1  g713(.A1(new_n876), .A2(KEYINPUT58), .A3(G475), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(new_n410), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n410), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n885), .B1(new_n901), .B2(new_n902), .ZN(G60));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n904));
  XNOR2_X1  g718(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n349), .A2(new_n282), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n905), .B(new_n906), .Z(new_n907));
  OAI21_X1  g721(.A(new_n862), .B1(new_n890), .B2(KEYINPUT53), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n909), .B2(new_n893), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n641), .A2(new_n642), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n904), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n907), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n867), .B2(new_n863), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(KEYINPUT122), .A3(new_n911), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n911), .A2(new_n907), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n885), .B1(new_n894), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n913), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n913), .A2(new_n916), .A3(new_n918), .A4(KEYINPUT123), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT124), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT60), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n875), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n661), .ZN(new_n928));
  INV_X1    g742(.A(new_n606), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n928), .B(new_n884), .C1(new_n929), .C2(new_n927), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT61), .Z(G66));
  INV_X1    g745(.A(G224), .ZN(new_n932));
  OAI21_X1  g746(.A(G953), .B1(new_n298), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT125), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n852), .B1(new_n839), .B2(new_n844), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(G953), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n224), .B1(G898), .B2(new_n254), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G69));
  OAI21_X1  g752(.A(new_n544), .B1(new_n540), .B2(KEYINPUT30), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n405), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n669), .B2(new_n254), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n779), .B1(new_n785), .B2(new_n786), .ZN(new_n942));
  NOR4_X1   g756(.A1(new_n778), .A2(new_n576), .A3(new_n728), .A4(new_n823), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n821), .A2(new_n704), .ZN(new_n944));
  INV_X1    g758(.A(new_n751), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n945), .A3(new_n755), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n941), .B1(new_n948), .B2(new_n254), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n697), .A2(new_n699), .A3(new_n944), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n697), .A2(KEYINPUT62), .A3(new_n699), .A4(new_n944), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n681), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n753), .B1(new_n834), .B2(new_n835), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n955), .B(new_n956), .C1(new_n841), .C2(new_n840), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n942), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n940), .B1(new_n958), .B2(new_n254), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n949), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n471), .B2(new_n669), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G72));
  NAND3_X1  g776(.A1(new_n942), .A2(new_n935), .A3(new_n947), .ZN(new_n963));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n963), .A2(KEYINPUT127), .A3(new_n965), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n572), .A2(new_n510), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n965), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n692), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n885), .B1(new_n908), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n954), .A2(new_n942), .A3(new_n935), .A4(new_n957), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n965), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n977), .B2(new_n692), .ZN(new_n978));
  AOI211_X1 g792(.A(KEYINPUT126), .B(new_n691), .C1(new_n976), .C2(new_n965), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n971), .B(new_n974), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(G57));
endmodule


