//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT77), .B(KEYINPUT22), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n190), .B(new_n191), .Z(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT78), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  XNOR2_X1  g009(.A(G125), .B(G140), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(KEYINPUT16), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT74), .B1(new_n197), .B2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT74), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n202));
  OR2_X1    g016(.A1(G125), .A2(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(G125), .A2(G140), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n200), .B(new_n201), .C1(new_n205), .C2(new_n195), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n198), .A2(new_n199), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G128), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(KEYINPUT70), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT70), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n212), .B1(new_n216), .B2(G119), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n210), .B1(new_n217), .B2(new_n208), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G110), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(G119), .ZN(new_n220));
  INV_X1    g034(.A(new_n212), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT24), .B(G110), .ZN(new_n223));
  OR2_X1    g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n207), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT76), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT75), .B(G110), .Z(new_n227));
  OAI211_X1 g041(.A(new_n210), .B(new_n227), .C1(new_n217), .C2(new_n208), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n223), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n196), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(G146), .B2(new_n197), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n225), .A2(new_n226), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n226), .B1(new_n225), .B2(new_n234), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n193), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n225), .A2(new_n234), .A3(new_n192), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n239), .A2(new_n240), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n237), .A2(new_n238), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT80), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT25), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT25), .B1(new_n243), .B2(new_n244), .ZN(new_n246));
  INV_X1    g060(.A(G217), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(G234), .B2(new_n238), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n245), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n248), .A2(G902), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n237), .A2(new_n241), .A3(new_n242), .A4(new_n251), .ZN(new_n252));
  XOR2_X1   g066(.A(new_n252), .B(KEYINPUT81), .Z(new_n253));
  OAI21_X1  g067(.A(new_n187), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n243), .A2(new_n244), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT25), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n248), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n252), .B(KEYINPUT81), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(KEYINPUT82), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT0), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(new_n211), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(G146), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(G146), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n201), .A2(KEYINPUT65), .A3(G143), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n201), .A2(G143), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n264), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G131), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(G137), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(G137), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT11), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n283), .B2(G137), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n284), .A2(KEYINPUT11), .A3(new_n288), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n281), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT11), .ZN(new_n293));
  INV_X1    g107(.A(G137), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT67), .B1(new_n294), .B2(G134), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(G134), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT66), .B1(new_n294), .B2(G134), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n281), .B(new_n291), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n280), .B1(new_n292), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(G143), .B2(new_n201), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n275), .B1(new_n305), .B2(new_n216), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n278), .A2(new_n304), .A3(G128), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n283), .A2(G137), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n285), .B2(KEYINPUT69), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n296), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G131), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n308), .A2(new_n300), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n276), .A2(new_n279), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n295), .A2(new_n296), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n316), .A2(KEYINPUT11), .B1(new_n284), .B2(new_n288), .ZN(new_n317));
  INV_X1    g131(.A(new_n291), .ZN(new_n318));
  OAI21_X1  g132(.A(G131), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n315), .B1(new_n319), .B2(new_n300), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n303), .A2(new_n314), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n324));
  INV_X1    g138(.A(G116), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(G119), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n209), .A2(KEYINPUT71), .A3(G116), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT2), .B(G113), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n332));
  INV_X1    g146(.A(new_n330), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT72), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n335));
  NOR3_X1   g149(.A1(new_n329), .A2(new_n335), .A3(new_n330), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n331), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n323), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(G237), .A2(G953), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G210), .ZN(new_n340));
  INV_X1    g154(.A(G101), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n343));
  XOR2_X1   g157(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g158(.A(new_n337), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n302), .A2(new_n345), .A3(new_n314), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT28), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n302), .A2(KEYINPUT28), .A3(new_n345), .A4(new_n314), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n338), .A2(new_n344), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n346), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n308), .A2(new_n300), .A3(new_n313), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT30), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n320), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n323), .B2(new_n353), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n351), .B1(new_n355), .B2(new_n337), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n263), .B(new_n350), .C1(new_n356), .C2(new_n344), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT73), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n337), .B1(new_n320), .B2(new_n352), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n348), .A2(new_n349), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n344), .ZN(new_n361));
  OR3_X1    g175(.A1(new_n360), .A2(new_n263), .A3(new_n361), .ZN(new_n362));
  AOI211_X1 g176(.A(new_n345), .B(new_n354), .C1(new_n323), .C2(new_n353), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n361), .B1(new_n363), .B2(new_n351), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n263), .A4(new_n350), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n358), .A2(new_n238), .A3(new_n362), .A4(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n367), .A2(G472), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n369));
  NOR2_X1   g183(.A1(G472), .A2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n354), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n320), .A2(new_n321), .ZN(new_n372));
  AOI211_X1 g186(.A(KEYINPUT68), .B(new_n315), .C1(new_n319), .C2(new_n300), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n372), .A2(new_n373), .A3(new_n352), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n337), .B(new_n371), .C1(new_n374), .C2(KEYINPUT30), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT31), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n346), .A4(new_n344), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n338), .A2(new_n348), .A3(new_n349), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n361), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n376), .B1(new_n356), .B2(new_n344), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n369), .B(new_n370), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n375), .A2(new_n346), .A3(new_n344), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT31), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n377), .A3(new_n379), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n369), .B1(new_n386), .B2(new_n370), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n262), .B1(new_n368), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n319), .A2(new_n300), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n273), .A2(new_n277), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n305), .B2(new_n211), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n307), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G104), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT3), .B1(new_n395), .B2(G107), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(G107), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n396), .A2(new_n399), .A3(new_n341), .A4(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n398), .A2(G104), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n395), .A2(G107), .ZN(new_n403));
  OAI21_X1  g217(.A(G101), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n394), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT10), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n308), .A2(KEYINPUT10), .A3(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n396), .A2(new_n399), .A3(KEYINPUT84), .A4(new_n400), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(G101), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n413), .A2(new_n417), .A3(G101), .A4(new_n414), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n280), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT85), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT85), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n416), .A2(new_n421), .A3(new_n280), .A4(new_n418), .ZN(new_n422));
  AOI211_X1 g236(.A(new_n391), .B(new_n410), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  INV_X1    g238(.A(G227), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G953), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n424), .B(new_n426), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n390), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n420), .A2(new_n422), .ZN(new_n430));
  INV_X1    g244(.A(new_n410), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n391), .ZN(new_n433));
  INV_X1    g247(.A(new_n391), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(new_n434), .A3(new_n431), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT86), .A3(new_n427), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n406), .B1(new_n308), .B2(new_n405), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n391), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n428), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n238), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(G469), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n434), .B1(new_n430), .B2(new_n431), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n428), .B1(new_n448), .B2(new_n423), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n435), .A2(new_n441), .A3(new_n427), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G469), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n238), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n437), .B2(new_n443), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT87), .B1(new_n454), .B2(new_n452), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n447), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G237), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n188), .A3(G214), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n271), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n339), .A2(G143), .A3(G214), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G131), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n281), .A3(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n281), .B1(new_n459), .B2(new_n460), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT17), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n468), .A2(new_n207), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n470));
  XNOR2_X1  g284(.A(G113), .B(G122), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n395), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n466), .A2(KEYINPUT18), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT18), .A2(G131), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n459), .A2(new_n460), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n196), .A2(KEYINPUT90), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n203), .A2(new_n477), .A3(new_n204), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n201), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n473), .B(new_n475), .C1(new_n232), .C2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n469), .A2(new_n470), .A3(new_n472), .A4(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n472), .B(new_n480), .C1(new_n468), .C2(new_n207), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT93), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n462), .A2(new_n464), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n199), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT19), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n476), .B2(new_n478), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n231), .A2(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n488), .A2(G146), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n480), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT92), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n472), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n480), .B(KEYINPUT92), .C1(new_n486), .C2(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n484), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT20), .ZN(new_n498));
  NOR2_X1   g312(.A1(G475), .A2(G902), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT94), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n481), .A2(new_n483), .B1(new_n494), .B2(new_n495), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT20), .B1(new_n503), .B2(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G116), .B(G122), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n506), .A2(KEYINPUT95), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(KEYINPUT95), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G107), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n508), .A3(new_n398), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n216), .A2(G143), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT13), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(G134), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n271), .A2(G128), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n513), .A2(new_n283), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n283), .B1(new_n513), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n513), .A2(new_n514), .A3(G134), .A4(new_n516), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n512), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n325), .A2(KEYINPUT14), .A3(G122), .ZN(new_n522));
  INV_X1    g336(.A(new_n506), .ZN(new_n523));
  OAI211_X1 g337(.A(G107), .B(new_n522), .C1(new_n523), .C2(KEYINPUT14), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n511), .B(new_n524), .C1(new_n517), .C2(new_n518), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT9), .B(G234), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT83), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n527), .A2(new_n247), .A3(G953), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n521), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n521), .B2(new_n525), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n238), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G478), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(KEYINPUT15), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n531), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n469), .A2(new_n480), .ZN(new_n536));
  INV_X1    g350(.A(new_n472), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n484), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n238), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G475), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n188), .A2(G952), .ZN(new_n542));
  INV_X1    g356(.A(G234), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n457), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(G902), .B(G953), .C1(new_n543), .C2(new_n457), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n546), .B(KEYINPUT96), .Z(new_n547));
  XOR2_X1   g361(.A(KEYINPUT21), .B(G898), .Z(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n505), .A2(new_n535), .A3(new_n541), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT97), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n531), .B(new_n533), .ZN(new_n554));
  INV_X1    g368(.A(G475), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n539), .B2(new_n238), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT97), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n551), .A4(new_n505), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G214), .B1(G237), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  MUX2_X1   g376(.A(new_n308), .B(new_n280), .S(G125), .Z(new_n563));
  INV_X1    g377(.A(G224), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G953), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT7), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT89), .B1(new_n280), .B2(new_n194), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n568), .A2(KEYINPUT89), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n569), .A2(new_n570), .B1(new_n563), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n416), .A2(new_n337), .A3(new_n418), .ZN(new_n573));
  XOR2_X1   g387(.A(G110), .B(G122), .Z(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n332), .A2(KEYINPUT72), .A3(new_n333), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n335), .B1(new_n329), .B2(new_n330), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT5), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n209), .A3(G116), .ZN(new_n580));
  OAI211_X1 g394(.A(G113), .B(new_n580), .C1(new_n329), .C2(new_n579), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n405), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n573), .A2(new_n575), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n574), .B(KEYINPUT8), .Z(new_n584));
  INV_X1    g398(.A(new_n582), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n405), .B1(new_n578), .B2(new_n581), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n572), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n573), .A2(new_n582), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT88), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n589), .A2(new_n574), .B1(new_n590), .B2(KEYINPUT6), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(KEYINPUT6), .ZN(new_n592));
  AOI211_X1 g406(.A(new_n575), .B(new_n592), .C1(new_n573), .C2(new_n582), .ZN(new_n593));
  INV_X1    g407(.A(new_n583), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n563), .B(new_n565), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n238), .B(new_n588), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G210), .B1(G237), .B2(G902), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n589), .A2(new_n574), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n592), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT6), .A4(new_n574), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n583), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n596), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n598), .A3(new_n588), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n562), .B1(new_n600), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(G221), .B1(new_n527), .B2(G902), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n456), .A2(new_n560), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n389), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT98), .B(G101), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G3));
  OAI21_X1  g427(.A(new_n238), .B1(new_n380), .B2(new_n381), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n614), .A2(G472), .B1(new_n370), .B2(new_n386), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n262), .A2(new_n456), .A3(new_n609), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n608), .A2(new_n551), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n556), .B1(new_n504), .B2(new_n502), .ZN(new_n618));
  OR3_X1    g432(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT33), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT33), .B1(new_n529), .B2(new_n530), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(G478), .A3(new_n620), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n531), .A2(G478), .ZN(new_n622));
  NAND2_X1  g436(.A1(G478), .A2(G902), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT99), .B1(new_n617), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n608), .A2(new_n625), .A3(new_n628), .A4(new_n551), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n616), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(new_n395), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND2_X1  g448(.A1(new_n618), .A2(new_n554), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n616), .A2(new_n617), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT101), .B(KEYINPUT102), .Z(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT35), .B(G107), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n636), .B(new_n639), .ZN(G9));
  OR3_X1    g454(.A1(new_n193), .A2(KEYINPUT103), .A3(KEYINPUT36), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT103), .B1(new_n193), .B2(KEYINPUT36), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n235), .A2(new_n236), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n643), .B(new_n644), .Z(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n251), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n259), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n615), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n610), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT37), .B(G110), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  NAND2_X1  g465(.A1(new_n367), .A2(G472), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n370), .B1(new_n380), .B2(new_n381), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT32), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n382), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n545), .B1(new_n547), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n635), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n656), .A2(new_n647), .A3(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n456), .A2(new_n608), .A3(new_n609), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  NOR2_X1   g477(.A1(new_n356), .A2(new_n361), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n351), .A2(new_n344), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n359), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n238), .ZN(new_n667));
  OAI21_X1  g481(.A(G472), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n655), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n647), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n600), .A2(new_n607), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT38), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n674), .A2(new_n535), .A3(new_n562), .A4(new_n618), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n456), .A2(new_n609), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n658), .B(KEYINPUT39), .Z(new_n677));
  AND2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n678), .A2(KEYINPUT104), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(KEYINPUT104), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n679), .A2(KEYINPUT40), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT40), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n671), .B(new_n675), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  AOI22_X1  g498(.A1(G472), .A2(new_n367), .B1(new_n654), .B2(new_n382), .ZN(new_n685));
  INV_X1    g499(.A(new_n647), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n626), .A2(new_n658), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n608), .A3(new_n676), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n427), .B1(new_n433), .B2(new_n435), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n435), .A2(new_n441), .A3(new_n427), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n238), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n609), .A3(new_n453), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n695), .A2(KEYINPUT105), .A3(new_n609), .A4(new_n453), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n656), .A3(new_n262), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n691), .B1(new_n701), .B2(new_n630), .ZN(new_n702));
  INV_X1    g516(.A(new_n630), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n259), .A2(KEYINPUT82), .A3(new_n260), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT82), .B1(new_n259), .B2(new_n260), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n685), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n703), .A2(new_n707), .A3(KEYINPUT106), .A4(new_n700), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND2_X1  g525(.A1(new_n698), .A2(new_n699), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n685), .A2(new_n712), .A3(new_n706), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n617), .A2(new_n635), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  NAND3_X1  g530(.A1(new_n698), .A2(new_n608), .A3(new_n699), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n698), .A2(new_n719), .A3(new_n608), .A4(new_n699), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n656), .A2(new_n560), .A3(new_n647), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n344), .B1(new_n360), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n726), .B2(new_n360), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n385), .A2(new_n728), .A3(new_n377), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n614), .A2(G472), .B1(new_n729), .B2(new_n370), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n250), .A2(new_n253), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n731), .B1(new_n730), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n618), .B2(new_n535), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n505), .A2(new_n541), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(KEYINPUT110), .A3(new_n554), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n617), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n698), .A4(new_n699), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n725), .B1(new_n735), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n730), .A2(new_n732), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AND4_X1   g561(.A1(new_n741), .A2(new_n740), .A3(new_n698), .A4(new_n699), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT111), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NAND3_X1  g565(.A1(new_n688), .A2(new_n647), .A3(new_n730), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n721), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  INV_X1    g569(.A(new_n732), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n685), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n453), .B1(new_n454), .B2(new_n452), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n758), .A2(new_n609), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n600), .A2(new_n607), .A3(new_n561), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n626), .A3(new_n658), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n758), .A2(new_n760), .A3(new_n609), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n656), .A2(new_n262), .A3(new_n688), .A4(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n763), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NAND3_X1  g585(.A1(new_n707), .A2(new_n659), .A3(new_n764), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n738), .A2(new_n624), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT43), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(KEYINPUT115), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(KEYINPUT115), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n686), .A2(new_n615), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n774), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n444), .B(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(G469), .ZN(new_n783));
  NAND2_X1  g597(.A1(G469), .A2(G902), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT113), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT114), .ZN(new_n790));
  INV_X1    g604(.A(new_n453), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n785), .B2(KEYINPUT113), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n793), .A3(new_n788), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n786), .A2(new_n790), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n609), .A2(new_n781), .A3(new_n795), .A4(new_n677), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n779), .A2(new_n780), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n761), .B1(new_n797), .B2(KEYINPUT44), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  AND3_X1   g614(.A1(new_n795), .A2(KEYINPUT47), .A3(new_n609), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT47), .B1(new_n795), .B2(new_n609), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n685), .A3(new_n706), .A4(new_n762), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  NAND2_X1  g621(.A1(new_n776), .A2(new_n545), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n808), .A2(new_n712), .A3(new_n761), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n757), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT48), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n735), .A2(new_n808), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n721), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n542), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n712), .A2(new_n761), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n262), .A3(new_n545), .A4(new_n670), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n618), .A2(new_n624), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n673), .A2(new_n561), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n812), .A2(new_n700), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n812), .A2(KEYINPUT50), .A3(new_n700), .A4(new_n820), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n819), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n695), .A2(new_n453), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n609), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n802), .A2(new_n804), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n812), .A2(new_n760), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT119), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n826), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n809), .A2(new_n647), .A3(new_n730), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(KEYINPUT120), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n801), .A2(new_n803), .A3(new_n828), .ZN(new_n837));
  INV_X1    g651(.A(new_n832), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n835), .B(new_n825), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n834), .A2(KEYINPUT120), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n834), .A2(KEYINPUT120), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n814), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n658), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n760), .A2(new_n505), .A3(new_n557), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n687), .A2(new_n676), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n764), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT116), .B1(new_n752), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n772), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n770), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n721), .A2(new_n722), .B1(new_n713), .B2(new_n714), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n625), .B1(new_n554), .B2(new_n618), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n616), .A2(new_n617), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n610), .B1(new_n389), .B2(new_n648), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n709), .A2(new_n750), .A3(new_n851), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n753), .A2(new_n764), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(KEYINPUT116), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n850), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n737), .A2(new_n608), .A3(new_n739), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(new_n759), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n686), .A3(new_n844), .A4(new_n669), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n754), .A2(new_n662), .A3(new_n689), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n866), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n721), .A2(new_n753), .B1(new_n660), .B2(new_n661), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT52), .A3(new_n689), .A4(new_n863), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n867), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n709), .A2(new_n750), .A3(new_n851), .A4(new_n855), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n846), .A2(new_n772), .A3(new_n848), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n765), .A2(new_n767), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT112), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n875), .B1(new_n879), .B2(new_n763), .ZN(new_n880));
  INV_X1    g694(.A(new_n858), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n868), .A2(new_n870), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n873), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n872), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n882), .A2(new_n884), .A3(new_n873), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n859), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n882), .A2(KEYINPUT117), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n891), .A3(new_n867), .A4(new_n871), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n888), .B1(new_n892), .B2(new_n873), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n843), .B(new_n887), .C1(new_n886), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n816), .A2(new_n626), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n894), .A2(new_n895), .B1(G952), .B2(G953), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n827), .B(KEYINPUT49), .Z(new_n897));
  NOR2_X1   g711(.A1(new_n673), .A2(new_n756), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n775), .A2(new_n561), .A3(new_n609), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n670), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n896), .A2(new_n900), .ZN(G75));
  AOI21_X1  g715(.A(new_n238), .B1(new_n872), .B2(new_n885), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(G210), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n604), .B(new_n605), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n905), .A2(KEYINPUT121), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n188), .A2(G952), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n905), .B2(KEYINPUT121), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n905), .B2(KEYINPUT121), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(G51));
  XOR2_X1   g727(.A(new_n784), .B(KEYINPUT57), .Z(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT53), .B1(new_n859), .B2(new_n883), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n871), .A2(new_n867), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n874), .A2(new_n880), .A3(KEYINPUT53), .A4(new_n881), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT54), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n915), .B1(new_n920), .B2(new_n887), .ZN(new_n921));
  INV_X1    g735(.A(new_n451), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT122), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n872), .A2(new_n886), .A3(new_n885), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n886), .B1(new_n872), .B2(new_n885), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n914), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n927), .A3(new_n451), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n902), .A2(G469), .A3(new_n782), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n923), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n910), .ZN(G54));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT58), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n933), .A2(new_n555), .A3(KEYINPUT123), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n238), .B(new_n934), .C1(new_n872), .C2(new_n885), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT123), .B1(new_n933), .B2(new_n555), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n932), .B1(new_n937), .B2(new_n503), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n935), .A2(KEYINPUT124), .A3(new_n497), .A4(new_n936), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n503), .ZN(new_n940));
  AND4_X1   g754(.A1(new_n910), .A2(new_n938), .A3(new_n939), .A4(new_n940), .ZN(G60));
  NAND2_X1  g755(.A1(new_n619), .A2(new_n620), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n887), .B1(new_n893), .B2(new_n886), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n623), .B(KEYINPUT59), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n944), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n920), .B2(new_n887), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n945), .A2(new_n909), .A3(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(new_n872), .A2(new_n885), .ZN(new_n949));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT60), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n237), .A2(new_n241), .A3(new_n242), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n645), .A3(new_n951), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n910), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT61), .B1(new_n955), .B2(KEYINPUT125), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G66));
  AOI21_X1  g772(.A(new_n188), .B1(new_n548), .B2(G224), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n856), .B2(new_n188), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n595), .B1(G898), .B2(new_n188), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(G69));
  NOR2_X1   g776(.A1(new_n488), .A2(new_n490), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n355), .B(new_n963), .Z(new_n964));
  AND2_X1   g778(.A1(new_n869), .A2(new_n689), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n795), .A2(new_n609), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n966), .A2(new_n677), .A3(new_n757), .A4(new_n861), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n799), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(new_n806), .A3(new_n770), .A4(new_n772), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n964), .B1(new_n969), .B2(new_n188), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n425), .A2(G900), .A3(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n683), .A2(KEYINPUT126), .A3(new_n973), .A4(new_n965), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n973), .A2(KEYINPUT126), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n679), .A2(new_n680), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n976), .A2(new_n389), .A3(new_n852), .ZN(new_n977));
  AOI22_X1  g791(.A1(new_n977), .A2(new_n760), .B1(new_n796), .B2(new_n798), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n974), .A2(new_n806), .A3(new_n975), .A4(new_n978), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n683), .A2(new_n965), .B1(KEYINPUT126), .B2(new_n973), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n964), .B1(new_n981), .B2(G953), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n425), .A2(new_n657), .A3(new_n188), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n972), .B1(new_n982), .B2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n364), .A2(new_n384), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n893), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n986), .B1(new_n969), .B2(new_n856), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n375), .A2(new_n665), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n909), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n979), .A2(new_n856), .A3(new_n980), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n664), .B1(new_n994), .B2(new_n987), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(KEYINPUT127), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n997), .B(new_n664), .C1(new_n994), .C2(new_n987), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n993), .B1(new_n996), .B2(new_n998), .ZN(G57));
endmodule


