//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n527, new_n528,
    new_n529, new_n530, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n543, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(new_n465), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n468), .B1(new_n473), .B2(G2105), .ZN(G160));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n461), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n478), .A2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(G136), .B2(new_n484), .ZN(G162));
  NOR2_X1   g060(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n466), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n475), .B2(new_n476), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n461), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n488), .ZN(new_n496));
  INV_X1    g071(.A(new_n486), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n477), .A2(new_n496), .A3(new_n461), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  OAI21_X1  g075(.A(KEYINPUT5), .B1(KEYINPUT71), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(KEYINPUT72), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n504), .A2(KEYINPUT71), .A3(KEYINPUT5), .A4(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(G88), .B1(G50), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n506), .A2(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  XOR2_X1   g088(.A(new_n513), .B(KEYINPUT73), .Z(new_n514));
  OAI21_X1  g089(.A(G651), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n510), .A2(G51), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n508), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  AOI22_X1  g101(.A1(new_n508), .A2(G90), .B1(G52), .B2(new_n510), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT74), .ZN(G171));
  NAND2_X1  g106(.A1(new_n506), .A2(new_n507), .ZN(new_n532));
  INV_X1    g107(.A(G81), .ZN(new_n533));
  INV_X1    g108(.A(G43), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n509), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT75), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n528), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT76), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  NAND2_X1  g121(.A1(G78), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(new_n506), .ZN(new_n548));
  INV_X1    g123(.A(G65), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G651), .B1(new_n508), .B2(G91), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OR3_X1    g127(.A1(new_n509), .A2(KEYINPUT9), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT9), .B1(new_n509), .B2(new_n552), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n551), .B1(new_n557), .B2(new_n558), .ZN(G299));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n530), .B(new_n560), .ZN(G301));
  OAI21_X1  g136(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n508), .A2(G87), .B1(G49), .B2(new_n510), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(G288));
  NAND3_X1  g141(.A1(new_n507), .A2(G48), .A3(G543), .ZN(new_n567));
  INV_X1    g142(.A(G86), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n532), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  AND2_X1   g145(.A1(G73), .A2(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n506), .B2(G61), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n528), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n528), .ZN(new_n576));
  XNOR2_X1  g151(.A(KEYINPUT79), .B(G85), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n508), .A2(new_n577), .B1(new_n510), .B2(G47), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(new_n508), .A2(G92), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT10), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n548), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(G868), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g164(.A(new_n588), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g165(.A1(G286), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(G299), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G280));
  XOR2_X1   g168(.A(G280), .B(KEYINPUT80), .Z(G297));
  NOR2_X1   g169(.A1(new_n587), .A2(G559), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n582), .A2(new_n586), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n595), .B1(G860), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT81), .ZN(G148));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n539), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n595), .B2(new_n599), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n477), .A2(new_n462), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT83), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT13), .Z(new_n607));
  INV_X1    g182(.A(G2100), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n484), .A2(G135), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n479), .A2(G123), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n461), .A2(G111), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2096), .Z(new_n616));
  NAND3_X1  g191(.A1(new_n609), .A2(new_n610), .A3(new_n616), .ZN(G156));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2427), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(new_n620), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n623), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  AND3_X1   g206(.A1(new_n630), .A2(G14), .A3(new_n631), .ZN(G401));
  XNOR2_X1  g207(.A(G2067), .B(G2678), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT84), .ZN(new_n634));
  NOR2_X1   g209(.A1(G2072), .A2(G2078), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n442), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2084), .B(G2090), .ZN(new_n637));
  NOR3_X1   g212(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT18), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n636), .A2(KEYINPUT85), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(KEYINPUT85), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(new_n636), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n642), .B(new_n637), .C1(new_n644), .C2(new_n634), .ZN(new_n645));
  INV_X1    g220(.A(new_n637), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n634), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n639), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2096), .B(G2100), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n651));
  XNOR2_X1  g226(.A(G1971), .B(G1976), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT20), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n654), .B(new_n655), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n658), .B(new_n659), .C1(new_n653), .C2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1991), .B(G1996), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n665), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(G229));
  NOR2_X1   g246(.A1(G6), .A2(G16), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n572), .A2(new_n528), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n673), .A2(new_n569), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n672), .B1(new_n674), .B2(G16), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT32), .ZN(new_n676));
  INV_X1    g251(.A(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n679), .A2(G23), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G288), .B2(G16), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(G22), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n679), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G1971), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n678), .A2(new_n683), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n690));
  OR2_X1    g265(.A1(G25), .A2(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n479), .A2(G119), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n461), .A2(G107), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n484), .A2(KEYINPUT88), .A3(G131), .ZN(new_n695));
  AOI21_X1  g270(.A(KEYINPUT88), .B1(new_n484), .B2(G131), .ZN(new_n696));
  OAI221_X1 g271(.A(new_n692), .B1(new_n693), .B2(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n691), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT35), .B(G1991), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1986), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n689), .A2(new_n690), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(KEYINPUT36), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n689), .A2(new_n708), .A3(new_n690), .A4(new_n705), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n484), .A2(G139), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT95), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n711), .B(new_n714), .C1(new_n461), .C2(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(G33), .B(new_n716), .S(G29), .Z(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(G2072), .ZN(new_n718));
  INV_X1    g293(.A(G28), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT30), .ZN(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n719), .B2(KEYINPUT30), .ZN(new_n721));
  OR2_X1    g296(.A1(KEYINPUT31), .A2(G11), .ZN(new_n722));
  NAND2_X1  g297(.A1(KEYINPUT31), .A2(G11), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n615), .B2(new_n698), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n698), .B1(new_n726), .B2(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G160), .B2(G29), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G2084), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n718), .A2(new_n725), .A3(new_n730), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n679), .A2(G21), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G286), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT96), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n734), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n698), .A2(G27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n698), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n737), .B1(G2078), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G2078), .B2(new_n739), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n731), .A2(new_n736), .A3(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n698), .A2(G32), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n484), .A2(G141), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n479), .A2(G129), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT26), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n748), .A2(new_n749), .B1(G105), .B2(new_n462), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n744), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n743), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n717), .A2(G2072), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n679), .A2(G5), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G171), .B2(new_n679), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n754), .B1(new_n752), .B2(new_n753), .C1(G1961), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n742), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(G1961), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT97), .Z(new_n760));
  AND3_X1   g335(.A1(new_n758), .A2(KEYINPUT98), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(KEYINPUT98), .B1(new_n758), .B2(new_n760), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n698), .A2(G26), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n484), .A2(G140), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n479), .A2(G128), .ZN(new_n768));
  OAI21_X1  g343(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g345(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n771));
  OAI221_X1 g346(.A(G2104), .B1(G116), .B2(new_n461), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT91), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n767), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n766), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2067), .ZN(new_n780));
  NOR2_X1   g355(.A1(G4), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n596), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT89), .B(G1348), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n679), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n540), .B2(new_n679), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G1341), .Z(new_n787));
  NAND3_X1  g362(.A1(new_n780), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n698), .A2(G35), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT99), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n698), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT29), .B(G2090), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n679), .A2(G20), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT23), .Z(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G299), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT100), .B(G1956), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  AOI211_X1 g375(.A(new_n795), .B(new_n800), .C1(new_n788), .C2(new_n789), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n710), .A2(new_n763), .A3(new_n790), .A4(new_n801), .ZN(G150));
  INV_X1    g377(.A(G150), .ZN(G311));
  NAND2_X1  g378(.A1(new_n596), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT38), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n508), .A2(G93), .B1(G55), .B2(new_n510), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n528), .B2(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n539), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n539), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n805), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n813));
  AOI21_X1  g388(.A(G860), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n808), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT37), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(G145));
  INV_X1    g393(.A(G37), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT101), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n491), .B2(new_n494), .ZN(new_n821));
  OR2_X1    g396(.A1(G102), .A2(G2105), .ZN(new_n822));
  INV_X1    g397(.A(G114), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G2105), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n824), .A3(G2104), .ZN(new_n825));
  AND2_X1   g400(.A1(G126), .A2(G2105), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n464), .B2(new_n465), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n825), .A2(new_n827), .A3(KEYINPUT101), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n821), .A2(new_n489), .A3(new_n498), .A4(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n778), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n832));
  INV_X1    g407(.A(new_n751), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n716), .A2(KEYINPUT102), .A3(new_n751), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n778), .A2(new_n835), .A3(new_n834), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n830), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n484), .A2(G142), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n479), .A2(G130), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(G118), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n843), .A2(KEYINPUT103), .B1(new_n844), .B2(G2105), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(KEYINPUT103), .B2(new_n843), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n606), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(new_n697), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n837), .A2(new_n830), .A3(new_n838), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n840), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n851), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n849), .B1(new_n853), .B2(new_n839), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n615), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G162), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NOR4_X1   g432(.A1(new_n853), .A2(new_n839), .A3(KEYINPUT104), .A4(new_n850), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n850), .A2(KEYINPUT104), .B1(new_n853), .B2(new_n839), .ZN(new_n859));
  INV_X1    g434(.A(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n819), .B(new_n857), .C1(new_n858), .C2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(G395));
  XNOR2_X1  g439(.A(G288), .B(G290), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(KEYINPUT107), .ZN(new_n866));
  XNOR2_X1  g441(.A(G303), .B(KEYINPUT106), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n674), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(KEYINPUT107), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n867), .B(G305), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(KEYINPUT107), .A3(new_n865), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n595), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n811), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n596), .A2(new_n592), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n587), .A2(G299), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n809), .A2(new_n810), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(new_n876), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n811), .A2(new_n595), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n878), .A2(new_n886), .A3(new_n879), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n886), .B1(new_n878), .B2(new_n879), .ZN(new_n889));
  OAI22_X1  g464(.A1(new_n884), .A2(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT108), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n599), .B1(new_n875), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n882), .A2(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n873), .B(KEYINPUT42), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n882), .A2(new_n890), .A3(KEYINPUT108), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT109), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n808), .A2(new_n599), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n892), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(G295));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(G331));
  NAND2_X1  g480(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT111), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n887), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n888), .A2(KEYINPUT111), .ZN(new_n909));
  NAND2_X1  g484(.A1(G301), .A2(G286), .ZN(new_n910));
  NAND2_X1  g485(.A1(G171), .A2(G168), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(new_n811), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n910), .A2(new_n911), .B1(new_n809), .B2(new_n810), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n908), .B(new_n909), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n883), .A2(new_n910), .A3(new_n911), .ZN(new_n916));
  INV_X1    g491(.A(new_n914), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n881), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n873), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n870), .A2(new_n872), .ZN(new_n921));
  OAI22_X1  g496(.A1(new_n913), .A2(new_n914), .B1(new_n888), .B2(new_n889), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n924));
  NAND4_X1  g499(.A1(new_n920), .A2(new_n819), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n819), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n921), .B1(new_n922), .B2(new_n918), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n925), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n921), .B1(new_n915), .B2(new_n918), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n918), .A2(new_n922), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n873), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n935), .A2(new_n819), .A3(new_n923), .A4(new_n924), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n930), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n931), .A2(new_n937), .ZN(G397));
  INV_X1    g513(.A(G2067), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n831), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n778), .A2(G2067), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n833), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G1384), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n829), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(G160), .A2(G40), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n948), .ZN(new_n950));
  NAND2_X1  g525(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n950), .A2(G1996), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n948), .B(new_n953), .C1(KEYINPUT124), .C2(KEYINPUT46), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n954), .B2(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT125), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n949), .A2(new_n958), .A3(new_n955), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(KEYINPUT47), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n751), .B(new_n953), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n940), .A2(new_n941), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n700), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n697), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n940), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n948), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n697), .B(new_n963), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n950), .ZN(new_n969));
  NOR2_X1   g544(.A1(G290), .A2(G1986), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT112), .Z(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n948), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n972), .B(KEYINPUT48), .Z(new_n973));
  OAI211_X1 g548(.A(new_n960), .B(new_n966), .C1(new_n969), .C2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT47), .B1(new_n957), .B2(new_n959), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(G305), .B2(G1981), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n674), .A2(KEYINPUT114), .A3(new_n677), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n981));
  NAND3_X1  g556(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n674), .B2(new_n677), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n981), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n978), .A2(new_n979), .B1(new_n982), .B2(new_n984), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT49), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n944), .A2(KEYINPUT113), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n829), .A2(new_n990), .A3(new_n943), .ZN(new_n991));
  AND2_X1   g566(.A1(G160), .A2(G40), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n986), .A2(new_n988), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n564), .A2(new_n998), .A3(new_n565), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n980), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n996), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n564), .A2(G1976), .A3(new_n565), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1003), .A2(G8), .A3(new_n993), .A4(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n993), .A2(G8), .A3(new_n1004), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT52), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n997), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G303), .A2(G8), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT55), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n499), .A2(new_n943), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n989), .A2(new_n991), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n1014), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1017), .A2(G2090), .A3(new_n947), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n945), .A2(G1384), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n947), .B1(new_n829), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1013), .A2(new_n945), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1971), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(G8), .B(new_n1012), .C1(new_n1018), .C2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1001), .A2(new_n1002), .B1(new_n1009), .B2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1025));
  AND3_X1   g600(.A1(new_n829), .A2(new_n990), .A3(new_n943), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n990), .B1(new_n829), .B2(new_n943), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT50), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1013), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n947), .B1(new_n1029), .B2(new_n1014), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G2090), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1022), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1011), .B1(new_n1033), .B2(new_n995), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(new_n1023), .A3(new_n997), .A4(new_n1008), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT45), .B1(new_n989), .B2(new_n991), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n499), .A2(new_n1019), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n992), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n734), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n947), .A2(G2084), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT50), .B1(new_n989), .B2(new_n991), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(new_n1015), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(G8), .A3(G168), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1025), .B1(new_n1035), .B2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n997), .A2(new_n1008), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1011), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1047), .A2(new_n1023), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1024), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n945), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n947), .B1(new_n499), .B2(new_n1019), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1966), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1014), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1015), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1040), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT121), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1039), .A2(new_n1043), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(new_n1062), .A3(G168), .ZN(new_n1063));
  AND2_X1   g638(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1044), .A2(G8), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(G8), .A3(G286), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1063), .A2(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n995), .B(G168), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT62), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT119), .B1(new_n1017), .B2(new_n947), .ZN(new_n1077));
  INV_X1    g652(.A(G1961), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n992), .C1(new_n1042), .C2(new_n1015), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G2078), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1054), .A2(KEYINPUT53), .A3(new_n1082), .A4(new_n1055), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(G2078), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1081), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G171), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1035), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1073), .A2(new_n1076), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1053), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1081), .A2(G301), .A3(new_n1083), .A4(new_n1086), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1020), .A2(KEYINPUT53), .A3(new_n1082), .A4(new_n946), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1081), .A2(new_n1086), .A3(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT54), .B(new_n1092), .C1(new_n1094), .C2(G301), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1035), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1348), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1077), .A2(new_n1099), .A3(new_n1080), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n993), .A2(KEYINPUT118), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n989), .A2(new_n1102), .A3(new_n991), .A4(new_n992), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n939), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n596), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1100), .A2(new_n1105), .A3(KEYINPUT60), .A4(new_n587), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n592), .A2(KEYINPUT57), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n553), .A2(new_n555), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n551), .A2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(G1956), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1020), .A2(new_n1021), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1114), .B(new_n1118), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1118), .B1(G299), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1020), .A2(new_n1021), .A3(new_n1120), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1124), .B(new_n1125), .C1(new_n1031), .C2(G1956), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(new_n1126), .A3(KEYINPUT61), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1122), .A2(new_n1126), .A3(KEYINPUT120), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1122), .B2(KEYINPUT120), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1127), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT58), .B(G1341), .Z(new_n1132));
  NAND3_X1  g707(.A1(new_n1101), .A2(new_n1103), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1020), .A2(new_n953), .A3(new_n1021), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n539), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT59), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1113), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n587), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1122), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1126), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1098), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1081), .A2(G301), .A3(new_n1086), .A4(new_n1093), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1088), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT123), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1148), .A3(new_n1145), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1091), .B1(new_n1142), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n971), .B1(G1986), .B2(G290), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n950), .B1(new_n968), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n976), .B1(new_n1151), .B2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g729(.A1(new_n925), .A2(new_n929), .ZN(new_n1156));
  INV_X1    g730(.A(G319), .ZN(new_n1157));
  NOR3_X1   g731(.A1(G401), .A2(new_n1157), .A3(G227), .ZN(new_n1158));
  OAI21_X1  g732(.A(new_n1158), .B1(new_n669), .B2(new_n670), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n1159), .A2(KEYINPUT126), .ZN(new_n1160));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n1161));
  OAI211_X1 g735(.A(new_n1161), .B(new_n1158), .C1(new_n669), .C2(new_n670), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g737(.A1(new_n1156), .A2(new_n862), .A3(new_n1163), .ZN(G225));
  INV_X1    g738(.A(G225), .ZN(G308));
endmodule


