//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1148, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1203,
    new_n1204;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n203), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n210), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n202), .A2(new_n203), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT64), .ZN(new_n229));
  INV_X1    g0029(.A(G13), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n229), .B1(new_n207), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n232));
  AND2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OR3_X1    g0033(.A1(new_n228), .A2(new_n208), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n213), .A2(new_n225), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n220), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G58), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  OAI21_X1  g0053(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n254), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n256), .B1(new_n261), .B2(G226), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n257), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n264), .A2(new_n265), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n267), .A2(G223), .B1(G77), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G222), .ZN(new_n270));
  XOR2_X1   g0070(.A(KEYINPUT68), .B(G1698), .Z(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n266), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n269), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n231), .A2(new_n232), .B1(G33), .B2(G41), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(new_n273), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n262), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n278), .A2(G200), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n280));
  INV_X1    g0080(.A(G190), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n231), .A2(new_n232), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(G33), .B2(new_n209), .ZN(new_n285));
  AND2_X1   g0085(.A1(KEYINPUT8), .A2(G58), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT8), .A2(G58), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n208), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n288), .A2(new_n290), .B1(G150), .B2(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n292), .A2(KEYINPUT70), .B1(G20), .B2(new_n204), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n285), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n230), .A2(new_n208), .A3(G1), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n201), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n207), .A2(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n285), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n300), .B2(new_n201), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(KEYINPUT71), .B2(new_n295), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT73), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(KEYINPUT9), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n296), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n303), .A2(KEYINPUT9), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n283), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n283), .B(new_n307), .C1(KEYINPUT74), .C2(KEYINPUT10), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n278), .A2(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n296), .A2(new_n302), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n278), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n310), .A2(new_n311), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n297), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n285), .A2(G68), .A3(new_n318), .A4(new_n299), .ZN(new_n319));
  XOR2_X1   g0119(.A(new_n319), .B(KEYINPUT76), .Z(new_n320));
  NAND2_X1  g0120(.A1(new_n209), .A2(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n233), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n291), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n323));
  INV_X1    g0123(.A(G77), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n289), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n297), .A2(new_n203), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT12), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n327), .A2(KEYINPUT12), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n326), .A2(KEYINPUT11), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n320), .B(new_n330), .C1(KEYINPUT11), .C2(new_n326), .ZN(new_n331));
  INV_X1    g0131(.A(new_n256), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n260), .B2(new_n215), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT75), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n266), .A2(G1698), .ZN(new_n337));
  INV_X1    g0137(.A(G226), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n336), .B1(new_n337), .B2(new_n220), .C1(new_n272), .C2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n339), .B2(new_n276), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n340), .A2(new_n341), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT14), .B1(new_n345), .B2(new_n314), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(G179), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n345), .A2(KEYINPUT14), .A3(new_n314), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n331), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n331), .B1(new_n345), .B2(G190), .ZN(new_n351));
  OAI21_X1  g0151(.A(G200), .B1(new_n343), .B2(new_n344), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n256), .B1(new_n261), .B2(G244), .ZN(new_n355));
  INV_X1    g0155(.A(G107), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n337), .A2(new_n215), .B1(new_n356), .B2(new_n266), .ZN(new_n357));
  OR3_X1    g0157(.A1(new_n272), .A2(KEYINPUT72), .A3(new_n220), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT72), .B1(new_n272), .B2(new_n220), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n276), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(new_n281), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n297), .A2(new_n324), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n300), .B2(new_n324), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n288), .A2(new_n291), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT15), .B(G87), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(new_n208), .B2(new_n324), .C1(new_n289), .C2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n365), .B1(new_n322), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n362), .A2(G200), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n369), .B1(new_n362), .B2(new_n314), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n362), .A2(G179), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n317), .A2(new_n354), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n233), .A2(new_n321), .A3(new_n318), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n288), .A2(new_n299), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n379), .A2(new_n380), .B1(new_n318), .B2(new_n288), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT78), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n264), .A2(new_n208), .A3(new_n265), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT7), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n264), .A2(new_n386), .A3(new_n208), .A4(new_n265), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(G68), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(G58), .B(G68), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(G20), .B1(G159), .B2(new_n291), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(KEYINPUT16), .A3(new_n390), .ZN(new_n394));
  AND4_X1   g0194(.A1(KEYINPUT77), .A2(new_n393), .A3(new_n394), .A4(new_n322), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n285), .B1(new_n391), .B2(new_n392), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT77), .B1(new_n396), .B2(new_n394), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n383), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT79), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(KEYINPUT79), .B(new_n383), .C1(new_n395), .C2(new_n397), .ZN(new_n401));
  OR2_X1    g0201(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n402));
  NAND2_X1  g0202(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(G223), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G226), .A2(G1698), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n268), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n257), .A2(new_n216), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n276), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n256), .B1(new_n261), .B2(G232), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  MUX2_X1   g0210(.A(G179), .B(G169), .S(new_n410), .Z(new_n411));
  NAND3_X1  g0211(.A1(new_n400), .A2(new_n401), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT18), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n400), .A2(new_n401), .A3(new_n414), .A4(new_n411), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n408), .A2(G190), .A3(new_n409), .ZN(new_n416));
  INV_X1    g0216(.A(G200), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n408), .B2(new_n409), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n383), .C1(new_n395), .C2(new_n397), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT17), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n413), .A2(new_n415), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n378), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT82), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT5), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT81), .B1(new_n425), .B2(G41), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT81), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n258), .A3(KEYINPUT5), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(G41), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G45), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(G1), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n259), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n424), .B1(new_n434), .B2(new_n222), .ZN(new_n435));
  INV_X1    g0235(.A(new_n259), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n430), .B2(new_n432), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(KEYINPUT82), .A3(G257), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n272), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(KEYINPUT4), .A3(G244), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n267), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT4), .ZN(new_n443));
  INV_X1    g0243(.A(G244), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n272), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n276), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n430), .A2(G274), .A3(new_n259), .A4(new_n432), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n439), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G169), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n439), .A2(new_n447), .A3(G179), .A4(new_n448), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n379), .B1(new_n207), .B2(G33), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT80), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n318), .B2(G97), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n297), .A2(KEYINPUT80), .A3(new_n221), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n452), .A2(G97), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n356), .A2(KEYINPUT6), .A3(G97), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n221), .A2(new_n356), .ZN(new_n458));
  NOR2_X1   g0258(.A1(G97), .A2(G107), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n460), .B2(KEYINPUT6), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n461), .A2(G20), .B1(G77), .B2(new_n291), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n385), .A2(G107), .A3(new_n387), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n322), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n456), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT85), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT85), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n456), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n450), .A2(new_n451), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n439), .A2(new_n447), .A3(new_n448), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n466), .B1(new_n471), .B2(G190), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n449), .A2(KEYINPUT83), .A3(G200), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT83), .B1(new_n449), .B2(G200), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT84), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n472), .B(KEYINPUT84), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n266), .A2(new_n208), .A3(G87), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT22), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n481), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT23), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(new_n356), .A3(G20), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n289), .ZN(new_n489));
  XOR2_X1   g0289(.A(new_n489), .B(KEYINPUT90), .Z(new_n490));
  NAND2_X1  g0290(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(KEYINPUT24), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT24), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n484), .B2(new_n490), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n322), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT25), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n318), .B2(G107), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n356), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n452), .A2(G107), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G294), .ZN(new_n501));
  OAI221_X1 g0301(.A(new_n501), .B1(new_n337), .B2(new_n222), .C1(new_n272), .C2(new_n217), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(new_n276), .B1(G264), .B2(new_n437), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n448), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n314), .ZN(new_n505));
  INV_X1    g0305(.A(G179), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n506), .A3(new_n448), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n432), .A2(G274), .ZN(new_n511));
  OAI21_X1  g0311(.A(G250), .B1(new_n431), .B2(G1), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n436), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  OAI221_X1 g0314(.A(new_n514), .B1(new_n337), .B2(new_n444), .C1(new_n272), .C2(new_n215), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n513), .B1(new_n515), .B2(new_n276), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT86), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(KEYINPUT86), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n506), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n516), .A2(KEYINPUT86), .ZN(new_n522));
  AOI211_X1 g0322(.A(new_n518), .B(new_n513), .C1(new_n515), .C2(new_n276), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n314), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n525));
  XOR2_X1   g0325(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n526));
  NAND2_X1  g0326(.A1(new_n335), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n525), .B1(new_n527), .B2(new_n208), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n266), .A2(new_n208), .A3(G68), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n289), .A2(new_n221), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n322), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n367), .A2(new_n297), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT88), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n285), .B(new_n318), .C1(G1), .C2(new_n257), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n367), .ZN(new_n537));
  OR3_X1    g0337(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n535), .B1(new_n534), .B2(new_n537), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n521), .A2(new_n524), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n519), .A2(G190), .A3(new_n520), .ZN(new_n541));
  OAI21_X1  g0341(.A(G200), .B1(new_n522), .B2(new_n523), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n534), .B1(G87), .B2(new_n452), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n503), .A2(G190), .A3(new_n448), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n504), .A2(G200), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n495), .A2(new_n499), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n510), .A2(new_n540), .A3(new_n544), .A4(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n230), .A2(G1), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n208), .A2(G116), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n257), .A2(G97), .ZN(new_n552));
  AOI21_X1  g0352(.A(G20), .B1(G33), .B2(G283), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n322), .A2(KEYINPUT20), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT20), .B1(new_n322), .B2(new_n554), .ZN(new_n556));
  OAI221_X1 g0356(.A(new_n551), .B1(new_n555), .B2(new_n556), .C1(new_n488), .C2(new_n536), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n437), .A2(G270), .ZN(new_n558));
  XNOR2_X1  g0358(.A(KEYINPUT89), .B(G303), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n267), .A2(G264), .B1(new_n268), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n440), .A2(G257), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n448), .B(new_n558), .C1(new_n562), .C2(new_n361), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n557), .B1(G200), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n281), .B2(new_n563), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n557), .A2(new_n563), .A3(G169), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n557), .A2(new_n563), .A3(KEYINPUT21), .A4(G169), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n563), .A2(new_n506), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n557), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n565), .A2(new_n568), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n548), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n423), .A2(new_n479), .A3(new_n573), .ZN(G372));
  NAND3_X1  g0374(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n499), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n491), .B(KEYINPUT24), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(new_n322), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n579), .A2(new_n508), .A3(KEYINPUT91), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT91), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n500), .B2(new_n509), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n576), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n517), .A2(new_n314), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n521), .A2(new_n539), .A3(new_n538), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n517), .A2(G200), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n541), .A2(new_n543), .A3(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n585), .A2(new_n547), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n479), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n470), .A2(new_n540), .A3(new_n544), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n590), .A2(KEYINPUT26), .ZN(new_n591));
  INV_X1    g0391(.A(new_n466), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n450), .B2(new_n451), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n585), .A2(new_n593), .A3(new_n587), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n585), .B1(new_n594), .B2(KEYINPUT26), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n423), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT92), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n398), .A2(new_n411), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n600), .B(KEYINPUT18), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n353), .A2(new_n376), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n350), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n604), .B2(new_n421), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n310), .A2(new_n311), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n316), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT93), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(KEYINPUT93), .B(new_n316), .C1(new_n605), .C2(new_n606), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n599), .A2(new_n611), .ZN(G369));
  NAND2_X1  g0412(.A1(new_n549), .A2(new_n208), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(G213), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n616), .B(KEYINPUT94), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT95), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n618), .A2(G343), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(G343), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n622), .A2(new_n557), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT96), .B1(new_n575), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n572), .B2(new_n623), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n575), .A2(KEYINPUT96), .A3(new_n623), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G330), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n622), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n510), .B(new_n547), .C1(new_n579), .C2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n510), .B2(new_n631), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n575), .A2(new_n510), .A3(new_n547), .A4(new_n631), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n580), .A2(new_n582), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n622), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n635), .A2(new_n638), .ZN(G399));
  INV_X1    g0439(.A(new_n211), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G41), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n525), .A2(new_n488), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n641), .A2(new_n642), .A3(new_n207), .ZN(new_n643));
  INV_X1    g0443(.A(new_n227), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(new_n641), .ZN(new_n645));
  XOR2_X1   g0445(.A(new_n645), .B(KEYINPUT28), .Z(new_n646));
  INV_X1    g0446(.A(KEYINPUT29), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n594), .A2(KEYINPUT26), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n470), .A2(new_n540), .A3(new_n649), .A4(new_n544), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n585), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT97), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n576), .A2(new_n510), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n479), .A2(new_n588), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT97), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n648), .A2(new_n655), .A3(new_n585), .A4(new_n650), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n647), .B1(new_n657), .B2(new_n631), .ZN(new_n658));
  AOI211_X1 g0458(.A(KEYINPUT29), .B(new_n622), .C1(new_n589), .C2(new_n596), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n573), .A2(new_n479), .A3(new_n631), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n522), .A2(new_n523), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n570), .A2(new_n662), .A3(new_n471), .A4(new_n503), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT30), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n506), .A2(new_n563), .A3(new_n504), .A4(new_n517), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n663), .A2(new_n664), .B1(new_n665), .B2(new_n449), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n471), .A2(new_n503), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(KEYINPUT30), .A3(new_n570), .A4(new_n662), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n622), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT31), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n631), .B1(new_n666), .B2(new_n668), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT31), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n661), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n660), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n646), .B1(new_n678), .B2(G1), .ZN(G364));
  NOR2_X1   g0479(.A1(new_n230), .A2(G20), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n207), .B1(new_n680), .B2(G45), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n641), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n629), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n627), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(G330), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(G13), .A2(G33), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G20), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n640), .A2(new_n268), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n692), .A2(G355), .B1(new_n488), .B2(new_n640), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n640), .A2(new_n266), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n228), .B2(G45), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n252), .A2(new_n431), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n233), .B1(G20), .B2(new_n314), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n689), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n506), .A2(G200), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n208), .A2(G190), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n281), .A2(G179), .A3(G200), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n208), .ZN(new_n705));
  OAI221_X1 g0505(.A(new_n266), .B1(new_n703), .B2(new_n324), .C1(new_n705), .C2(new_n221), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n208), .A2(new_n281), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n506), .A2(new_n417), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n417), .A2(G179), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n702), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n710), .A2(G50), .B1(new_n713), .B2(G107), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n707), .A2(new_n701), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n708), .A2(new_n702), .ZN(new_n716));
  OAI221_X1 g0516(.A(new_n714), .B1(new_n202), .B2(new_n715), .C1(new_n203), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n707), .A2(new_n711), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT99), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(KEYINPUT99), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n706), .B(new_n717), .C1(G87), .C2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n702), .A2(new_n506), .A3(new_n417), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT98), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G159), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT32), .ZN(new_n731));
  INV_X1    g0531(.A(G283), .ZN(new_n732));
  INV_X1    g0532(.A(G311), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n712), .A2(new_n732), .B1(new_n703), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n266), .B1(new_n710), .B2(G326), .ZN(new_n735));
  INV_X1    g0535(.A(G294), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(new_n705), .ZN(new_n737));
  INV_X1    g0537(.A(new_n715), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n734), .B(new_n737), .C1(G322), .C2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G329), .ZN(new_n740));
  INV_X1    g0540(.A(G303), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n740), .A2(new_n728), .B1(new_n721), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(KEYINPUT33), .B(G317), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT100), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n716), .B1(new_n744), .B2(KEYINPUT100), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n723), .A2(new_n731), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n698), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n700), .B(new_n683), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n686), .B1(new_n691), .B2(new_n750), .ZN(G396));
  NOR2_X1   g0551(.A1(new_n631), .A2(new_n369), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT103), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n375), .B1(new_n753), .B2(new_n372), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n375), .A2(new_n622), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n688), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n733), .A2(new_n728), .B1(new_n721), .B2(new_n356), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n709), .A2(new_n741), .B1(new_n716), .B2(new_n732), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n713), .A2(G87), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(new_n736), .B2(new_n715), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n268), .B1(new_n703), .B2(new_n488), .C1(new_n705), .C2(new_n221), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n760), .A2(new_n761), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n712), .A2(new_n203), .ZN(new_n766));
  INV_X1    g0566(.A(new_n705), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(G58), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n716), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G137), .A2(new_n710), .B1(new_n769), .B2(G150), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G143), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n715), .A2(new_n772), .B1(new_n703), .B2(new_n729), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(KEYINPUT101), .B(KEYINPUT34), .Z(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n768), .B1(new_n201), .B2(new_n721), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n776), .B2(new_n774), .ZN(new_n778));
  INV_X1    g0578(.A(G132), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n266), .B1(new_n728), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT102), .Z(new_n781));
  AOI21_X1  g0581(.A(new_n765), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n749), .A2(new_n688), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n749), .B1(G77), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n683), .B1(new_n759), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n622), .B1(new_n589), .B2(new_n596), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(new_n757), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(new_n676), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n785), .B1(new_n788), .B2(new_n683), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT104), .ZN(G384));
  NOR2_X1   g0590(.A1(new_n680), .A2(new_n207), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n400), .A2(new_n401), .A3(new_n617), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT37), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n420), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n412), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n393), .A2(new_n394), .A3(new_n322), .ZN(new_n796));
  INV_X1    g0596(.A(new_n381), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n411), .B2(new_n617), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n420), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(KEYINPUT37), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT105), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n798), .A2(new_n617), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n422), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n795), .A2(KEYINPUT105), .A3(new_n801), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT38), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT106), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n808), .A2(KEYINPUT106), .A3(new_n809), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n804), .A2(new_n806), .A3(KEYINPUT38), .A4(new_n807), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OR3_X1    g0615(.A1(new_n673), .A2(KEYINPUT108), .A3(KEYINPUT31), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT108), .B1(new_n673), .B2(KEYINPUT31), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n816), .A2(new_n661), .A3(new_n817), .A4(new_n674), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n331), .A2(new_n622), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n354), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n331), .B(new_n622), .C1(new_n348), .C2(new_n349), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n818), .A2(new_n822), .A3(new_n758), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT40), .B1(new_n815), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT107), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n420), .A2(new_n825), .B1(new_n398), .B2(new_n411), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n792), .B(new_n826), .C1(new_n825), .C2(new_n420), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n412), .A2(new_n794), .ZN(new_n828));
  AOI22_X1  g0628(.A1(KEYINPUT37), .A2(new_n827), .B1(new_n828), .B2(new_n792), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n792), .B1(new_n601), .B2(new_n421), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n809), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n814), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n823), .A2(KEYINPUT40), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n824), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n423), .A2(new_n818), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n628), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT109), .Z(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n601), .A2(new_n617), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n755), .B1(new_n786), .B2(new_n758), .ZN(new_n841));
  INV_X1    g0641(.A(new_n822), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n840), .B1(new_n843), .B2(new_n815), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n815), .B2(KEYINPUT39), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n350), .A2(new_n622), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n423), .B1(new_n658), .B2(new_n659), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n611), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n848), .B(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n791), .B1(new_n839), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n839), .B2(new_n851), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n233), .A2(new_n208), .A3(new_n488), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n461), .A2(KEYINPUT35), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n461), .A2(KEYINPUT35), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT36), .ZN(new_n858));
  OAI21_X1  g0658(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n227), .A2(new_n859), .B1(G50), .B2(new_n203), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(G1), .A3(new_n230), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n853), .A2(new_n858), .A3(new_n861), .ZN(G367));
  OAI21_X1  g0662(.A(new_n479), .B1(new_n592), .B2(new_n631), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n593), .A2(new_n622), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n636), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n510), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n631), .B1(new_n868), .B2(new_n470), .ZN(new_n869));
  OR3_X1    g0669(.A1(new_n585), .A2(new_n543), .A3(new_n631), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n585), .B(new_n587), .C1(new_n543), .C2(new_n631), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n867), .A2(new_n869), .B1(KEYINPUT43), .B2(new_n872), .ZN(new_n873));
  OR3_X1    g0673(.A1(new_n873), .A2(KEYINPUT43), .A3(new_n872), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(KEYINPUT43), .B2(new_n872), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n635), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n877), .B2(new_n865), .ZN(new_n878));
  INV_X1    g0678(.A(new_n865), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n874), .A2(new_n635), .A3(new_n879), .A4(new_n875), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n641), .B(KEYINPUT41), .Z(new_n881));
  NAND2_X1  g0681(.A1(new_n865), .A2(new_n638), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT44), .Z(new_n883));
  NOR2_X1   g0683(.A1(new_n865), .A2(new_n638), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT45), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n877), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n877), .A3(new_n885), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n576), .A2(new_n622), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n636), .B1(new_n633), .B2(new_n889), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n629), .B(new_n890), .Z(new_n891));
  NOR2_X1   g0691(.A1(new_n677), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n881), .B1(new_n893), .B2(new_n678), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n878), .B(new_n880), .C1(new_n682), .C2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n694), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n240), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n699), .B1(new_n211), .B2(new_n367), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n683), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n769), .A2(G159), .B1(new_n713), .B2(G77), .ZN(new_n900));
  INV_X1    g0700(.A(G150), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n900), .B1(new_n772), .B2(new_n709), .C1(new_n901), .C2(new_n715), .ZN(new_n902));
  INV_X1    g0702(.A(G137), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n903), .A2(new_n728), .B1(new_n721), .B2(new_n202), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n767), .A2(G68), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(new_n266), .C1(new_n201), .C2(new_n703), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n902), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT110), .Z(new_n908));
  OAI221_X1 g0708(.A(new_n268), .B1(new_n703), .B2(new_n732), .C1(new_n705), .C2(new_n356), .ZN(new_n909));
  INV_X1    g0709(.A(new_n559), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n910), .A2(new_n715), .B1(new_n716), .B2(new_n736), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n709), .A2(new_n733), .B1(new_n712), .B2(new_n221), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(G317), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n914), .B2(new_n728), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n721), .A2(new_n488), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT46), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n908), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT47), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n899), .B1(new_n919), .B2(new_n698), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n872), .B2(new_n690), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n895), .A2(new_n921), .ZN(G387));
  INV_X1    g0722(.A(new_n891), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n634), .A2(new_n689), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n244), .A2(new_n431), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT111), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n288), .A2(new_n201), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT50), .Z(new_n928));
  AOI211_X1 g0728(.A(G45), .B(new_n642), .C1(G68), .C2(G77), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n896), .B(new_n926), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n692), .A2(new_n642), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(G107), .B2(new_n211), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n699), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n683), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n722), .A2(G77), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n268), .B1(new_n713), .B2(G97), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n901), .C2(new_n728), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT112), .Z(new_n938));
  NOR2_X1   g0738(.A1(new_n705), .A2(new_n367), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n769), .A2(new_n288), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n201), .B2(new_n715), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n709), .A2(new_n729), .B1(new_n703), .B2(new_n203), .ZN(new_n942));
  NOR4_X1   g0742(.A1(new_n938), .A2(new_n939), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT113), .ZN(new_n944));
  INV_X1    g0744(.A(new_n703), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G317), .A2(new_n738), .B1(new_n945), .B2(new_n559), .ZN(new_n946));
  INV_X1    g0746(.A(G322), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n946), .B1(new_n733), .B2(new_n716), .C1(new_n947), .C2(new_n709), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT48), .Z(new_n949));
  OAI22_X1  g0749(.A1(new_n721), .A2(new_n736), .B1(new_n732), .B2(new_n705), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n950), .A2(KEYINPUT114), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(KEYINPUT114), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(KEYINPUT49), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(KEYINPUT49), .ZN(new_n955));
  INV_X1    g0755(.A(new_n728), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(G326), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n266), .B1(new_n713), .B2(G116), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n944), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n934), .B1(new_n960), .B2(new_n698), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n923), .A2(new_n682), .B1(new_n924), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n892), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n641), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n678), .A2(new_n923), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G393));
  INV_X1    g0766(.A(new_n888), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n963), .B1(new_n967), .B2(new_n886), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n893), .A3(new_n641), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT115), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n967), .B2(new_n886), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n887), .A2(KEYINPUT115), .A3(new_n888), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n972), .A3(new_n682), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n249), .A2(new_n896), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n699), .B1(new_n221), .B2(new_n211), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n683), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT51), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n709), .A2(new_n901), .B1(new_n715), .B2(new_n729), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n722), .A2(G68), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n977), .B2(new_n978), .C1(new_n772), .C2(new_n728), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G50), .A2(new_n769), .B1(new_n945), .B2(new_n288), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n767), .A2(G77), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n981), .A2(new_n266), .A3(new_n762), .A4(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n559), .A2(new_n769), .B1(new_n945), .B2(G294), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n266), .B1(new_n713), .B2(G107), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n984), .B(new_n985), .C1(new_n488), .C2(new_n705), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n709), .A2(new_n914), .B1(new_n715), .B2(new_n733), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT52), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n732), .B2(new_n721), .C1(new_n947), .C2(new_n728), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n980), .A2(new_n983), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n976), .B1(new_n990), .B2(new_n698), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n879), .B2(new_n690), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n969), .A2(new_n973), .A3(new_n992), .ZN(G390));
  INV_X1    g0793(.A(new_n845), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n847), .B1(new_n841), .B2(new_n842), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n808), .A2(KEYINPUT106), .A3(new_n809), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT106), .B1(new_n808), .B2(new_n809), .ZN(new_n997));
  INV_X1    g0797(.A(new_n814), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT39), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n994), .B(new_n995), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n832), .A2(new_n847), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n657), .A2(new_n631), .A3(new_n754), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n756), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1002), .B1(new_n1004), .B2(new_n822), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n822), .A2(new_n675), .A3(G330), .A4(new_n758), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1001), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1005), .B1(new_n846), .B2(new_n995), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n818), .A2(new_n822), .A3(G330), .A4(new_n758), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n681), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n846), .A2(new_n687), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n683), .B1(new_n783), .B2(new_n288), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G294), .A2(new_n956), .B1(new_n722), .B2(G87), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G283), .A2(new_n710), .B1(new_n945), .B2(G97), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G107), .A2(new_n769), .B1(new_n738), .B2(G116), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n266), .B(new_n766), .C1(G77), .C2(new_n767), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n722), .A2(G150), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT53), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(KEYINPUT54), .B(G143), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n266), .B1(new_n703), .B2(new_n1022), .C1(new_n705), .C2(new_n729), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n715), .A2(new_n779), .B1(new_n712), .B2(new_n201), .ZN(new_n1024));
  INV_X1    g0824(.A(G128), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n709), .A2(new_n1025), .B1(new_n716), .B2(new_n903), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(G125), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n1028), .B2(new_n728), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1019), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1014), .B1(new_n1030), .B2(new_n698), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1012), .B1(new_n1013), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n423), .A2(G330), .A3(new_n818), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n849), .A2(new_n611), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n842), .B1(new_n676), .B2(new_n757), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n1010), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n841), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n818), .A2(G330), .A3(new_n758), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n842), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1003), .A2(new_n756), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n1041), .A3(new_n1007), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1034), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1011), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1008), .B(new_n1043), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n641), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1032), .A2(new_n1047), .ZN(G378));
  NAND2_X1  g0848(.A1(new_n313), .A2(new_n617), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n317), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n317), .A2(new_n1049), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  OR3_X1    g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1053), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n687), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n683), .B1(new_n783), .B2(G50), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n935), .B1(new_n732), .B2(new_n728), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G116), .A2(new_n710), .B1(new_n769), .B2(G97), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n356), .B2(new_n715), .C1(new_n367), .C2(new_n703), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n713), .A2(G58), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n905), .A2(new_n258), .A3(new_n268), .A4(new_n1063), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1060), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT58), .Z(new_n1066));
  AOI21_X1  g0866(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n716), .A2(new_n779), .B1(new_n703), .B2(new_n903), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n709), .A2(new_n1028), .B1(new_n715), .B2(new_n1025), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(G150), .C2(new_n767), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n721), .B2(new_n1022), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(KEYINPUT59), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(KEYINPUT59), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n956), .A2(G124), .ZN(new_n1074));
  AOI211_X1 g0874(.A(G33), .B(G41), .C1(new_n713), .C2(G159), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1066), .B1(G50), .B2(new_n1067), .C1(new_n1072), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT116), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n749), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1059), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1058), .A2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT117), .Z(new_n1083));
  INV_X1    g0883(.A(KEYINPUT118), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n848), .A2(new_n1057), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n824), .A2(new_n833), .A3(new_n628), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n844), .B(new_n1056), .C1(new_n846), .C2(new_n847), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1086), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1084), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1086), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n847), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1056), .B1(new_n1094), .B2(new_n844), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1087), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1091), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(KEYINPUT118), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1090), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1083), .B1(new_n1100), .B2(new_n682), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1034), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1046), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(KEYINPUT57), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n641), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT119), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT119), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1107), .A3(new_n641), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT57), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1101), .B1(new_n1109), .B2(new_n1110), .ZN(G375));
  AND2_X1   g0911(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1034), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n881), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n1044), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n741), .A2(new_n728), .B1(new_n721), .B2(new_n221), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n268), .B1(new_n712), .B2(new_n324), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G116), .A2(new_n769), .B1(new_n945), .B2(G107), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n736), .B2(new_n709), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n939), .B1(G283), .B2(new_n738), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT120), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1063), .B(new_n266), .C1(new_n201), .C2(new_n705), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n716), .A2(new_n1022), .B1(new_n703), .B2(new_n901), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n709), .A2(new_n779), .B1(new_n715), .B2(new_n903), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G128), .A2(new_n956), .B1(new_n722), .B2(G159), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1120), .A2(new_n1122), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n683), .B1(G68), .B2(new_n783), .C1(new_n1128), .C2(new_n749), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n842), .B2(new_n687), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1112), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n682), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1115), .A2(new_n1132), .ZN(G381));
  NAND2_X1  g0933(.A1(new_n1100), .A2(new_n682), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1083), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1104), .A2(new_n1107), .A3(new_n641), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1107), .B1(new_n1104), .B2(new_n641), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1136), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(G378), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OR4_X1    g0945(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1146));
  OR4_X1    g0946(.A1(G387), .A2(new_n1145), .A3(G381), .A4(new_n1146), .ZN(G407));
  NAND3_X1  g0947(.A1(new_n619), .A2(new_n620), .A3(G213), .ZN(new_n1148));
  OAI211_X1 g0948(.A(G407), .B(G213), .C1(new_n1145), .C2(new_n1148), .ZN(G409));
  NAND2_X1  g0949(.A1(G375), .A2(G378), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1148), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n681), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1082), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n1047), .A3(new_n1032), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1100), .A2(new_n1114), .A3(new_n1103), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1151), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT60), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1113), .B1(new_n1160), .B2(new_n1043), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1112), .A2(KEYINPUT60), .A3(new_n1034), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n641), .A3(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(new_n1132), .B1(G384), .B2(KEYINPUT121), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(G384), .A2(KEYINPUT121), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1164), .B(new_n1165), .Z(new_n1166));
  NAND2_X1  g0966(.A1(new_n1151), .A2(G2897), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1159), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT61), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(G393), .B(G396), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT123), .Z(new_n1175));
  AND3_X1   g0975(.A1(new_n895), .A2(new_n921), .A3(G390), .ZN(new_n1176));
  AOI21_X1  g0976(.A(G390), .B1(new_n895), .B2(new_n921), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1176), .B(KEYINPUT125), .Z(new_n1179));
  OR2_X1    g0979(.A1(new_n1177), .A2(KEYINPUT124), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(KEYINPUT124), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1174), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1178), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1158), .B(new_n1166), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT122), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1157), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1148), .B1(new_n1187), .B2(new_n1155), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G375), .B2(G378), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(KEYINPUT122), .A3(new_n1166), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT63), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1186), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1189), .A2(KEYINPUT63), .A3(new_n1166), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1173), .A2(new_n1183), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT62), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT126), .B1(new_n1184), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT126), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1189), .A2(new_n1197), .A3(KEYINPUT62), .A4(new_n1166), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1186), .A2(new_n1190), .A3(new_n1195), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1172), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1194), .B1(new_n1201), .B2(new_n1183), .ZN(G405));
  NAND2_X1  g1002(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(new_n1166), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(new_n1183), .ZN(G402));
endmodule


