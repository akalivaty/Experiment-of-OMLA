//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  INV_X1    g000(.A(G134gat), .ZN(new_n202));
  NOR3_X1   g001(.A1(new_n202), .A2(KEYINPUT66), .A3(G127gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(KEYINPUT66), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G113gat), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT67), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT67), .B1(new_n207), .B2(new_n209), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT68), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n205), .B(new_n216), .C1(new_n212), .C2(new_n213), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(KEYINPUT2), .ZN(new_n223));
  INV_X1    g022(.A(G148gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G141gat), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT76), .B(G148gat), .Z(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G141gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n219), .B1(new_n228), .B2(new_n220), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n223), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n209), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n207), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n209), .A2(new_n232), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n211), .B(new_n204), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n239), .A3(new_n231), .A4(new_n236), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(KEYINPUT77), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n237), .A2(new_n242), .A3(KEYINPUT4), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n217), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n207), .A2(new_n209), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(new_n211), .A3(new_n210), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n216), .B1(new_n249), .B2(new_n205), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n236), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n252), .B(new_n223), .C1(new_n227), .C2(new_n229), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n241), .A2(new_n243), .A3(new_n244), .A4(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n230), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n237), .ZN(new_n259));
  INV_X1    g058(.A(new_n244), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n255), .A2(new_n244), .A3(new_n257), .ZN(new_n263));
  OR3_X1    g062(.A1(new_n237), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n238), .A2(KEYINPUT79), .A3(new_n240), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT0), .ZN(new_n269));
  XNOR2_X1  g068(.A(G57gat), .B(G85gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n262), .A2(new_n271), .A3(new_n266), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n267), .A2(KEYINPUT6), .A3(new_n272), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT23), .ZN(new_n284));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT24), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT24), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(G183gat), .A3(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n288), .B(new_n289), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n302), .B2(new_n294), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n297), .B1(new_n289), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n283), .A2(KEYINPUT26), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n290), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n285), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(new_n283), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G183gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n313), .ZN(new_n317));
  INV_X1    g116(.A(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n311), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G183gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT27), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n323), .A2(new_n311), .A3(G190gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n310), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n304), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n282), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n306), .A2(new_n309), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(KEYINPUT65), .ZN(new_n330));
  AOI21_X1  g129(.A(G190gat), .B1(new_n316), .B2(new_n313), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT28), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n329), .B1(new_n332), .B2(new_n324), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n300), .A2(new_n301), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n295), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT25), .B1(new_n335), .B2(new_n298), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n336), .A3(new_n297), .ZN(new_n337));
  INV_X1    g136(.A(new_n282), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT22), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n341), .A2(new_n342), .B1(G211gat), .B2(G218gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n343), .B(KEYINPUT73), .C1(new_n341), .C2(new_n342), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345));
  INV_X1    g144(.A(G211gat), .ZN(new_n346));
  INV_X1    g145(.A(G218gat), .ZN(new_n347));
  OAI22_X1  g146(.A1(new_n346), .A2(new_n347), .B1(KEYINPUT72), .B2(KEYINPUT22), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n341), .A2(new_n342), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n344), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G211gat), .B(G218gat), .Z(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n337), .A2(KEYINPUT75), .A3(new_n338), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT75), .B1(new_n337), .B2(new_n338), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n361), .B(new_n328), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n281), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT30), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n360), .A2(new_n365), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n281), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n367), .A3(new_n281), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n278), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT88), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n327), .A2(new_n251), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n337), .A2(new_n218), .A3(new_n236), .ZN(new_n378));
  INV_X1    g177(.A(G227gat), .ZN(new_n379));
  INV_X1    g178(.A(G233gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT33), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT70), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT70), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n386), .A3(new_n383), .ZN(new_n387));
  XNOR2_X1  g186(.A(G15gat), .B(G43gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G71gat), .B(G99gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n382), .B2(KEYINPUT32), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n385), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n381), .B1(new_n377), .B2(new_n378), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT34), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI211_X1 g194(.A(KEYINPUT34), .B(new_n381), .C1(new_n377), .C2(new_n378), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n382), .B(KEYINPUT32), .C1(new_n383), .C2(new_n390), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n392), .B2(new_n398), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n376), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n391), .A2(new_n387), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n386), .B1(new_n382), .B2(new_n383), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n397), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT88), .A3(new_n399), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n375), .A2(new_n409), .A3(KEYINPUT35), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n253), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n359), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G228gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n380), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n356), .A2(new_n411), .A3(new_n358), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n231), .B1(new_n417), .B2(new_n252), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n352), .A2(new_n357), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n344), .A2(new_n350), .A3(new_n355), .A4(new_n351), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n411), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n231), .B1(new_n422), .B2(new_n252), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n415), .B1(new_n424), .B2(new_n413), .ZN(new_n425));
  OAI21_X1  g224(.A(G22gat), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n356), .A2(new_n358), .B1(new_n411), .B2(new_n253), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n423), .A2(new_n427), .B1(new_n414), .B2(new_n380), .ZN(new_n428));
  INV_X1    g227(.A(G22gat), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n428), .B(new_n429), .C1(new_n418), .C2(new_n416), .ZN(new_n430));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT31), .B(G50gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n426), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n426), .A2(new_n436), .A3(new_n430), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  OAI211_X1 g237(.A(KEYINPUT80), .B(G22gat), .C1(new_n419), .C2(new_n425), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n433), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n439), .A2(new_n433), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n436), .A3(new_n430), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT81), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n435), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n410), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT71), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n407), .A2(new_n447), .A3(new_n399), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n401), .A2(KEYINPUT71), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n445), .A2(new_n450), .A3(new_n278), .A4(new_n374), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT35), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(KEYINPUT38), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n340), .B2(new_n361), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n359), .B(new_n328), .C1(new_n363), .C2(new_n364), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n281), .A2(new_n456), .ZN(new_n461));
  INV_X1    g260(.A(new_n281), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(new_n369), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT86), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n459), .B(new_n465), .C1(new_n366), .C2(new_n461), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n464), .A2(new_n371), .A3(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n467), .A2(KEYINPUT87), .A3(new_n277), .A4(new_n276), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n464), .A2(new_n371), .A3(new_n466), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n278), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n369), .A2(KEYINPUT37), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n455), .B1(new_n473), .B2(new_n463), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n468), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n435), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n438), .B1(new_n437), .B2(new_n440), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n442), .A2(KEYINPUT81), .A3(new_n443), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n372), .A2(new_n373), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n259), .A2(new_n260), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n481), .A2(KEYINPUT83), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(KEYINPUT83), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n265), .A2(new_n264), .A3(new_n255), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n260), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT84), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(KEYINPUT40), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n484), .A3(new_n260), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n488), .A2(new_n271), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n480), .A2(new_n493), .A3(new_n273), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n488), .A2(new_n271), .A3(new_n492), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n490), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n479), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n475), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n450), .A2(KEYINPUT36), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT36), .B1(new_n407), .B2(new_n399), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n445), .A2(KEYINPUT82), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n479), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n375), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n453), .B1(new_n498), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n510), .A2(G1gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G8gat), .ZN(new_n515));
  INV_X1    g314(.A(G8gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n511), .A2(new_n516), .A3(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G43gat), .B(G50gat), .Z(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  AND2_X1   g320(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G29gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n520), .B1(new_n527), .B2(KEYINPUT15), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n527), .A2(KEYINPUT15), .A3(new_n520), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n531), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n519), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n518), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n519), .A2(KEYINPUT90), .A3(new_n531), .A4(new_n533), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n538), .B2(new_n518), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n537), .B(KEYINPUT13), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n537), .A4(new_n539), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT12), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n542), .A2(new_n548), .A3(new_n549), .A4(new_n556), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT21), .ZN(new_n561));
  INV_X1    g360(.A(G64gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(G57gat), .ZN(new_n563));
  INV_X1    g362(.A(G57gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(G64gat), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT9), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  INV_X1    g366(.A(G71gat), .ZN(new_n568));
  INV_X1    g367(.A(G78gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n562), .B2(G57gat), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT92), .B1(new_n564), .B2(G64gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(new_n562), .A3(G57gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n564), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n573), .A2(new_n574), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT9), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n567), .B1(new_n570), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n571), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n519), .B1(new_n561), .B2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT20), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n583), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n582), .A2(new_n561), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT93), .Z(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT95), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n590), .B(KEYINPUT93), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n593), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n595), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n597), .B1(new_n595), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n589), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n595), .A2(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n596), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(new_n588), .A3(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  OR2_X1    g408(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n610));
  AND3_X1   g409(.A1(KEYINPUT96), .A2(KEYINPUT97), .A3(KEYINPUT7), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT97), .B1(KEYINPUT96), .B2(KEYINPUT7), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n609), .B1(KEYINPUT96), .B2(KEYINPUT7), .ZN(new_n614));
  NAND2_X1  g413(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(KEYINPUT96), .A2(KEYINPUT97), .A3(KEYINPUT7), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT8), .ZN(new_n622));
  OAI22_X1  g421(.A1(new_n621), .A2(new_n622), .B1(G85gat), .B2(G92gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(G99gat), .A2(G106gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n571), .A2(new_n581), .ZN(new_n629));
  INV_X1    g428(.A(new_n627), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n620), .A2(new_n630), .A3(new_n624), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n620), .B2(new_n624), .ZN(new_n633));
  AOI211_X1 g432(.A(new_n627), .B(new_n623), .C1(new_n613), .C2(new_n619), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n582), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT98), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n632), .A2(new_n635), .A3(new_n639), .A4(new_n636), .ZN(new_n640));
  NOR4_X1   g439(.A1(new_n634), .A2(new_n633), .A3(new_n582), .A4(new_n636), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT99), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n635), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(G120gat), .B(G148gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT100), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n647), .A2(new_n649), .A3(new_n654), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI22_X1  g457(.A1(new_n534), .A2(new_n535), .B1(new_n634), .B2(new_n633), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n633), .A2(new_n634), .ZN(new_n660));
  AND2_X1   g459(.A1(G232gat), .A2(G233gat), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n660), .A2(new_n538), .B1(KEYINPUT41), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(G190gat), .B(G218gat), .Z(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n659), .A2(new_n666), .A3(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n661), .A2(KEYINPUT41), .ZN(new_n669));
  XNOR2_X1  g468(.A(G134gat), .B(G162gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n665), .A2(new_n671), .A3(new_n667), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n608), .A2(new_n658), .A3(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n509), .A2(new_n560), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n278), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n480), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n682), .A2(KEYINPUT101), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n516), .B1(new_n677), .B2(new_n480), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n682), .B1(new_n688), .B2(new_n683), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n684), .B1(new_n687), .B2(new_n689), .ZN(G1325gat));
  INV_X1    g489(.A(new_n677), .ZN(new_n691));
  AOI211_X1 g490(.A(KEYINPUT102), .B(new_n500), .C1(new_n450), .C2(KEYINPUT36), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n502), .A2(KEYINPUT102), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G15gat), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n409), .A2(G15gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n691), .B2(new_n697), .ZN(G1326gat));
  NAND2_X1  g497(.A1(new_n477), .A2(new_n478), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n504), .B1(new_n699), .B2(new_n435), .ZN(new_n700));
  AOI211_X1 g499(.A(KEYINPUT82), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n677), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT43), .B(G22gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n410), .A2(new_n445), .B1(KEYINPUT35), .B2(new_n451), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n475), .A2(new_n497), .B1(new_n702), .B2(new_n375), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(new_n695), .ZN(new_n709));
  INV_X1    g508(.A(new_n675), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n706), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n607), .B1(new_n509), .B2(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n560), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n658), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n278), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n475), .A2(new_n497), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n719), .B(new_n502), .C1(new_n507), .C2(new_n506), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n715), .B1(new_n720), .B2(new_n453), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n710), .A2(new_n607), .A3(new_n658), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n721), .A2(new_n525), .A3(new_n678), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n718), .A2(new_n724), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n374), .A2(G36gat), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n721), .A2(new_n726), .A3(new_n722), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n509), .A2(new_n560), .A3(new_n722), .A4(new_n727), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT103), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n728), .A2(new_n730), .A3(KEYINPUT105), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G36gat), .B1(new_n717), .B2(new_n374), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n728), .A2(new_n730), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT104), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n738), .A2(KEYINPUT104), .A3(KEYINPUT46), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n736), .B(new_n737), .C1(new_n739), .C2(new_n740), .ZN(G1329gat));
  INV_X1    g540(.A(G43gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n721), .A2(new_n722), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(new_n409), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT102), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n499), .B2(new_n501), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n692), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n744), .B1(new_n717), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT47), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n744), .C1(new_n717), .C2(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1330gat));
  NAND3_X1  g552(.A1(new_n721), .A2(KEYINPUT106), .A3(new_n722), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n506), .A2(G50gat), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n743), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n711), .A2(new_n713), .A3(new_n479), .A4(new_n716), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G50gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(KEYINPUT48), .A3(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n711), .A2(new_n713), .A3(new_n702), .A4(new_n716), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n756), .A2(new_n758), .B1(G50gat), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(KEYINPUT48), .B2(new_n764), .ZN(G1331gat));
  NAND2_X1  g564(.A1(new_n708), .A2(new_n695), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n453), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768));
  INV_X1    g567(.A(new_n658), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n560), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n607), .A3(new_n710), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT107), .Z(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n767), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT108), .B1(new_n709), .B2(new_n772), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n278), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n564), .ZN(G1332gat));
  NAND2_X1  g577(.A1(new_n480), .A2(KEYINPUT109), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n374), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n562), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT110), .Z(new_n785));
  NAND3_X1  g584(.A1(new_n774), .A2(new_n775), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT111), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n774), .A2(new_n775), .A3(new_n788), .A4(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n783), .A2(new_n562), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1333gat));
  OAI21_X1  g591(.A(G71gat), .B1(new_n776), .B2(new_n695), .ZN(new_n793));
  INV_X1    g592(.A(new_n409), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n568), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n776), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n793), .B(KEYINPUT50), .C1(new_n776), .C2(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1334gat));
  NOR2_X1   g599(.A1(new_n776), .A2(new_n506), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(new_n569), .ZN(G1335gat));
  NAND2_X1  g601(.A1(new_n714), .A2(new_n770), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n278), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n710), .B1(new_n766), .B2(new_n453), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n608), .B1(KEYINPUT112), .B2(KEYINPUT51), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n560), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n811), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n805), .A2(new_n813), .A3(new_n807), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OR3_X1    g614(.A1(new_n278), .A2(G85gat), .A3(new_n769), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n804), .B1(new_n815), .B2(new_n816), .ZN(G1336gat));
  AOI21_X1  g616(.A(new_n813), .B1(new_n805), .B2(new_n807), .ZN(new_n818));
  INV_X1    g617(.A(new_n807), .ZN(new_n819));
  NOR4_X1   g618(.A1(new_n709), .A2(new_n710), .A3(new_n811), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI211_X1 g620(.A(G92gat), .B(new_n769), .C1(new_n779), .C2(new_n781), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n711), .A2(new_n713), .A3(new_n770), .A4(new_n782), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT114), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G92gat), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n824), .A2(KEYINPUT114), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n711), .A2(new_n713), .A3(new_n480), .A4(new_n770), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G92gat), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n822), .B(KEYINPUT113), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n815), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n828), .A2(new_n833), .ZN(G1337gat));
  OAI21_X1  g633(.A(G99gat), .B1(new_n803), .B2(new_n695), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n409), .A2(G99gat), .A3(new_n769), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n815), .B2(new_n836), .ZN(G1338gat));
  NOR3_X1   g636(.A1(new_n445), .A2(G106gat), .A3(new_n769), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT115), .Z(new_n839));
  NAND4_X1  g638(.A1(new_n812), .A2(new_n814), .A3(KEYINPUT116), .A4(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n711), .A2(new_n713), .A3(new_n702), .A4(new_n770), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G106gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n821), .A2(new_n839), .B1(KEYINPUT116), .B2(KEYINPUT53), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n711), .A2(new_n713), .A3(new_n479), .A4(new_n770), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(G106gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n844), .A2(new_n849), .ZN(G1339gat));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n641), .B1(new_n637), .B2(KEYINPUT98), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n852), .A2(new_n645), .A3(new_n640), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n645), .B1(new_n852), .B2(new_n640), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n655), .B1(new_n647), .B2(KEYINPUT54), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n851), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n654), .B1(new_n854), .B2(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n647), .A2(KEYINPUT54), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n859), .B(KEYINPUT55), .C1(new_n860), .C2(new_n853), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n858), .A2(new_n560), .A3(new_n657), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n546), .A2(new_n547), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n537), .B1(new_n536), .B2(new_n539), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n555), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(new_n559), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n675), .B1(new_n658), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n858), .A2(new_n657), .A3(new_n861), .A4(new_n866), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n675), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n870), .A3(new_n608), .ZN(new_n871));
  NOR4_X1   g670(.A1(new_n608), .A2(new_n658), .A3(new_n675), .A4(new_n560), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n506), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT117), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n782), .A2(new_n278), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n794), .A3(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(new_n208), .A3(new_n715), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n607), .B1(new_n869), .B2(new_n675), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n872), .B1(new_n880), .B2(new_n868), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n278), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n479), .B1(new_n449), .B2(new_n448), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n782), .ZN(new_n885));
  AOI21_X1  g684(.A(G113gat), .B1(new_n885), .B2(new_n560), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n879), .A2(new_n886), .ZN(G1340gat));
  OAI21_X1  g686(.A(G120gat), .B1(new_n878), .B2(new_n769), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n658), .A2(new_n206), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT118), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(G1341gat));
  OAI21_X1  g691(.A(G127gat), .B1(new_n878), .B2(new_n608), .ZN(new_n893));
  INV_X1    g692(.A(G127gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n885), .A2(new_n894), .A3(new_n607), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1342gat));
  OAI21_X1  g695(.A(G134gat), .B1(new_n878), .B2(new_n710), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n374), .A2(new_n675), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n884), .A2(G134gat), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT56), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(G1343gat));
  NOR2_X1   g700(.A1(new_n747), .A2(new_n445), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n882), .ZN(new_n903));
  NOR4_X1   g702(.A1(new_n903), .A2(G141gat), .A3(new_n715), .A4(new_n782), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n877), .B1(new_n746), .B2(new_n692), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n881), .A2(new_n506), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n874), .A2(KEYINPUT57), .A3(new_n702), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n907), .B1(new_n881), .B2(new_n445), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT119), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n560), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G141gat), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n905), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n911), .A2(KEYINPUT119), .A3(new_n912), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n874), .A2(new_n909), .A3(KEYINPUT57), .A4(new_n702), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n695), .A3(new_n877), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT120), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n910), .A2(new_n922), .A3(new_n913), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n560), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n904), .B1(new_n924), .B2(G141gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n917), .B1(new_n925), .B2(new_n916), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g727(.A(KEYINPUT121), .B(new_n917), .C1(new_n925), .C2(new_n916), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1344gat));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n921), .A2(new_n923), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(new_n658), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n931), .B1(new_n933), .B2(new_n226), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n907), .B1(new_n874), .B2(new_n479), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n881), .A2(new_n506), .A3(KEYINPUT57), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n769), .B1(new_n906), .B2(KEYINPUT122), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n937), .B(new_n938), .C1(KEYINPUT122), .C2(new_n906), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n931), .A2(new_n224), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n903), .A2(new_n782), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n658), .A2(new_n226), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n939), .A2(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n934), .A2(new_n943), .ZN(G1345gat));
  AOI21_X1  g743(.A(G155gat), .B1(new_n941), .B2(new_n607), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n607), .A2(G155gat), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT123), .Z(new_n947));
  AOI21_X1  g746(.A(new_n945), .B1(new_n932), .B2(new_n947), .ZN(G1346gat));
  NOR3_X1   g747(.A1(new_n903), .A2(G162gat), .A3(new_n898), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT124), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n932), .A2(new_n675), .ZN(new_n951));
  INV_X1    g750(.A(G162gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(G1347gat));
  NOR2_X1   g752(.A1(new_n881), .A2(new_n678), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(new_n883), .A3(new_n782), .ZN(new_n955));
  AOI21_X1  g754(.A(G169gat), .B1(new_n955), .B2(new_n560), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n678), .A2(new_n374), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n876), .A2(new_n794), .A3(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n560), .A2(G169gat), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1348gat));
  AOI21_X1  g760(.A(G176gat), .B1(new_n955), .B2(new_n658), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n658), .A2(G176gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n959), .B2(new_n963), .ZN(G1349gat));
  NAND3_X1  g763(.A1(new_n955), .A2(new_n312), .A3(new_n607), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969));
  AOI22_X1  g768(.A1(new_n967), .A2(new_n968), .B1(new_n969), .B2(KEYINPUT60), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n969), .A2(KEYINPUT60), .ZN(new_n971));
  OAI21_X1  g770(.A(G183gat), .B1(new_n958), .B2(new_n608), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n970), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(G1350gat));
  NAND3_X1  g774(.A1(new_n955), .A2(new_n318), .A3(new_n675), .ZN(new_n976));
  OAI21_X1  g775(.A(G190gat), .B1(new_n958), .B2(new_n710), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n977), .A2(KEYINPUT61), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n977), .A2(KEYINPUT61), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G1351gat));
  AND3_X1   g779(.A1(new_n902), .A2(new_n782), .A3(new_n954), .ZN(new_n981));
  AOI21_X1  g780(.A(G197gat), .B1(new_n981), .B2(new_n560), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n747), .A2(new_n678), .A3(new_n374), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n937), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n560), .A2(G197gat), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1352gat));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n987));
  AOI21_X1  g786(.A(G204gat), .B1(new_n987), .B2(KEYINPUT62), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n981), .A2(new_n658), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(new_n984), .ZN(new_n992));
  OAI21_X1  g791(.A(G204gat), .B1(new_n992), .B2(new_n769), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1353gat));
  NAND3_X1  g793(.A1(new_n981), .A2(new_n346), .A3(new_n607), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n984), .A2(new_n607), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n996), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n992), .B2(new_n710), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n981), .A2(new_n347), .A3(new_n675), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1355gat));
endmodule


