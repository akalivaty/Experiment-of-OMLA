//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT69), .B(G113gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  OR2_X1    g008(.A1(G113gat), .A2(G120gat), .ZN(new_n210));
  XOR2_X1   g009(.A(KEYINPUT70), .B(KEYINPUT1), .Z(new_n211));
  XNOR2_X1  g010(.A(G127gat), .B(G134gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(G127gat), .A2(G134gat), .ZN(new_n216));
  XOR2_X1   g015(.A(KEYINPUT68), .B(G134gat), .Z(new_n217));
  INV_X1    g016(.A(G127gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G141gat), .B(G148gat), .Z(new_n222));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  INV_X1    g025(.A(G162gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT74), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT74), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G155gat), .B2(G162gat), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n224), .A2(new_n225), .A3(new_n228), .A4(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n226), .B(new_n227), .C1(new_n223), .C2(KEYINPUT75), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n225), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n225), .A2(KEYINPUT2), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT75), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n222), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n213), .A2(new_n231), .A3(new_n219), .A4(new_n236), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT4), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n237), .A2(KEYINPUT3), .B1(new_n219), .B2(new_n213), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n231), .A2(new_n245), .A3(new_n236), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n207), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT39), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n206), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n220), .A2(new_n237), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(new_n207), .A3(new_n241), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n252), .A2(KEYINPUT77), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n249), .B1(new_n252), .B2(KEYINPUT77), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n240), .A2(new_n242), .B1(new_n244), .B2(new_n246), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n253), .B(new_n254), .C1(new_n255), .C2(new_n207), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(new_n256), .A3(KEYINPUT40), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT40), .B1(new_n250), .B2(new_n256), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(KEYINPUT78), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT78), .ZN(new_n260));
  AOI211_X1 g059(.A(new_n260), .B(KEYINPUT40), .C1(new_n250), .C2(new_n256), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G8gat), .B(G36gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G64gat), .B(G92gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT72), .B(G197gat), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n266), .A2(G204gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268));
  INV_X1    g067(.A(G211gat), .ZN(new_n269));
  INV_X1    g068(.A(G218gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(G204gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT73), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n273), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(KEYINPUT24), .ZN(new_n283));
  AND2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  INV_X1    g085(.A(G190gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT24), .A3(new_n282), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n281), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n279), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n293), .A2(KEYINPUT26), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n284), .B1(new_n293), .B2(KEYINPUT26), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n294), .A2(new_n295), .B1(G183gat), .B2(G190gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT27), .B(G183gat), .Z(new_n298));
  OAI21_X1  g097(.A(KEYINPUT65), .B1(new_n298), .B2(G190gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(new_n287), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n297), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n287), .A2(KEYINPUT28), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n296), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n292), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G226gat), .ZN(new_n310));
  INV_X1    g109(.A(G233gat), .ZN(new_n311));
  OAI22_X1  g110(.A1(new_n309), .A2(KEYINPUT29), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n308), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(G226gat), .A3(G233gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n278), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n313), .A2(new_n316), .B1(G226gat), .B2(G233gat), .ZN(new_n317));
  AOI211_X1 g116(.A(new_n310), .B(new_n311), .C1(new_n292), .C2(new_n308), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n317), .A2(new_n318), .A3(new_n277), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n265), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n312), .A2(new_n278), .A3(new_n314), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n277), .B1(new_n317), .B2(new_n318), .ZN(new_n322));
  INV_X1    g121(.A(new_n265), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(KEYINPUT30), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT30), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n321), .A2(new_n322), .A3(new_n326), .A4(new_n323), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT5), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n243), .A2(new_n207), .A3(new_n247), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n207), .B1(new_n251), .B2(new_n241), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n330), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT5), .B1(new_n255), .B2(new_n207), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n330), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n332), .B1(new_n255), .B2(new_n207), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n337), .B(KEYINPUT79), .C1(new_n338), .C2(new_n330), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n336), .A2(new_n206), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n262), .A2(new_n328), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT29), .B1(new_n273), .B2(new_n274), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n274), .B2(new_n273), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n238), .B1(new_n343), .B2(new_n245), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n246), .A2(new_n316), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n277), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G228gat), .ZN(new_n347));
  OAI22_X1  g146(.A1(new_n344), .A2(new_n346), .B1(new_n347), .B2(new_n311), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT76), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n346), .A2(new_n347), .A3(new_n311), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT3), .B1(new_n278), .B2(new_n316), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n238), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G78gat), .B(G106gat), .ZN(new_n354));
  INV_X1    g153(.A(G22gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT31), .B(G50gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n353), .B(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n337), .B1(new_n338), .B2(new_n330), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  INV_X1    g161(.A(new_n206), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT6), .B1(new_n361), .B2(new_n363), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n340), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT37), .B1(new_n315), .B2(new_n319), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT38), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT37), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n321), .A2(new_n322), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n367), .A2(new_n368), .A3(new_n265), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n367), .A2(new_n265), .A3(new_n370), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT38), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n366), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n372), .B1(new_n371), .B2(new_n324), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n341), .B(new_n360), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n360), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n365), .B1(new_n363), .B2(new_n361), .ZN(new_n380));
  INV_X1    g179(.A(new_n364), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n325), .A2(new_n327), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n313), .A2(new_n220), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n292), .A2(new_n308), .A3(new_n221), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G227gat), .A2(G233gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT64), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n387), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n221), .B1(new_n292), .B2(new_n308), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G15gat), .B(G43gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT33), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(KEYINPUT32), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT71), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT32), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n404), .B1(new_n388), .B2(new_n391), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT71), .A3(new_n400), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT34), .ZN(new_n408));
  INV_X1    g207(.A(new_n399), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n396), .B2(KEYINPUT32), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n407), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n408), .B1(new_n407), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n393), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT71), .B1(new_n405), .B2(new_n400), .ZN(new_n417));
  AND4_X1   g216(.A1(KEYINPUT71), .A2(new_n396), .A3(KEYINPUT32), .A4(new_n400), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT34), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n407), .A2(new_n408), .A3(new_n413), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n420), .A2(new_n392), .A3(new_n389), .A4(new_n421), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n416), .A2(KEYINPUT36), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT36), .B1(new_n416), .B2(new_n422), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n378), .B(new_n385), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n416), .A2(new_n360), .A3(new_n422), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n416), .A2(new_n360), .A3(new_n422), .A4(KEYINPUT82), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT35), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n384), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n340), .A2(new_n365), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n433), .B(new_n383), .C1(new_n434), .C2(new_n364), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT81), .B1(new_n366), .B2(new_n328), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n430), .B1(new_n437), .B2(new_n426), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n425), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  OR2_X1    g238(.A1(G71gat), .A2(G78gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(G71gat), .A2(G78gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G57gat), .B(G64gat), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(KEYINPUT91), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT9), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(KEYINPUT90), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n445), .ZN(new_n448));
  INV_X1    g247(.A(G64gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(G57gat), .ZN(new_n450));
  INV_X1    g249(.A(G57gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(G64gat), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n447), .A2(new_n448), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n444), .A2(new_n446), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n452), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT91), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n455), .A2(new_n456), .B1(new_n441), .B2(new_n440), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n448), .A2(new_n447), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n455), .A3(new_n446), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(KEYINPUT21), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT93), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n454), .A2(new_n460), .A3(KEYINPUT93), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n462), .B1(new_n466), .B2(KEYINPUT21), .ZN(new_n467));
  NOR2_X1   g266(.A1(G15gat), .A2(G22gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n470));
  NAND2_X1  g269(.A1(G15gat), .A2(G22gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT86), .B1(new_n473), .B2(new_n468), .ZN(new_n474));
  INV_X1    g273(.A(G1gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT16), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(G1gat), .B1(new_n472), .B2(new_n474), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n478), .A2(new_n479), .A3(G8gat), .ZN(new_n480));
  INV_X1    g279(.A(G8gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n474), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n475), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(new_n477), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  MUX2_X1   g284(.A(new_n462), .B(new_n467), .S(new_n485), .Z(new_n486));
  NAND2_X1  g285(.A1(G231gat), .A2(G233gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT92), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(new_n286), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(new_n269), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n486), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G127gat), .B(G155gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n491), .B(new_n494), .ZN(new_n495));
  OR3_X1    g294(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n496), .A2(new_n497), .B1(G29gat), .B2(G36gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(G43gat), .B(G50gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(KEYINPUT15), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505));
  INV_X1    g304(.A(G50gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(KEYINPUT84), .A3(G43gat), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(G43gat), .ZN(new_n509));
  INV_X1    g308(.A(G43gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G50gat), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n509), .A2(new_n511), .A3(new_n502), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n505), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT85), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n508), .A2(new_n514), .A3(new_n498), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n499), .A2(KEYINPUT15), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n501), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518));
  INV_X1    g317(.A(G92gat), .ZN(new_n519));
  AOI22_X1  g318(.A1(KEYINPUT8), .A2(new_n518), .B1(new_n203), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n203), .B2(new_n519), .ZN(new_n522));
  NAND3_X1  g321(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G99gat), .B(G106gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(G232gat), .A2(G233gat), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n517), .A2(new_n526), .B1(KEYINPUT41), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n526), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n517), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g330(.A(KEYINPUT17), .B(new_n501), .C1(new_n515), .C2(new_n516), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT95), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n533), .B(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n527), .A2(KEYINPUT41), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT94), .ZN(new_n538));
  XNOR2_X1  g337(.A(G134gat), .B(G162gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n495), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT96), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n454), .A2(new_n460), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(new_n454), .B2(new_n460), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n526), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT10), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n461), .A2(KEYINPUT96), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n529), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n464), .A2(KEYINPUT10), .A3(new_n465), .A4(new_n526), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n548), .A2(new_n551), .ZN(new_n557));
  INV_X1    g356(.A(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n556), .A2(new_n559), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n544), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G169gat), .B(G197gat), .Z(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT12), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n577));
  OAI21_X1  g376(.A(G8gat), .B1(new_n478), .B2(new_n479), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n483), .A2(new_n481), .A3(new_n477), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n577), .B1(new_n517), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n517), .A2(new_n580), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT13), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT88), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n485), .B1(new_n517), .B2(new_n530), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n584), .B(new_n582), .C1(new_n589), .C2(new_n532), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT87), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT18), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n590), .B2(new_n588), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n587), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI211_X1 g394(.A(new_n588), .B(new_n593), .C1(new_n590), .C2(new_n591), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n576), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n591), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT88), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n590), .A2(new_n588), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT18), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n592), .A2(KEYINPUT18), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n602), .A2(new_n575), .A3(new_n603), .A4(new_n587), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n569), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n439), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n382), .B(KEYINPUT97), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(new_n475), .ZN(G1324gat));
  NOR2_X1   g410(.A1(new_n608), .A2(new_n383), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT42), .B1(new_n612), .B2(new_n481), .ZN(new_n613));
  NAND2_X1  g412(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n614));
  OR2_X1    g413(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  MUX2_X1   g415(.A(KEYINPUT42), .B(new_n613), .S(new_n616), .Z(G1325gat));
  INV_X1    g416(.A(new_n608), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n423), .A2(new_n424), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n618), .A2(G15gat), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n416), .A2(new_n422), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(G15gat), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n623), .ZN(G1326gat));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n360), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT43), .B(G22gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(G1327gat));
  AND2_X1   g426(.A1(new_n439), .A2(new_n543), .ZN(new_n628));
  INV_X1    g427(.A(new_n495), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n629), .A2(new_n606), .A3(new_n567), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(G29gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n382), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT45), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n543), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT99), .B1(new_n541), .B2(new_n542), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(KEYINPUT44), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n439), .A2(KEYINPUT98), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n425), .A2(new_n432), .A3(new_n645), .A4(new_n438), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n439), .B2(new_n543), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n630), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n635), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n637), .B1(new_n654), .B2(new_n633), .ZN(G1328gat));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n328), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(G36gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n631), .A2(G36gat), .A3(new_n383), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT46), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(G1329gat));
  NAND3_X1  g459(.A1(new_n652), .A2(G43gat), .A3(new_n619), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n662), .A2(KEYINPUT47), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n632), .A2(new_n622), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n664), .A2(new_n510), .B1(new_n662), .B2(KEYINPUT47), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n661), .B2(new_n665), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(G1330gat));
  NOR3_X1   g467(.A1(new_n631), .A2(G50gat), .A3(new_n360), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n379), .B(new_n630), .C1(new_n647), .C2(new_n649), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n671), .A2(KEYINPUT102), .ZN(new_n672));
  OAI21_X1  g471(.A(G50gat), .B1(new_n671), .B2(KEYINPUT102), .ZN(new_n673));
  OAI211_X1 g472(.A(KEYINPUT48), .B(new_n670), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n671), .A2(new_n675), .A3(G50gat), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n671), .B2(G50gat), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n676), .A2(new_n677), .A3(new_n669), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n674), .B1(new_n678), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g478(.A1(new_n605), .A2(new_n568), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n544), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n644), .B2(new_n646), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n635), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n609), .A2(KEYINPUT103), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g487(.A(new_n383), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT104), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n691), .B(new_n692), .Z(G1333gat));
  NAND3_X1  g492(.A1(new_n682), .A2(G71gat), .A3(new_n619), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n682), .A2(new_n622), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(G71gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n379), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT105), .B(G78gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1335gat));
  NAND4_X1  g499(.A1(new_n439), .A2(new_n606), .A3(new_n495), .A4(new_n543), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT106), .B(KEYINPUT51), .Z(new_n702));
  OR2_X1    g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT51), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n609), .A2(G85gat), .A3(new_n568), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT107), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n680), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n629), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n647), .B2(new_n649), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n635), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n710), .B1(new_n716), .B2(new_n203), .ZN(G1336gat));
  NOR3_X1   g516(.A1(new_n383), .A2(new_n568), .A3(G92gat), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT52), .B1(new_n707), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G92gat), .B1(new_n713), .B2(new_n383), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n701), .A2(KEYINPUT108), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n705), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n701), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(new_n724), .A3(new_n718), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(G1337gat));
  INV_X1    g527(.A(G99gat), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n707), .A2(new_n729), .A3(new_n622), .A4(new_n567), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n619), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n732), .B2(new_n729), .ZN(G1338gat));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n379), .B(new_n712), .C1(new_n647), .C2(new_n649), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G106gat), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n360), .A2(G106gat), .A3(new_n568), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n707), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n738), .ZN(new_n740));
  AOI211_X1 g539(.A(KEYINPUT110), .B(new_n740), .C1(new_n703), .C2(new_n706), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n734), .B(new_n736), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n724), .A3(new_n738), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT109), .B1(new_n744), .B2(KEYINPUT53), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n746), .B(new_n734), .C1(new_n736), .C2(new_n743), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n742), .B1(new_n745), .B2(new_n747), .ZN(G1339gat));
  NOR2_X1   g547(.A1(new_n639), .A2(new_n640), .ZN(new_n749));
  INV_X1    g548(.A(new_n556), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n565), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n552), .A2(new_n558), .A3(new_n553), .ZN(new_n754));
  AND4_X1   g553(.A1(new_n753), .A2(new_n556), .A3(KEYINPUT54), .A4(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n751), .B1(new_n554), .B2(new_n555), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n753), .B1(new_n756), .B2(new_n754), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT55), .B(new_n752), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n566), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(KEYINPUT112), .A3(new_n566), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n752), .B1(new_n755), .B2(new_n757), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n761), .A2(new_n605), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n574), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n581), .B1(new_n517), .B2(new_n580), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n515), .A2(new_n516), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n500), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n770), .A2(new_n485), .A3(new_n577), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n585), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n582), .B1(new_n589), .B2(new_n532), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(G229gat), .A3(G233gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n772), .B2(KEYINPUT113), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n767), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n604), .A3(new_n567), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n749), .B1(new_n766), .B2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n777), .A2(new_n604), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n761), .A2(new_n780), .A3(new_n762), .A4(new_n765), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n641), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n495), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n544), .A2(new_n606), .A3(new_n568), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n379), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n609), .A2(new_n328), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n622), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G113gat), .B1(new_n787), .B2(new_n606), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n783), .A2(new_n784), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(new_n686), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n428), .A2(new_n429), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n383), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n606), .A2(new_n208), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n788), .B1(new_n794), .B2(new_n795), .ZN(G1340gat));
  OAI21_X1  g595(.A(G120gat), .B1(new_n787), .B2(new_n568), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n568), .A2(G120gat), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n794), .B2(new_n798), .ZN(G1341gat));
  NOR3_X1   g598(.A1(new_n787), .A2(new_n218), .A3(new_n495), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n793), .A2(new_n383), .A3(new_n629), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(G127gat), .B1(new_n801), .B2(new_n802), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(G1342gat));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n543), .A2(new_n383), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT115), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n217), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n806), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n543), .ZN(new_n816));
  OAI21_X1  g615(.A(G134gat), .B1(new_n787), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(KEYINPUT56), .A3(new_n812), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(new_n817), .A3(new_n819), .ZN(G1343gat));
  INV_X1    g619(.A(new_n619), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n786), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n379), .A2(KEYINPUT57), .ZN(new_n824));
  INV_X1    g623(.A(new_n781), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n605), .A2(new_n566), .A3(new_n765), .A4(new_n758), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n543), .B1(new_n826), .B2(new_n778), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n749), .A2(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n827), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT118), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n629), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n784), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n824), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT57), .B1(new_n789), .B2(new_n379), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT117), .B(KEYINPUT57), .C1(new_n789), .C2(new_n379), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n605), .B(new_n823), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G141gat), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n619), .A2(new_n360), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n790), .A2(new_n383), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n606), .A2(G141gat), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT58), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n840), .A2(new_n848), .A3(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1344gat));
  INV_X1    g649(.A(G148gat), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(KEYINPUT59), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n823), .B1(new_n837), .B2(new_n838), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n568), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n789), .A2(new_n379), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT57), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n360), .A2(KEYINPUT57), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n784), .B(KEYINPUT120), .Z(new_n858));
  NAND2_X1  g657(.A1(new_n825), .A2(new_n543), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n629), .B1(new_n859), .B2(new_n830), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n857), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n856), .A2(new_n567), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G148gat), .B1(new_n862), .B2(new_n822), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT59), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n843), .A2(new_n851), .A3(new_n567), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1345gat));
  NAND2_X1  g666(.A1(new_n629), .A2(G155gat), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT121), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(G155gat), .B1(new_n843), .B2(new_n629), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(G1346gat));
  OAI21_X1  g671(.A(G162gat), .B1(new_n853), .B2(new_n641), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n790), .A2(new_n227), .A3(new_n809), .A4(new_n842), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1347gat));
  NAND3_X1  g674(.A1(new_n684), .A2(new_n685), .A3(new_n328), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(KEYINPUT125), .A3(new_n622), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n876), .B2(new_n621), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n785), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G169gat), .B1(new_n881), .B2(new_n606), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n791), .A2(new_n383), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT122), .B1(new_n789), .B2(new_n609), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n885), .B(new_n635), .C1(new_n783), .C2(new_n784), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(KEYINPUT123), .B(new_n883), .C1(new_n884), .C2(new_n886), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n606), .A2(G169gat), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n882), .B1(new_n894), .B2(new_n895), .ZN(G1348gat));
  INV_X1    g695(.A(G176gat), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n897), .A3(new_n568), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n891), .A2(new_n567), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n897), .ZN(G1349gat));
  OAI21_X1  g699(.A(G183gat), .B1(new_n881), .B2(new_n495), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n305), .A2(new_n306), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n629), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n901), .B1(new_n887), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g704(.A1(new_n891), .A2(new_n287), .A3(new_n749), .ZN(new_n906));
  OAI21_X1  g705(.A(G190gat), .B1(new_n881), .B2(new_n816), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(KEYINPUT126), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n908), .B2(KEYINPUT126), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n906), .B1(new_n909), .B2(new_n911), .ZN(G1351gat));
  NOR2_X1   g711(.A1(new_n876), .A2(new_n619), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n856), .A2(new_n861), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n606), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n884), .A2(new_n886), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n619), .A2(new_n360), .A3(new_n383), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n606), .A2(G197gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1352gat));
  INV_X1    g719(.A(G204gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n567), .A2(new_n921), .ZN(new_n922));
  OR3_X1    g721(.A1(new_n918), .A2(KEYINPUT62), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n913), .ZN(new_n924));
  OAI21_X1  g723(.A(G204gat), .B1(new_n862), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT62), .B1(new_n918), .B2(new_n922), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(G1353gat));
  INV_X1    g726(.A(new_n918), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n269), .A3(new_n629), .ZN(new_n929));
  INV_X1    g728(.A(new_n914), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n629), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n931), .B2(G211gat), .ZN(new_n932));
  OAI211_X1 g731(.A(KEYINPUT63), .B(G211gat), .C1(new_n914), .C2(new_n495), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n932), .B2(new_n934), .ZN(G1354gat));
  AOI21_X1  g734(.A(G218gat), .B1(new_n928), .B2(new_n749), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n543), .A2(G218gat), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT127), .Z(new_n938));
  AOI21_X1  g737(.A(new_n936), .B1(new_n930), .B2(new_n938), .ZN(G1355gat));
endmodule


