//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  OR3_X1    g0019(.A1(new_n218), .A2(new_n209), .A3(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n202), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n215), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT67), .B(G50), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT69), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G150), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n209), .A2(G33), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n254), .B1(new_n201), .B2(new_n209), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n219), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n209), .A3(G1), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n259), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n209), .A2(G1), .ZN(new_n264));
  INV_X1    g0064(.A(G50), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(new_n266), .B1(new_n265), .B2(new_n262), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n208), .A2(G274), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT70), .A2(G41), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT70), .A2(G41), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n278), .B1(G226), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n289), .A2(G223), .B1(G77), .B2(new_n287), .ZN(new_n290));
  INV_X1    g0090(.A(G222), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT3), .ZN(new_n292));
  INV_X1    g0092(.A(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n288), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n290), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n280), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n284), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n270), .B(new_n272), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n283), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT73), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n300), .B2(new_n301), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(KEYINPUT10), .B(new_n309), .C1(new_n302), .C2(new_n306), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g0113(.A(KEYINPUT8), .B(G58), .Z(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n253), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G20), .A2(G77), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT15), .B(G87), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n315), .B(new_n316), .C1(new_n256), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n259), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n263), .A2(KEYINPUT72), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT72), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n262), .B2(new_n259), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n264), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(G77), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n262), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(G77), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n296), .A2(G232), .A3(new_n288), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n296), .A2(G1698), .ZN(new_n332));
  INV_X1    g0132(.A(G238), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n331), .B1(new_n223), .B2(new_n296), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n299), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n278), .B1(G244), .B2(new_n282), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(G190), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n336), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G200), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n330), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n335), .A2(new_n341), .A3(new_n336), .ZN(new_n342));
  INV_X1    g0142(.A(G169), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n344), .C1(new_n321), .C2(new_n329), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n269), .B1(new_n304), .B2(new_n343), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(G179), .B2(new_n304), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n313), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n296), .A2(G232), .A3(G1698), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G97), .ZN(new_n353));
  INV_X1    g0153(.A(G226), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n352), .B(new_n353), .C1(new_n297), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n299), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n357));
  AOI21_X1  g0157(.A(new_n278), .B1(G238), .B2(new_n282), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT13), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n356), .A2(new_n358), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(G190), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n202), .B2(new_n256), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n259), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT11), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n325), .A2(G68), .A3(new_n326), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n261), .A2(G1), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(G20), .A3(new_n216), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT77), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g0172(.A(new_n372), .B(KEYINPUT12), .Z(new_n373));
  NAND3_X1  g0173(.A1(new_n367), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n363), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n362), .A2(new_n357), .ZN(new_n377));
  OAI21_X1  g0177(.A(G200), .B1(new_n377), .B2(new_n359), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT76), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT76), .B(G200), .C1(new_n377), .C2(new_n359), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(G169), .B1(new_n377), .B2(new_n359), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT78), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n384), .A2(new_n385), .ZN(new_n387));
  OAI211_X1 g0187(.A(G169), .B(new_n387), .C1(new_n377), .C2(new_n359), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n360), .B(G179), .C1(new_n361), .C2(new_n362), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n384), .A2(new_n385), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n382), .B1(new_n394), .B2(new_n374), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n313), .A2(new_n346), .A3(KEYINPUT74), .A4(new_n348), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n351), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n255), .A2(new_n264), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n263), .B1(new_n262), .B2(new_n255), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n259), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n294), .A2(new_n209), .A3(new_n295), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT7), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n294), .A2(new_n404), .A3(new_n209), .A4(new_n295), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(G68), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G58), .A2(G68), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT79), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(KEYINPUT79), .A2(G58), .A3(G68), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n217), .A3(new_n410), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(G20), .B1(G159), .B2(new_n253), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n401), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n406), .A2(new_n412), .A3(KEYINPUT16), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n400), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT80), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n280), .A2(G232), .A3(new_n281), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n418), .B1(new_n278), .B2(new_n419), .ZN(new_n420));
  OR2_X1    g0220(.A1(G223), .A2(G1698), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n354), .A2(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n421), .B(new_n422), .C1(new_n285), .C2(new_n286), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n299), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n280), .A2(G232), .A3(new_n281), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n274), .A2(new_n275), .A3(G45), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n427), .B(KEYINPUT80), .C1(new_n428), .C2(new_n273), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n420), .A2(new_n305), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n280), .B1(new_n423), .B2(new_n424), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n427), .B1(new_n428), .B2(new_n273), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n301), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT17), .B1(new_n417), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n413), .A2(new_n414), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(new_n416), .A3(new_n259), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n399), .A3(new_n434), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT82), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n417), .A2(KEYINPUT82), .A3(new_n434), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n435), .B1(new_n442), .B2(KEYINPUT17), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  AOI21_X1  g0244(.A(G179), .B1(new_n425), .B2(new_n299), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n420), .A3(new_n429), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n343), .B1(new_n431), .B2(new_n432), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n437), .A2(new_n399), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n444), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n417), .A2(new_n449), .A3(new_n450), .A4(KEYINPUT18), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n443), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n397), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n296), .A2(new_n209), .A3(G87), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n458), .B(KEYINPUT22), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT24), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT23), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(new_n223), .A3(G20), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n461), .B(new_n463), .C1(new_n464), .C2(new_n256), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n465), .B(KEYINPUT88), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n459), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n460), .B1(new_n459), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n259), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n208), .A2(G33), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n263), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n262), .A2(KEYINPUT25), .A3(new_n223), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT25), .B1(new_n262), .B2(new_n223), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n471), .A2(new_n223), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n296), .A2(G250), .A3(new_n288), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n296), .A2(G257), .A3(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G294), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n299), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT89), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT89), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n484), .A3(new_n299), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n208), .B(G45), .C1(new_n486), .C2(G41), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT70), .B(G41), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(new_n486), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n299), .ZN(new_n490));
  INV_X1    g0290(.A(G274), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n299), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n490), .A2(G264), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n483), .A2(new_n485), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT90), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n495), .A3(G169), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n493), .A2(new_n482), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G179), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n494), .B2(G169), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n477), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n494), .A2(G190), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n497), .A2(G200), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n469), .B(new_n476), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT21), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n296), .A2(G257), .A3(new_n288), .ZN(new_n507));
  INV_X1    g0307(.A(G303), .ZN(new_n508));
  OAI221_X1 g0308(.A(new_n507), .B1(new_n508), .B2(new_n296), .C1(new_n332), .C2(new_n224), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n299), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n492), .A2(new_n489), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n490), .A2(G270), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G169), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n464), .B1(new_n208), .B2(G33), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n322), .A2(new_n324), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G116), .B2(new_n328), .ZN(new_n517));
  AOI21_X1  g0317(.A(G20), .B1(new_n293), .B2(G97), .ZN(new_n518));
  INV_X1    g0318(.A(G283), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n293), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n464), .A2(G20), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n259), .A2(KEYINPUT86), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT86), .B1(new_n259), .B2(new_n521), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(KEYINPUT20), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n517), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n506), .B1(new_n514), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(new_n527), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(new_n516), .C1(G116), .C2(new_n328), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(KEYINPUT21), .A3(G169), .A4(new_n513), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n513), .A2(new_n341), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n531), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n529), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n513), .A2(new_n305), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n513), .A2(G200), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n528), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n536), .A2(KEYINPUT87), .A3(new_n528), .A4(new_n537), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n208), .A2(G45), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G250), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n299), .A2(new_n544), .B1(new_n491), .B2(new_n543), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  OAI221_X1 g0346(.A(new_n546), .B1(new_n297), .B2(new_n333), .C1(new_n222), .C2(new_n332), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n547), .B2(new_n299), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n301), .ZN(new_n549));
  AOI211_X1 g0349(.A(new_n305), .B(new_n545), .C1(new_n547), .C2(new_n299), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G87), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n471), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT85), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n296), .A2(new_n209), .A3(G68), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n209), .B1(new_n353), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G87), .B2(new_n206), .ZN(new_n558));
  INV_X1    g0358(.A(G97), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n556), .B1(new_n256), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n555), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n259), .B1(new_n262), .B2(new_n317), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n548), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n343), .ZN(new_n565));
  INV_X1    g0365(.A(new_n317), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n263), .A2(new_n566), .A3(new_n470), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n548), .A2(new_n341), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n551), .A2(new_n563), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT4), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n297), .A2(new_n222), .B1(KEYINPUT84), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n289), .A2(G250), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n570), .A2(KEYINPUT84), .B1(G33), .B2(G283), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NOR4_X1   g0374(.A1(new_n297), .A2(KEYINPUT84), .A3(new_n570), .A4(new_n222), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n299), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n490), .A2(G257), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n511), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n343), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n471), .A2(G97), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G97), .B2(new_n262), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT83), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT83), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n580), .B(new_n583), .C1(G97), .C2(new_n262), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT6), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n559), .A2(new_n223), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(new_n205), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n223), .A2(KEYINPUT6), .A3(G97), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n403), .A2(G107), .A3(new_n405), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n259), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n579), .B(new_n595), .C1(G179), .C2(new_n578), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n578), .A2(G200), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n582), .A2(new_n584), .B1(new_n259), .B2(new_n593), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n598), .C1(new_n305), .C2(new_n578), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n569), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n457), .A2(new_n505), .A3(new_n542), .A4(new_n600), .ZN(G372));
  INV_X1    g0401(.A(new_n348), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT92), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n453), .B2(new_n454), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n446), .A2(new_n448), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n452), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT18), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n451), .A2(new_n444), .A3(new_n452), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(KEYINPUT92), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n380), .A2(new_n381), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n375), .A3(new_n363), .ZN(new_n614));
  INV_X1    g0414(.A(new_n345), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n374), .A2(new_n394), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n443), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n612), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n602), .B1(new_n618), .B2(new_n313), .ZN(new_n619));
  INV_X1    g0419(.A(new_n457), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n569), .A2(new_n596), .A3(new_n599), .A4(new_n504), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n501), .A2(KEYINPUT91), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT91), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n477), .B(new_n623), .C1(new_n499), .C2(new_n500), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n535), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n621), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n547), .A2(new_n299), .ZN(new_n629));
  INV_X1    g0429(.A(new_n545), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n341), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n562), .A2(new_n567), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n631), .B(new_n632), .C1(G169), .C2(new_n548), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n548), .A2(G190), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n301), .B2(new_n548), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n554), .A2(new_n562), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n628), .B1(new_n596), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n598), .B1(new_n343), .B2(new_n578), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n576), .A2(new_n577), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n341), .A3(new_n511), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n569), .A2(KEYINPUT26), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n633), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n627), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n619), .B1(new_n620), .B2(new_n645), .ZN(G369));
  AND2_X1   g0446(.A1(new_n622), .A2(new_n624), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n369), .A2(new_n209), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n626), .A2(new_n653), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n505), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n542), .B1(new_n528), .B2(new_n654), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n535), .A2(new_n531), .A3(new_n653), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n477), .A2(new_n653), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n505), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n501), .A2(new_n654), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(G330), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n659), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(new_n212), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n488), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G1), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n218), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n505), .A2(new_n600), .A3(new_n542), .A4(new_n654), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT31), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n548), .A2(new_n482), .A3(new_n493), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(new_n533), .A3(new_n640), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n497), .A2(G179), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n513), .A3(new_n578), .A4(new_n564), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n654), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n678), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n682), .A3(new_n684), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n676), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  AND4_X1   g0494(.A1(new_n501), .A2(new_n532), .A3(new_n529), .A4(new_n534), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n643), .B(new_n633), .C1(new_n695), .C2(new_n621), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n694), .B1(new_n696), .B2(new_n654), .ZN(new_n697));
  INV_X1    g0497(.A(new_n621), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n647), .B2(new_n535), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n643), .A2(new_n633), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n653), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n697), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT93), .B1(new_n693), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n693), .A2(new_n702), .A3(KEYINPUT93), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n675), .B1(new_n706), .B2(G1), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT94), .ZN(G364));
  AOI21_X1  g0508(.A(new_n219), .B1(G20), .B2(new_n343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G179), .A2(G200), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G190), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n559), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n209), .A2(new_n305), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n301), .A2(G179), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n209), .A2(G190), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n716), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n717), .A2(new_n552), .B1(new_n719), .B2(new_n223), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n341), .A2(new_n301), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n718), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n296), .B1(new_n722), .B2(new_n216), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n714), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(KEYINPUT99), .B(G159), .Z(new_n725));
  NAND2_X1  g0525(.A1(new_n718), .A2(new_n710), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT101), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT100), .B(KEYINPUT32), .Z(new_n729));
  OAI21_X1  g0529(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n341), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n715), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n718), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n732), .A2(new_n215), .B1(new_n733), .B2(new_n202), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n721), .A2(new_n715), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT97), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n735), .A2(new_n736), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n734), .B1(new_n741), .B2(G50), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT98), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n730), .B(new_n743), .C1(new_n729), .C2(new_n728), .ZN(new_n744));
  INV_X1    g0544(.A(new_n717), .ZN(new_n745));
  INV_X1    g0545(.A(new_n732), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G303), .A2(new_n745), .B1(new_n746), .B2(G322), .ZN(new_n747));
  INV_X1    g0547(.A(G311), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n748), .B2(new_n733), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(G326), .B2(new_n741), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n712), .A2(G294), .ZN(new_n751));
  INV_X1    g0551(.A(new_n722), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT33), .B(G317), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n296), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n719), .ZN(new_n755));
  INV_X1    g0555(.A(new_n726), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G283), .A2(new_n755), .B1(new_n756), .B2(G329), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n750), .A2(new_n751), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT102), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n709), .B1(new_n744), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n261), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n208), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OR3_X1    g0563(.A1(new_n670), .A2(KEYINPUT95), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT95), .B1(new_n670), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n212), .A2(new_n296), .ZN(new_n768));
  INV_X1    g0568(.A(G355), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(new_n769), .B1(G116), .B2(new_n212), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n246), .A2(new_n277), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n669), .A2(new_n296), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n218), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n773), .B1(new_n277), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n770), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n709), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n767), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT96), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n760), .A2(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n785), .B1(KEYINPUT96), .B2(new_n783), .C1(new_n662), .C2(new_n780), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n662), .A2(G330), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n660), .A2(new_n676), .A3(new_n661), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n787), .A2(new_n788), .A3(new_n766), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  OR2_X1    g0591(.A1(new_n345), .A2(KEYINPUT104), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n345), .A2(KEYINPUT104), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n794), .A2(new_n340), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n654), .B(new_n795), .C1(new_n627), .C2(new_n644), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n653), .B1(new_n321), .B2(new_n329), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n792), .A2(new_n340), .A3(new_n797), .A4(new_n793), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n615), .A2(new_n653), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n796), .B1(new_n701), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n767), .B1(new_n693), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n693), .B2(new_n801), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n781), .A2(new_n778), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n767), .B1(G77), .B2(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n722), .A2(new_n519), .B1(new_n733), .B2(new_n464), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n741), .B2(G303), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT103), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G107), .A2(new_n745), .B1(new_n746), .B2(G294), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n748), .B2(new_n726), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n287), .B1(new_n719), .B2(new_n552), .ZN(new_n811));
  OR3_X1    g0611(.A1(new_n810), .A2(new_n714), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n733), .ZN(new_n813));
  INV_X1    g0613(.A(new_n725), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n813), .A2(new_n814), .B1(new_n746), .B2(G143), .ZN(new_n815));
  INV_X1    g0615(.A(G150), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(new_n722), .C1(new_n740), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n296), .B1(new_n717), .B2(new_n265), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n719), .A2(new_n216), .B1(new_n726), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n821), .B(new_n823), .C1(G58), .C2(new_n712), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT34), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n818), .B2(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n808), .A2(new_n812), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n805), .B1(new_n827), .B2(new_n709), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n800), .B2(new_n778), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n803), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G384));
  OR2_X1    g0631(.A1(new_n794), .A2(new_n653), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n796), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  INV_X1    g0635(.A(new_n651), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n452), .A2(KEYINPUT106), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT106), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n417), .B2(new_n651), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(KEYINPUT37), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n440), .A2(new_n608), .A3(new_n441), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n452), .A2(new_n836), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n440), .A2(new_n608), .A3(new_n441), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n844), .B1(new_n443), .B2(new_n455), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n835), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n843), .A2(new_n846), .ZN(new_n850));
  INV_X1    g0650(.A(new_n456), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n850), .B(KEYINPUT38), .C1(new_n851), .C2(new_n844), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n375), .A2(new_n654), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n392), .B1(new_n386), .B2(new_n388), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n614), .B(new_n855), .C1(new_n856), .C2(new_n375), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n394), .A2(new_n854), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n834), .A2(new_n853), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n612), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n651), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT107), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n604), .A2(new_n443), .A3(new_n611), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n608), .A2(KEYINPUT92), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n451), .A2(new_n603), .A3(new_n452), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n438), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT37), .B1(new_n868), .B2(new_n840), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n840), .A2(new_n865), .B1(new_n869), .B2(new_n843), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n864), .B1(new_n870), .B2(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n865), .A2(new_n840), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n843), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(KEYINPUT107), .A3(new_n835), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n871), .A2(new_n875), .A3(new_n852), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n394), .A2(new_n374), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(new_n653), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n863), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n702), .A2(new_n620), .ZN(new_n884));
  INV_X1    g0684(.A(new_n619), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n883), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n876), .A2(KEYINPUT109), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT109), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n871), .A2(new_n875), .A3(new_n889), .A4(new_n852), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n857), .A2(new_n858), .B1(new_n798), .B2(new_n799), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT108), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n687), .A2(new_n892), .A3(KEYINPUT31), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n687), .B1(new_n677), .B2(KEYINPUT31), .ZN(new_n896));
  OAI211_X1 g0696(.A(KEYINPUT40), .B(new_n891), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n888), .A2(new_n890), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n900), .B1(new_n901), .B2(new_n853), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n457), .B1(new_n896), .B2(new_n895), .ZN(new_n904));
  OAI21_X1  g0704(.A(G330), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n904), .B2(new_n903), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n887), .A2(new_n906), .B1(new_n208), .B2(new_n761), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n887), .B2(new_n906), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n774), .A2(G77), .A3(new_n409), .A4(new_n410), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n265), .A2(G68), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n208), .B(G13), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n590), .A2(KEYINPUT35), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n590), .A2(KEYINPUT35), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n219), .A2(new_n209), .A3(new_n464), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT105), .Z(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT36), .ZN(new_n917));
  OR3_X1    g0717(.A1(new_n908), .A2(new_n911), .A3(new_n917), .ZN(G367));
  NOR2_X1   g0718(.A1(new_n713), .A2(new_n216), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(G150), .B2(new_n746), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT115), .Z(new_n921));
  NAND2_X1  g0721(.A1(new_n741), .A2(G143), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n755), .A2(G77), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n215), .B2(new_n717), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n296), .B1(new_n733), .B2(new_n265), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n725), .A2(new_n722), .B1(new_n726), .B2(new_n817), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n921), .A2(new_n922), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT46), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n717), .B2(new_n464), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT114), .Z(new_n931));
  OAI21_X1  g0731(.A(new_n287), .B1(new_n732), .B2(new_n508), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n717), .A2(new_n929), .A3(new_n464), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n932), .B(new_n933), .C1(G107), .C2(new_n712), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n559), .A2(new_n719), .B1(new_n733), .B2(new_n519), .ZN(new_n935));
  INV_X1    g0735(.A(G294), .ZN(new_n936));
  INV_X1    g0736(.A(G317), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n722), .A2(new_n936), .B1(new_n726), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n934), .B(new_n939), .C1(new_n748), .C2(new_n740), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n928), .B1(new_n931), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT47), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n709), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n212), .A2(new_n317), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n782), .B(new_n944), .C1(new_n772), .C2(new_n240), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n766), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n636), .A2(new_n653), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n569), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n633), .B2(new_n947), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n943), .B(new_n946), .C1(new_n949), .C2(new_n780), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n596), .B(new_n599), .C1(new_n598), .C2(new_n654), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n639), .A2(new_n641), .A3(new_n653), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n658), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT44), .Z(new_n956));
  NAND2_X1  g0756(.A1(new_n667), .A2(KEYINPUT113), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n667), .A2(KEYINPUT113), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n659), .A2(KEYINPUT45), .A3(new_n953), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT45), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n658), .B2(new_n954), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n956), .A2(new_n957), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n957), .B1(new_n956), .B2(new_n962), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n657), .B1(new_n666), .B2(new_n656), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(new_n787), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n704), .B2(new_n705), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT112), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n706), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n670), .B(KEYINPUT41), .Z(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n763), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT110), .Z(new_n978));
  INV_X1    g0778(.A(KEYINPUT111), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n978), .A2(new_n979), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n953), .A2(new_n505), .A3(new_n656), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(KEYINPUT42), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT42), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n596), .B1(new_n951), .B2(new_n501), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n654), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n980), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n667), .A2(new_n954), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n978), .A2(new_n979), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n950), .B1(new_n976), .B2(new_n992), .ZN(G387));
  INV_X1    g0793(.A(new_n967), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n664), .A2(new_n665), .A3(new_n779), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n768), .A2(new_n672), .B1(G107), .B2(new_n212), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n237), .A2(new_n277), .ZN(new_n997));
  INV_X1    g0797(.A(new_n672), .ZN(new_n998));
  AOI211_X1 g0798(.A(G45), .B(new_n998), .C1(G68), .C2(G77), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n255), .A2(G50), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT50), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n773), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n996), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n767), .B1(new_n1003), .B2(new_n782), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n741), .A2(G159), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n732), .A2(new_n265), .B1(new_n726), .B2(new_n816), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n287), .B(new_n1006), .C1(G97), .C2(new_n755), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n566), .A2(new_n712), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n733), .A2(new_n216), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n717), .A2(new_n202), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(new_n314), .C2(new_n752), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n296), .B1(new_n756), .B2(G326), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n713), .A2(new_n519), .B1(new_n717), .B2(new_n936), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G311), .A2(new_n752), .B1(new_n813), .B2(G303), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n937), .B2(new_n732), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G322), .B2(new_n741), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1014), .B1(new_n1017), .B2(KEYINPUT48), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT48), .B2(new_n1017), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1013), .B1(new_n464), .B2(new_n719), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1012), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1004), .B1(new_n1023), .B2(new_n709), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n994), .A2(new_n763), .B1(new_n995), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n706), .A2(new_n994), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n670), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n706), .A2(new_n994), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(G393));
  NOR2_X1   g0829(.A1(new_n963), .A2(new_n964), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n1026), .B2(KEYINPUT112), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n971), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n671), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n965), .A2(new_n763), .ZN(new_n1035));
  AOI21_X1  g0835(.A(KEYINPUT116), .B1(new_n954), .B2(new_n779), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n741), .A2(G150), .B1(G159), .B2(new_n746), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT51), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G50), .A2(new_n752), .B1(new_n756), .B2(G143), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n216), .B2(new_n717), .C1(new_n255), .C2(new_n733), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n296), .B1(new_n719), .B2(new_n552), .C1(new_n713), .C2(new_n202), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n740), .A2(new_n937), .B1(new_n748), .B2(new_n732), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  AOI22_X1  g0844(.A1(G283), .A2(new_n745), .B1(new_n756), .B2(G322), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n936), .B2(new_n733), .C1(new_n508), .C2(new_n722), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n287), .B1(new_n719), .B2(new_n223), .C1(new_n713), .C2(new_n464), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n709), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n251), .A2(new_n772), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n782), .B1(G97), .B2(new_n669), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n766), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT117), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT118), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n954), .A2(KEYINPUT116), .A3(new_n779), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1035), .B1(new_n1036), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1034), .A2(new_n1058), .ZN(G390));
  OAI211_X1 g0859(.A(G330), .B(new_n891), .C1(new_n895), .C2(new_n896), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT119), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n696), .A2(new_n654), .A3(new_n795), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n832), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n880), .B1(new_n1064), .B2(new_n859), .ZN(new_n1065));
  AND3_X1   g0865(.A1(new_n888), .A2(new_n1065), .A3(new_n890), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n880), .B1(new_n833), .B2(new_n859), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n878), .B2(new_n881), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1062), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n878), .A2(new_n881), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1067), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n691), .ZN(new_n1073));
  OAI211_X1 g0873(.A(G330), .B(new_n800), .C1(new_n896), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n859), .C1(KEYINPUT119), .C2(new_n1060), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n888), .A2(new_n1065), .A3(new_n890), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1069), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1079), .A2(new_n762), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n287), .B1(new_n756), .B2(G125), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n265), .B2(new_n719), .C1(new_n822), .C2(new_n732), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n745), .A2(G150), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT53), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1082), .B(new_n1084), .C1(G128), .C2(new_n741), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT54), .B(G143), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n722), .A2(new_n817), .B1(new_n733), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G159), .B2(new_n712), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT121), .Z(new_n1089));
  OAI21_X1  g0889(.A(new_n287), .B1(new_n717), .B2(new_n552), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n719), .A2(new_n216), .B1(new_n726), .B2(new_n936), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(G77), .C2(new_n712), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G107), .A2(new_n752), .B1(new_n813), .B2(G97), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n464), .B2(new_n732), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G283), .B2(new_n741), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1085), .A2(new_n1089), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n767), .B1(new_n314), .B2(new_n804), .C1(new_n1096), .C2(new_n781), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1070), .B2(new_n777), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1080), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n457), .B(G330), .C1(new_n896), .C2(new_n895), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n619), .C1(new_n620), .C2(new_n702), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1074), .A2(new_n860), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1060), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n833), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n692), .A2(new_n800), .A3(new_n859), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1064), .ZN(new_n1106));
  OAI211_X1 g0906(.A(G330), .B(new_n800), .C1(new_n895), .C2(new_n896), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n860), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1101), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n671), .B1(new_n1079), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1069), .A2(new_n1078), .A3(new_n1110), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1112), .A2(KEYINPUT120), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT120), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1099), .B1(new_n1114), .B2(new_n1115), .ZN(G378));
  INV_X1    g0916(.A(new_n1101), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n899), .A2(G330), .A3(new_n902), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n313), .A2(new_n348), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n268), .A2(new_n836), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1119), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT123), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1124), .A2(KEYINPUT123), .A3(new_n1125), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1132), .A2(new_n899), .A3(G330), .A4(new_n902), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n883), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n883), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1118), .A2(new_n1136), .A3(KEYINPUT57), .A4(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(KEYINPUT124), .A3(new_n670), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1118), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT124), .B1(new_n1138), .B2(new_n670), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n767), .B1(G50), .B2(new_n804), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1132), .A2(new_n778), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n287), .A2(new_n276), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(new_n265), .C1(G33), .C2(G41), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT122), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n722), .A2(new_n559), .B1(new_n726), .B2(new_n519), .ZN(new_n1151));
  NOR4_X1   g0951(.A1(new_n919), .A2(new_n1151), .A3(new_n1010), .A4(new_n1148), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n732), .A2(new_n223), .B1(new_n719), .B2(new_n215), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n566), .B2(new_n813), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(new_n464), .C2(new_n740), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT58), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1150), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n741), .A2(G125), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n717), .A2(new_n1086), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n722), .A2(new_n822), .B1(new_n733), .B2(new_n817), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(G128), .C2(new_n746), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1158), .B(new_n1161), .C1(new_n816), .C2(new_n713), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n814), .A2(new_n755), .ZN(new_n1164));
  AOI211_X1 g0964(.A(G33), .B(G41), .C1(new_n756), .C2(G124), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1157), .B1(new_n1156), .B2(new_n1155), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1146), .B(new_n1147), .C1(new_n709), .C2(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n1170), .B2(new_n763), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1145), .A2(new_n1171), .ZN(G375));
  NAND2_X1  g0972(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(new_n1117), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1174), .A2(new_n974), .A3(new_n1110), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT125), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n860), .A2(new_n777), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n767), .B1(G68), .B2(new_n804), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G283), .A2(new_n746), .B1(new_n756), .B2(G303), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1179), .A2(new_n287), .A3(new_n923), .A4(new_n1008), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G97), .A2(new_n745), .B1(new_n813), .B2(G107), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n464), .B2(new_n722), .C1(new_n740), .C2(new_n936), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G159), .A2(new_n745), .B1(new_n813), .B2(G150), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n722), .B2(new_n1086), .C1(new_n740), .C2(new_n822), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G137), .A2(new_n746), .B1(new_n756), .B2(G128), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n287), .B1(new_n755), .B2(G58), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n265), .C2(new_n713), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n1180), .A2(new_n1182), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1178), .B1(new_n1188), .B2(new_n709), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1173), .A2(new_n763), .B1(new_n1177), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1176), .A2(new_n1190), .ZN(G381));
  AOI211_X1 g0991(.A(new_n1098), .B(new_n1080), .C1(new_n1113), .C2(new_n1112), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1145), .A2(new_n1171), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n950), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n706), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1031), .B2(new_n971), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n762), .B1(new_n1197), .B2(new_n974), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1195), .B1(new_n1198), .B2(new_n991), .ZN(new_n1199));
  OR2_X1    g0999(.A1(G393), .A2(G396), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1194), .A2(new_n1199), .A3(new_n1201), .ZN(G407));
  OAI211_X1 g1002(.A(G407), .B(G213), .C1(G343), .C2(new_n1193), .ZN(G409));
  OAI211_X1 g1003(.A(G378), .B(new_n1171), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1171), .B1(new_n974), .B2(new_n1140), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1192), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n652), .A2(G213), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1208), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n1111), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n670), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1174), .B1(KEYINPUT60), .B2(new_n1111), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1190), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n830), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1214), .A2(new_n830), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G2897), .B(new_n1210), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1217), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1210), .A2(G2897), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1215), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT61), .B1(new_n1209), .B2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1034), .A2(new_n1058), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G387), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1199), .A2(G390), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(G393), .B(new_n790), .ZN(new_n1228));
  AND4_X1   g1028(.A1(KEYINPUT126), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT126), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1199), .B2(G390), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1231), .A2(new_n1228), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT63), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1234), .B1(new_n1209), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1210), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(KEYINPUT63), .A3(new_n1235), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1224), .A2(new_n1233), .A3(new_n1237), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT62), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1238), .A2(new_n1241), .A3(new_n1235), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1238), .B2(new_n1222), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1241), .B1(new_n1238), .B2(new_n1235), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1242), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1240), .B1(new_n1246), .B2(new_n1233), .ZN(G405));
  OAI21_X1  g1047(.A(KEYINPUT127), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1231), .A2(new_n1228), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT127), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1226), .A2(new_n1227), .A3(KEYINPUT126), .A4(new_n1228), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G375), .A2(new_n1192), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1255), .A2(new_n1236), .A3(new_n1204), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1236), .B1(new_n1255), .B2(new_n1204), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1248), .B(new_n1254), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n1204), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1235), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1255), .A2(new_n1236), .A3(new_n1204), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(new_n1252), .A3(new_n1233), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1262), .ZN(G402));
endmodule


