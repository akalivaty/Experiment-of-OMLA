

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(n517), .A2(G2104), .ZN(n535) );
  NOR2_X1 U551 ( .A1(KEYINPUT33), .A2(n753), .ZN(n755) );
  BUF_X1 U552 ( .A(n615), .Z(n616) );
  BUF_X1 U553 ( .A(n535), .Z(n515) );
  XNOR2_X1 U554 ( .A(KEYINPUT31), .B(n700), .ZN(n739) );
  AND2_X1 U555 ( .A1(n742), .A2(G8), .ZN(n516) );
  OR2_X1 U556 ( .A1(n677), .A2(G1384), .ZN(n681) );
  INV_X1 U557 ( .A(n691), .ZN(n692) );
  NAND2_X1 U558 ( .A1(n692), .A2(G8), .ZN(n804) );
  INV_X1 U559 ( .A(KEYINPUT65), .ZN(n751) );
  OR2_X1 U560 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U561 ( .A1(G651), .A2(n635), .ZN(n642) );
  INV_X1 U562 ( .A(G2105), .ZN(n517) );
  AND2_X1 U563 ( .A1(n517), .A2(G2104), .ZN(n615) );
  NAND2_X1 U564 ( .A1(G101), .A2(n615), .ZN(n518) );
  XNOR2_X1 U565 ( .A(n518), .B(KEYINPUT23), .ZN(n519) );
  XNOR2_X1 U566 ( .A(n519), .B(KEYINPUT67), .ZN(n521) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n886) );
  NAND2_X1 U568 ( .A1(G113), .A2(n886), .ZN(n520) );
  NAND2_X1 U569 ( .A1(n521), .A2(n520), .ZN(n526) );
  NAND2_X1 U570 ( .A1(G125), .A2(n515), .ZN(n524) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n522), .Z(n883) );
  NAND2_X1 U573 ( .A1(G137), .A2(n883), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X2 U575 ( .A1(n526), .A2(n525), .ZN(G160) );
  NOR2_X1 U576 ( .A1(G651), .A2(G543), .ZN(n646) );
  NAND2_X1 U577 ( .A1(n646), .A2(G85), .ZN(n528) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  XOR2_X1 U579 ( .A(G651), .B(KEYINPUT68), .Z(n529) );
  NOR2_X1 U580 ( .A1(n635), .A2(n529), .ZN(n647) );
  NAND2_X1 U581 ( .A1(G72), .A2(n647), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n534) );
  NAND2_X1 U583 ( .A1(n642), .A2(G47), .ZN(n532) );
  NOR2_X1 U584 ( .A1(G543), .A2(n529), .ZN(n530) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n530), .Z(n586) );
  BUF_X1 U586 ( .A(n586), .Z(n643) );
  NAND2_X1 U587 ( .A1(G60), .A2(n643), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n532), .A2(n531), .ZN(n533) );
  OR2_X1 U589 ( .A1(n534), .A2(n533), .ZN(G290) );
  AND2_X1 U590 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U591 ( .A1(n883), .A2(G138), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G126), .A2(n535), .ZN(n536) );
  XNOR2_X1 U593 ( .A(n536), .B(KEYINPUT93), .ZN(n540) );
  NAND2_X1 U594 ( .A1(G102), .A2(n615), .ZN(n538) );
  NAND2_X1 U595 ( .A1(G114), .A2(n886), .ZN(n537) );
  NAND2_X1 U596 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n677) );
  AND2_X1 U598 ( .A1(n541), .A2(n677), .ZN(G164) );
  INV_X1 U599 ( .A(G57), .ZN(G237) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  NAND2_X1 U601 ( .A1(n646), .A2(G88), .ZN(n543) );
  NAND2_X1 U602 ( .A1(G75), .A2(n647), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U604 ( .A(KEYINPUT90), .B(n544), .Z(n548) );
  NAND2_X1 U605 ( .A1(n643), .A2(G62), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n642), .A2(G50), .ZN(n545) );
  AND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(G303) );
  XNOR2_X1 U609 ( .A(KEYINPUT6), .B(KEYINPUT78), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n642), .A2(G51), .ZN(n550) );
  NAND2_X1 U611 ( .A1(G63), .A2(n643), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U613 ( .A(n552), .B(n551), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n646), .A2(G89), .ZN(n553) );
  XNOR2_X1 U615 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U616 ( .A1(G76), .A2(n647), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U618 ( .A(KEYINPUT5), .B(n556), .Z(n557) );
  NOR2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U620 ( .A(KEYINPUT79), .B(KEYINPUT7), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n560), .B(n559), .ZN(G168) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(n561) );
  XNOR2_X1 U623 ( .A(KEYINPUT80), .B(n561), .ZN(G286) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n562) );
  XOR2_X1 U625 ( .A(n562), .B(KEYINPUT10), .Z(n829) );
  NAND2_X1 U626 ( .A1(n829), .A2(G567), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(KEYINPUT11), .ZN(n564) );
  XNOR2_X1 U628 ( .A(KEYINPUT73), .B(n564), .ZN(G234) );
  NAND2_X1 U629 ( .A1(n646), .A2(G81), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G68), .A2(n647), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT13), .B(KEYINPUT74), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G56), .A2(n643), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n570), .Z(n571) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n642), .A2(G43), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n983) );
  INV_X1 U640 ( .A(G860), .ZN(n606) );
  OR2_X1 U641 ( .A1(n983), .A2(n606), .ZN(G153) );
  NAND2_X1 U642 ( .A1(G77), .A2(n647), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT69), .B(n575), .Z(n577) );
  NAND2_X1 U644 ( .A1(n646), .A2(G90), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U646 ( .A(KEYINPUT9), .B(n578), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n643), .A2(G64), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n642), .A2(G52), .ZN(n579) );
  AND2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(G301) );
  INV_X1 U651 ( .A(G301), .ZN(G171) );
  INV_X1 U652 ( .A(G868), .ZN(n660) );
  NOR2_X1 U653 ( .A1(n660), .A2(G171), .ZN(n583) );
  XNOR2_X1 U654 ( .A(n583), .B(KEYINPUT75), .ZN(n595) );
  NAND2_X1 U655 ( .A1(G54), .A2(n642), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n646), .A2(G92), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G79), .A2(n647), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n586), .A2(G66), .ZN(n587) );
  XOR2_X1 U660 ( .A(KEYINPUT76), .B(n587), .Z(n588) );
  NOR2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U663 ( .A(n592), .B(KEYINPUT15), .ZN(n593) );
  XOR2_X1 U664 ( .A(KEYINPUT77), .B(n593), .Z(n986) );
  INV_X1 U665 ( .A(n986), .ZN(n903) );
  NAND2_X1 U666 ( .A1(n660), .A2(n903), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U668 ( .A1(n642), .A2(G53), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G65), .A2(n643), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n646), .A2(G91), .ZN(n599) );
  NAND2_X1 U672 ( .A1(G78), .A2(n647), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U674 ( .A(KEYINPUT70), .B(n600), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U676 ( .A(n603), .B(KEYINPUT71), .Z(n991) );
  INV_X1 U677 ( .A(n991), .ZN(G299) );
  NAND2_X1 U678 ( .A1(G868), .A2(G286), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G299), .A2(n660), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U681 ( .A1(n606), .A2(G559), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n607), .A2(n986), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n983), .ZN(n609) );
  XOR2_X1 U685 ( .A(KEYINPUT81), .B(n609), .Z(n613) );
  NAND2_X1 U686 ( .A1(n986), .A2(G868), .ZN(n610) );
  NOR2_X1 U687 ( .A1(G559), .A2(n610), .ZN(n611) );
  XNOR2_X1 U688 ( .A(KEYINPUT82), .B(n611), .ZN(n612) );
  NOR2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U690 ( .A1(n886), .A2(G111), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n614), .B(KEYINPUT84), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G99), .A2(n616), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT85), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G135), .A2(n883), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G123), .A2(n515), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n622), .B(KEYINPUT18), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT83), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n930) );
  XOR2_X1 U701 ( .A(G2096), .B(n930), .Z(n626) );
  NOR2_X1 U702 ( .A1(G2100), .A2(n626), .ZN(n627) );
  XOR2_X1 U703 ( .A(KEYINPUT86), .B(n627), .Z(G156) );
  NAND2_X1 U704 ( .A1(G86), .A2(n646), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G48), .A2(n642), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n647), .A2(G73), .ZN(n630) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n630), .Z(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G61), .A2(n643), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U712 ( .A1(n642), .A2(G49), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G87), .A2(n635), .ZN(n637) );
  NAND2_X1 U714 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U716 ( .A1(n643), .A2(n638), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U718 ( .A(KEYINPUT89), .B(n641), .Z(G288) );
  XNOR2_X1 U719 ( .A(KEYINPUT19), .B(G288), .ZN(n653) );
  NAND2_X1 U720 ( .A1(n642), .A2(G55), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G67), .A2(n643), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n646), .A2(G93), .ZN(n649) );
  NAND2_X1 U724 ( .A1(G80), .A2(n647), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U727 ( .A(n652), .B(KEYINPUT88), .Z(n836) );
  XOR2_X1 U728 ( .A(n653), .B(n836), .Z(n654) );
  XOR2_X1 U729 ( .A(G303), .B(n654), .Z(n656) );
  XOR2_X1 U730 ( .A(n983), .B(G299), .Z(n655) );
  XNOR2_X1 U731 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U732 ( .A(n657), .B(G290), .Z(n658) );
  XNOR2_X1 U733 ( .A(G305), .B(n658), .ZN(n904) );
  NAND2_X1 U734 ( .A1(n986), .A2(G559), .ZN(n834) );
  XOR2_X1 U735 ( .A(n904), .B(n834), .Z(n659) );
  NOR2_X1 U736 ( .A1(n660), .A2(n659), .ZN(n662) );
  NOR2_X1 U737 ( .A1(G868), .A2(n836), .ZN(n661) );
  NOR2_X1 U738 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XOR2_X1 U744 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U746 ( .A1(G219), .A2(G220), .ZN(n668) );
  XNOR2_X1 U747 ( .A(KEYINPUT22), .B(KEYINPUT91), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U749 ( .A1(n669), .A2(G218), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G96), .A2(n670), .ZN(n839) );
  NAND2_X1 U751 ( .A1(n839), .A2(G2106), .ZN(n675) );
  NAND2_X1 U752 ( .A1(G108), .A2(G120), .ZN(n671) );
  NOR2_X1 U753 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n672), .A2(G69), .ZN(n673) );
  XNOR2_X1 U755 ( .A(n673), .B(KEYINPUT92), .ZN(n838) );
  NAND2_X1 U756 ( .A1(n838), .A2(G567), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n675), .A2(n674), .ZN(n841) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U759 ( .A1(n841), .A2(n676), .ZN(n832) );
  NAND2_X1 U760 ( .A1(n832), .A2(G36), .ZN(G176) );
  INV_X1 U761 ( .A(G303), .ZN(G166) );
  INV_X1 U762 ( .A(G1384), .ZN(n678) );
  AND2_X1 U763 ( .A1(G138), .A2(n678), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n883), .A2(n679), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n681), .A2(n680), .ZN(n683) );
  INV_X1 U766 ( .A(KEYINPUT66), .ZN(n682) );
  XNOR2_X1 U767 ( .A(n683), .B(n682), .ZN(n776) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n777) );
  NOR2_X1 U769 ( .A1(n776), .A2(n777), .ZN(n684) );
  XNOR2_X1 U770 ( .A(n684), .B(KEYINPUT64), .ZN(n691) );
  NOR2_X1 U771 ( .A1(n692), .A2(G2084), .ZN(n685) );
  NAND2_X1 U772 ( .A1(G8), .A2(n685), .ZN(n731) );
  NOR2_X1 U773 ( .A1(G1966), .A2(n804), .ZN(n729) );
  INV_X1 U774 ( .A(n685), .ZN(n686) );
  NAND2_X1 U775 ( .A1(G8), .A2(n686), .ZN(n687) );
  OR2_X1 U776 ( .A1(n729), .A2(n687), .ZN(n688) );
  XNOR2_X1 U777 ( .A(n688), .B(KEYINPUT30), .ZN(n689) );
  XOR2_X1 U778 ( .A(KEYINPUT99), .B(n689), .Z(n690) );
  NOR2_X1 U779 ( .A1(G168), .A2(n690), .ZN(n697) );
  XNOR2_X1 U780 ( .A(G2078), .B(KEYINPUT25), .ZN(n965) );
  NAND2_X1 U781 ( .A1(n693), .A2(n965), .ZN(n695) );
  INV_X1 U782 ( .A(n692), .ZN(n693) );
  INV_X1 U783 ( .A(n693), .ZN(n733) );
  XOR2_X1 U784 ( .A(G1961), .B(KEYINPUT96), .Z(n1004) );
  NAND2_X1 U785 ( .A1(n733), .A2(n1004), .ZN(n694) );
  NAND2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n701) );
  NOR2_X1 U787 ( .A1(G171), .A2(n701), .ZN(n696) );
  NOR2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U789 ( .A(n698), .B(KEYINPUT100), .ZN(n699) );
  INV_X1 U790 ( .A(n699), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n701), .A2(G171), .ZN(n727) );
  NAND2_X1 U792 ( .A1(G1956), .A2(n733), .ZN(n704) );
  NAND2_X1 U793 ( .A1(G2072), .A2(n693), .ZN(n702) );
  XOR2_X1 U794 ( .A(KEYINPUT27), .B(n702), .Z(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U796 ( .A(n705), .B(KEYINPUT97), .ZN(n719) );
  NOR2_X1 U797 ( .A1(n991), .A2(n719), .ZN(n706) );
  XOR2_X1 U798 ( .A(n706), .B(KEYINPUT28), .Z(n723) );
  NAND2_X1 U799 ( .A1(n693), .A2(G1996), .ZN(n707) );
  XNOR2_X1 U800 ( .A(n707), .B(KEYINPUT26), .ZN(n709) );
  NAND2_X1 U801 ( .A1(n733), .A2(G1341), .ZN(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U803 ( .A1(n983), .A2(n710), .ZN(n715) );
  NAND2_X1 U804 ( .A1(G2067), .A2(n693), .ZN(n712) );
  NAND2_X1 U805 ( .A1(n733), .A2(G1348), .ZN(n711) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n716) );
  INV_X1 U807 ( .A(n716), .ZN(n713) );
  AND2_X1 U808 ( .A1(n986), .A2(n713), .ZN(n714) );
  OR2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n903), .A2(n716), .ZN(n717) );
  NAND2_X1 U811 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n991), .A2(n719), .ZN(n720) );
  NAND2_X1 U813 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n725) );
  XOR2_X1 U815 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n724) );
  XNOR2_X1 U816 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n737) );
  AND2_X1 U818 ( .A1(n739), .A2(n737), .ZN(n728) );
  NOR2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n796) );
  NAND2_X1 U821 ( .A1(G1976), .A2(G288), .ZN(n980) );
  AND2_X1 U822 ( .A1(n796), .A2(n980), .ZN(n745) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n804), .ZN(n732) );
  XNOR2_X1 U824 ( .A(KEYINPUT101), .B(n732), .ZN(n736) );
  NOR2_X1 U825 ( .A1(n733), .A2(G2090), .ZN(n734) );
  NOR2_X1 U826 ( .A1(G166), .A2(n734), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n740) );
  AND2_X1 U828 ( .A1(n737), .A2(n740), .ZN(n738) );
  NAND2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n743) );
  INV_X1 U830 ( .A(n740), .ZN(n741) );
  OR2_X1 U831 ( .A1(n741), .A2(G286), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n743), .A2(n516), .ZN(n744) );
  XNOR2_X1 U833 ( .A(n744), .B(KEYINPUT32), .ZN(n797) );
  NAND2_X1 U834 ( .A1(n745), .A2(n797), .ZN(n749) );
  INV_X1 U835 ( .A(n980), .ZN(n747) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n746) );
  NOR2_X1 U838 ( .A1(n756), .A2(n746), .ZN(n990) );
  OR2_X1 U839 ( .A1(n747), .A2(n990), .ZN(n748) );
  AND2_X1 U840 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n804), .A2(n750), .ZN(n752) );
  XNOR2_X1 U842 ( .A(n752), .B(n751), .ZN(n753) );
  INV_X1 U843 ( .A(KEYINPUT102), .ZN(n754) );
  XNOR2_X1 U844 ( .A(n755), .B(n754), .ZN(n793) );
  NAND2_X1 U845 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n804), .A2(n757), .ZN(n759) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n994) );
  INV_X1 U848 ( .A(n994), .ZN(n758) );
  NOR2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n790) );
  NAND2_X1 U850 ( .A1(G95), .A2(n616), .ZN(n761) );
  NAND2_X1 U851 ( .A1(G107), .A2(n886), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U853 ( .A1(G131), .A2(n883), .ZN(n762) );
  XNOR2_X1 U854 ( .A(KEYINPUT95), .B(n762), .ZN(n763) );
  NOR2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n515), .A2(G119), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n880) );
  AND2_X1 U858 ( .A1(n880), .A2(G1991), .ZN(n775) );
  NAND2_X1 U859 ( .A1(G141), .A2(n883), .ZN(n768) );
  NAND2_X1 U860 ( .A1(G117), .A2(n886), .ZN(n767) );
  NAND2_X1 U861 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n616), .A2(G105), .ZN(n769) );
  XOR2_X1 U863 ( .A(KEYINPUT38), .B(n769), .Z(n770) );
  NOR2_X1 U864 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U865 ( .A1(n515), .A2(G129), .ZN(n772) );
  NAND2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n893) );
  AND2_X1 U867 ( .A1(n893), .A2(G1996), .ZN(n774) );
  NOR2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n933) );
  INV_X1 U869 ( .A(n933), .ZN(n779) );
  INV_X1 U870 ( .A(n776), .ZN(n778) );
  NOR2_X1 U871 ( .A1(n778), .A2(n777), .ZN(n822) );
  NAND2_X1 U872 ( .A1(n779), .A2(n822), .ZN(n811) );
  NAND2_X1 U873 ( .A1(G104), .A2(n616), .ZN(n781) );
  NAND2_X1 U874 ( .A1(G140), .A2(n883), .ZN(n780) );
  NAND2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n782), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n515), .A2(G128), .ZN(n783) );
  XNOR2_X1 U878 ( .A(n783), .B(KEYINPUT94), .ZN(n785) );
  NAND2_X1 U879 ( .A1(G116), .A2(n886), .ZN(n784) );
  NAND2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U881 ( .A(KEYINPUT35), .B(n786), .Z(n787) );
  NOR2_X1 U882 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U883 ( .A(KEYINPUT36), .B(n789), .ZN(n900) );
  XNOR2_X1 U884 ( .A(KEYINPUT37), .B(G2067), .ZN(n820) );
  NOR2_X1 U885 ( .A1(n900), .A2(n820), .ZN(n940) );
  NAND2_X1 U886 ( .A1(n822), .A2(n940), .ZN(n818) );
  AND2_X1 U887 ( .A1(n811), .A2(n818), .ZN(n795) );
  AND2_X1 U888 ( .A1(n790), .A2(n795), .ZN(n791) );
  XNOR2_X1 U889 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U890 ( .A1(n982), .A2(n822), .ZN(n794) );
  AND2_X1 U891 ( .A1(n791), .A2(n794), .ZN(n792) );
  NAND2_X1 U892 ( .A1(n793), .A2(n792), .ZN(n827) );
  INV_X1 U893 ( .A(n794), .ZN(n810) );
  INV_X1 U894 ( .A(n795), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n796), .A2(n797), .ZN(n800) );
  NOR2_X1 U896 ( .A1(G2090), .A2(G303), .ZN(n798) );
  NAND2_X1 U897 ( .A1(G8), .A2(n798), .ZN(n799) );
  NAND2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n801) );
  AND2_X1 U899 ( .A1(n801), .A2(n804), .ZN(n806) );
  NOR2_X1 U900 ( .A1(G1981), .A2(G305), .ZN(n802) );
  XOR2_X1 U901 ( .A(n802), .B(KEYINPUT24), .Z(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n825) );
  XOR2_X1 U905 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n817) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n893), .ZN(n927) );
  INV_X1 U907 ( .A(n811), .ZN(n814) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n880), .ZN(n931) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U910 ( .A1(n931), .A2(n812), .ZN(n813) );
  NOR2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n927), .A2(n815), .ZN(n816) );
  XNOR2_X1 U913 ( .A(n817), .B(n816), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n900), .A2(n820), .ZN(n941) );
  NAND2_X1 U916 ( .A1(n821), .A2(n941), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  AND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U920 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n829), .ZN(G217) );
  INV_X1 U922 ( .A(n829), .ZN(G223) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U924 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  XOR2_X1 U929 ( .A(KEYINPUT87), .B(n983), .Z(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n835) );
  NOR2_X1 U931 ( .A1(G860), .A2(n835), .ZN(n837) );
  XOR2_X1 U932 ( .A(n837), .B(n836), .Z(G145) );
  INV_X1 U933 ( .A(G108), .ZN(G238) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  NOR2_X1 U935 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U936 ( .A(n840), .B(KEYINPUT108), .Z(G261) );
  INV_X1 U937 ( .A(G261), .ZN(G325) );
  INV_X1 U938 ( .A(n841), .ZN(G319) );
  XOR2_X1 U939 ( .A(G1976), .B(G1971), .Z(n843) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n853) );
  XOR2_X1 U942 ( .A(KEYINPUT41), .B(G2474), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1956), .B(KEYINPUT109), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U945 ( .A(G1981), .B(G1961), .Z(n847) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1966), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U949 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n853), .B(n852), .Z(G229) );
  XOR2_X1 U952 ( .A(G2100), .B(G2096), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U955 ( .A(KEYINPUT43), .B(G2090), .Z(n857) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U959 ( .A(G2084), .B(G2078), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(G227) );
  NAND2_X1 U961 ( .A1(G100), .A2(n616), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G112), .A2(n886), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U964 ( .A(KEYINPUT114), .B(n864), .ZN(n871) );
  NAND2_X1 U965 ( .A1(n515), .A2(G124), .ZN(n865) );
  XOR2_X1 U966 ( .A(KEYINPUT44), .B(n865), .Z(n868) );
  NAND2_X1 U967 ( .A1(n883), .A2(G136), .ZN(n866) );
  XOR2_X1 U968 ( .A(KEYINPUT112), .B(n866), .Z(n867) );
  NOR2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n869), .B(KEYINPUT113), .ZN(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(G162) );
  NAND2_X1 U972 ( .A1(G130), .A2(n515), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G118), .A2(n886), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G106), .A2(n616), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G142), .A2(n883), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U978 ( .A(KEYINPUT45), .B(n876), .Z(n877) );
  NOR2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n930), .B(n879), .ZN(n899) );
  XOR2_X1 U981 ( .A(n880), .B(G162), .Z(n897) );
  XOR2_X1 U982 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n882) );
  XNOR2_X1 U983 ( .A(G164), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n882), .B(n881), .ZN(n892) );
  NAND2_X1 U985 ( .A1(G103), .A2(n616), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G139), .A2(n883), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G127), .A2(n515), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G115), .A2(n886), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n945) );
  XOR2_X1 U993 ( .A(n892), .B(n945), .Z(n895) );
  XOR2_X1 U994 ( .A(G160), .B(n893), .Z(n894) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U998 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U1000 ( .A(n903), .B(G286), .Z(n905) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1002 ( .A(n906), .B(G301), .Z(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G397) );
  XOR2_X1 U1004 ( .A(G2438), .B(G2435), .Z(n909) );
  XNOR2_X1 U1005 ( .A(G2430), .B(G2454), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n913) );
  XOR2_X1 U1007 ( .A(G2446), .B(KEYINPUT105), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G2451), .B(G2427), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1010 ( .A(n913), .B(n912), .Z(n915) );
  XNOR2_X1 U1011 ( .A(KEYINPUT104), .B(G2443), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n918) );
  XOR2_X1 U1013 ( .A(G1341), .B(G1348), .Z(n916) );
  XNOR2_X1 U1014 ( .A(KEYINPUT106), .B(n916), .ZN(n917) );
  XOR2_X1 U1015 ( .A(n918), .B(n917), .Z(n919) );
  NAND2_X1 U1016 ( .A1(G14), .A2(n919), .ZN(n925) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n925), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  INV_X1 U1025 ( .A(n925), .ZN(G401) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(KEYINPUT117), .B(n928), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(n929), .B(KEYINPUT51), .ZN(n938) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n936) );
  XOR2_X1 U1032 ( .A(G2084), .B(G160), .Z(n934) );
  XNOR2_X1 U1033 ( .A(KEYINPUT116), .B(n934), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(KEYINPUT118), .B(n943), .ZN(n952) );
  XNOR2_X1 U1039 ( .A(G164), .B(G2078), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n944), .B(KEYINPUT120), .ZN(n948) );
  XOR2_X1 U1041 ( .A(G2072), .B(n945), .Z(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT119), .B(n946), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1044 ( .A(KEYINPUT121), .B(n949), .Z(n950) );
  XNOR2_X1 U1045 ( .A(KEYINPUT50), .B(n950), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n953), .ZN(n954) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n975) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n975), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(G29), .ZN(n1034) );
  XNOR2_X1 U1051 ( .A(G2084), .B(G34), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n956), .B(KEYINPUT54), .ZN(n973) );
  XNOR2_X1 U1053 ( .A(G2090), .B(G35), .ZN(n970) );
  XNOR2_X1 U1054 ( .A(G2067), .B(G26), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(G33), .B(G2072), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n964) );
  XOR2_X1 U1057 ( .A(G32), .B(G1996), .Z(n959) );
  NAND2_X1 U1058 ( .A1(n959), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(G25), .B(G1991), .ZN(n960) );
  XNOR2_X1 U1060 ( .A(KEYINPUT122), .B(n960), .ZN(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1063 ( .A(G27), .B(n965), .Z(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n968), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(n971), .B(KEYINPUT123), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n975), .B(n974), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(G29), .A2(n976), .ZN(n977) );
  XOR2_X1 U1071 ( .A(KEYINPUT124), .B(n977), .Z(n978) );
  NAND2_X1 U1072 ( .A1(G11), .A2(n978), .ZN(n1032) );
  INV_X1 U1073 ( .A(G16), .ZN(n1028) );
  XOR2_X1 U1074 ( .A(n1028), .B(KEYINPUT56), .Z(n1003) );
  NAND2_X1 U1075 ( .A1(G1971), .A2(G303), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1078 ( .A(G1341), .B(n983), .Z(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1080 ( .A(G1348), .B(n986), .Z(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1083 ( .A(G1956), .B(n991), .Z(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n1001) );
  XOR2_X1 U1085 ( .A(G171), .B(G1961), .Z(n999) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G168), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(n996), .B(KEYINPUT125), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT57), .B(n997), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1030) );
  XNOR2_X1 U1093 ( .A(G5), .B(n1004), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(KEYINPUT126), .ZN(n1018) );
  XNOR2_X1 U1095 ( .A(G1348), .B(KEYINPUT59), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(G4), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(G1956), .B(G20), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(KEYINPUT127), .B(G1981), .Z(n1011) );
  XNOR2_X1 U1102 ( .A(G6), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1014), .Z(n1016) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G21), .ZN(n1015) );
  NOR2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(G1971), .B(G22), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(G23), .B(G1976), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XOR2_X1 U1111 ( .A(G1986), .B(G24), .Z(n1021) );
  NAND2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1113 ( .A(KEYINPUT58), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1035), .ZN(G150) );
  INV_X1 U1121 ( .A(G150), .ZN(G311) );
endmodule

