//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1275,
    new_n1276;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n465), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n476), .B1(new_n467), .B2(G2104), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n474), .A2(G137), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n465), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n472), .A2(new_n478), .A3(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n477), .A2(new_n473), .A3(new_n475), .A4(new_n468), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT67), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n474), .A2(G2105), .A3(new_n477), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n484), .B(new_n488), .C1(G124), .C2(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n477), .A2(new_n473), .A3(new_n493), .A4(new_n468), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT3), .B(G2104), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n477), .A2(new_n473), .A3(new_n468), .A4(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n497), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(new_n509), .B1(new_n506), .B2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(G88), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(G50), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n513), .A2(new_n517), .ZN(G166));
  XOR2_X1   g093(.A(KEYINPUT69), .B(KEYINPUT7), .Z(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n510), .A2(G89), .A3(new_n514), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n521), .A2(new_n522), .A3(new_n525), .A4(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND2_X1  g103(.A1(new_n510), .A2(new_n514), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n523), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n510), .A2(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n504), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  AND2_X1   g111(.A1(new_n510), .A2(new_n514), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n537), .A2(G81), .B1(G43), .B2(new_n524), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(KEYINPUT70), .B1(new_n539), .B2(new_n504), .ZN(new_n540));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n507), .A2(new_n509), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n506), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n546), .A2(new_n547), .A3(G651), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n538), .A2(new_n540), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n540), .A2(new_n538), .A3(new_n548), .A4(KEYINPUT71), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n523), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n514), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  AOI22_X1  g138(.A1(G91), .A2(new_n537), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n542), .A2(G65), .A3(new_n543), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(KEYINPUT72), .B1(new_n567), .B2(G651), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n569));
  AOI211_X1 g144(.A(new_n569), .B(new_n504), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n564), .B1(new_n568), .B2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G166), .ZN(G303));
  OAI21_X1  g148(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n510), .A2(G87), .A3(new_n514), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n514), .A2(G49), .A3(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT73), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n574), .A2(new_n575), .A3(new_n579), .A4(new_n576), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(G288));
  NAND3_X1  g156(.A1(new_n510), .A2(G86), .A3(new_n514), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n510), .A2(KEYINPUT74), .A3(G86), .A4(new_n514), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n544), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n504), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n529), .A2(new_n594), .B1(new_n595), .B2(new_n523), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n544), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G54), .B2(new_n524), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n529), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n510), .A2(KEYINPUT10), .A3(G92), .A4(new_n514), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n599), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n599), .B1(new_n610), .B2(G868), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT75), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n610), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n610), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n554), .B2(G868), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n495), .A2(new_n479), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n483), .A2(G135), .ZN(new_n630));
  INV_X1    g205(.A(G123), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n632));
  NOR3_X1   g207(.A1(new_n632), .A2(new_n475), .A3(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n475), .B2(G111), .ZN(new_n634));
  OR2_X1    g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(G2104), .A3(new_n635), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n630), .B1(new_n489), .B2(new_n631), .C1(new_n633), .C2(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n629), .A2(new_n638), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT79), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT80), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n651), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT81), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n652), .B2(new_n655), .ZN(new_n658));
  INV_X1    g233(.A(G14), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT82), .Z(new_n665));
  NOR2_X1   g240(.A1(G2072), .A2(G2078), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n444), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n663), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(KEYINPUT17), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n663), .B(new_n664), .C1(new_n444), .C2(new_n666), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n665), .A3(new_n663), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT83), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n679), .A2(new_n681), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(new_n684), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n684), .A3(new_n682), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n693), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n677), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(new_n677), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n698), .A2(new_n699), .A3(new_n694), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n697), .A2(new_n700), .A3(new_n702), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(KEYINPUT84), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(KEYINPUT84), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G35), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT100), .Z(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G2090), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT101), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G20), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT23), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n615), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT102), .B(G1956), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT103), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n715), .A2(G2090), .ZN(new_n727));
  INV_X1    g302(.A(new_n711), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(G27), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G164), .B2(new_n728), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT99), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(new_n443), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n443), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n719), .A2(G4), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n610), .B2(new_n719), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT93), .B(G1348), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n727), .A2(new_n732), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n719), .A2(G5), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G171), .B2(new_n719), .ZN(new_n740));
  INV_X1    g315(.A(G1961), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G28), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(KEYINPUT30), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n743), .B2(KEYINPUT30), .ZN(new_n746));
  OR2_X1    g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  NAND2_X1  g322(.A1(KEYINPUT31), .A2(G11), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n745), .A2(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n637), .B2(new_n711), .ZN(new_n750));
  NAND2_X1  g325(.A1(G286), .A2(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n719), .A2(G21), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n750), .B1(new_n753), .B2(G1966), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n742), .B(new_n754), .C1(G1966), .C2(new_n753), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n708), .A2(G32), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n759), .A2(new_n760), .B1(G105), .B2(new_n479), .ZN(new_n761));
  INV_X1    g336(.A(G129), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n489), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n483), .A2(G141), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n756), .B1(new_n765), .B2(new_n708), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n768), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT24), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(G34), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(G34), .ZN(new_n773));
  AND3_X1   g348(.A1(new_n711), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G160), .B2(G29), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G2084), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(G2084), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n769), .A2(new_n770), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n755), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n495), .A2(G127), .ZN(new_n780));
  INV_X1    g355(.A(G115), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n465), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n475), .B1(new_n782), .B2(KEYINPUT98), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(KEYINPUT98), .B2(new_n782), .ZN(new_n784));
  INV_X1    g359(.A(G139), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n482), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT97), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n788));
  NAND3_X1  g363(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n784), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G29), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G29), .B2(G33), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(new_n442), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n442), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n711), .A2(G26), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT28), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n483), .A2(G140), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n799));
  INV_X1    g374(.A(G116), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G2105), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT95), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n798), .B(new_n802), .C1(G128), .C2(new_n490), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n708), .ZN(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n794), .A2(new_n795), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n738), .A2(new_n779), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT103), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n718), .A2(new_n809), .A3(new_n724), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n719), .A2(G19), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n554), .B2(new_n719), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT94), .B(G1341), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n726), .A2(new_n808), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n574), .A2(new_n575), .A3(G16), .A4(new_n576), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT88), .ZN(new_n817));
  NOR2_X1   g392(.A1(G16), .A2(G23), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT87), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n817), .B1(new_n816), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT33), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n816), .A2(new_n819), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT88), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n822), .A2(new_n827), .A3(G1976), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT32), .B(G1981), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n719), .A2(G6), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n584), .A2(new_n585), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n524), .A2(G48), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n504), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n830), .B(new_n831), .C1(new_n836), .C2(new_n719), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n831), .B1(new_n836), .B2(new_n719), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n829), .ZN(new_n839));
  OAI21_X1  g414(.A(G16), .B1(new_n513), .B2(new_n517), .ZN(new_n840));
  INV_X1    g415(.A(G1971), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n719), .A2(G22), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT89), .Z(new_n843));
  AND3_X1   g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n841), .B1(new_n840), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n828), .A2(new_n837), .A3(new_n839), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(G1976), .B1(new_n822), .B2(new_n827), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT90), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n839), .A2(new_n846), .A3(new_n837), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT90), .ZN(new_n851));
  INV_X1    g426(.A(new_n848), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n828), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n849), .A2(new_n853), .A3(KEYINPUT34), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT36), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT91), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n849), .A2(new_n853), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT34), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n711), .A2(G25), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n483), .A2(G131), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT85), .ZN(new_n865));
  OR2_X1    g440(.A1(G95), .A2(G2105), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n866), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT86), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G119), .B2(new_n490), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n863), .B1(new_n870), .B2(new_n728), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G1991), .Z(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n719), .A2(G24), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n597), .B2(new_n719), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(G1986), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(G1986), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n873), .A2(new_n874), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n859), .B1(new_n862), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT34), .B1(new_n849), .B2(new_n853), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n882), .A2(KEYINPUT91), .A3(new_n879), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n858), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n855), .A2(KEYINPUT36), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n862), .A2(new_n859), .A3(new_n880), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT91), .B1(new_n882), .B2(new_n879), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n858), .A3(new_n885), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n815), .B1(new_n887), .B2(new_n891), .ZN(G311));
  NAND2_X1  g467(.A1(new_n808), .A2(new_n814), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n809), .B1(new_n718), .B2(new_n724), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n885), .B1(new_n890), .B2(new_n858), .ZN(new_n896));
  AOI211_X1 g471(.A(new_n857), .B(new_n886), .C1(new_n888), .C2(new_n889), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n810), .B(new_n895), .C1(new_n896), .C2(new_n897), .ZN(G150));
  AOI22_X1  g473(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(new_n504), .ZN(new_n900));
  INV_X1    g475(.A(G93), .ZN(new_n901));
  INV_X1    g476(.A(G55), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n529), .A2(new_n901), .B1(new_n902), .B2(new_n523), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n904), .B1(new_n551), .B2(new_n552), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(new_n549), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n610), .A2(G559), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n911), .A2(KEYINPUT39), .ZN(new_n912));
  INV_X1    g487(.A(G860), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(KEYINPUT39), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n904), .A2(new_n913), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(G145));
  NAND2_X1  g494(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n495), .A2(new_n496), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n499), .A2(new_n501), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n499), .B2(new_n501), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n803), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n490), .A2(G130), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n475), .A2(G118), .ZN(new_n930));
  OAI21_X1  g505(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n483), .A2(KEYINPUT107), .A3(G142), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT107), .B1(new_n483), .B2(G142), .ZN(new_n933));
  OAI221_X1 g508(.A(new_n929), .B1(new_n930), .B2(new_n931), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n928), .B(new_n934), .Z(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n791), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(new_n765), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n870), .B(new_n626), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n765), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n937), .B(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n939), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n935), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n943), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n939), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n928), .B(new_n934), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n637), .B(G160), .Z(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(G162), .Z(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  INV_X1    g529(.A(new_n952), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n945), .A2(new_n955), .A3(new_n949), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g533(.A(KEYINPUT41), .ZN(new_n959));
  NOR2_X1   g534(.A1(G299), .A2(new_n609), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n569), .B1(new_n961), .B2(new_n504), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n567), .A2(KEYINPUT72), .A3(G651), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n964), .A2(new_n564), .B1(new_n608), .B2(new_n603), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n959), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G299), .A2(new_n609), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n964), .A2(new_n564), .A3(new_n608), .A4(new_n603), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(KEYINPUT41), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n618), .B(new_n610), .C1(new_n905), .C2(new_n907), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n908), .A2(new_n620), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n960), .A2(new_n965), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n972), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n975), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n980));
  INV_X1    g555(.A(new_n577), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n597), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n597), .A2(new_n981), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n984), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(KEYINPUT108), .A3(new_n982), .ZN(new_n987));
  NAND2_X1  g562(.A1(G305), .A2(G303), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n836), .A2(G166), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n985), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n991), .A2(KEYINPUT108), .A3(new_n986), .A4(new_n982), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n978), .A2(new_n977), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT42), .B1(new_n994), .B2(new_n974), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n979), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n993), .B1(new_n979), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g572(.A(G868), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(G868), .B2(new_n904), .ZN(G295));
  OAI21_X1  g574(.A(new_n998), .B1(G868), .B2(new_n904), .ZN(G331));
  NAND2_X1  g575(.A1(new_n553), .A2(new_n906), .ZN(new_n1001));
  INV_X1    g576(.A(new_n532), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n533), .A2(new_n534), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G651), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT110), .B1(new_n532), .B2(new_n535), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(G286), .ZN(new_n1008));
  NAND3_X1  g583(.A1(G168), .A2(G171), .A3(new_n1005), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n907), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1001), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n905), .B2(new_n907), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1012), .A2(new_n977), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n970), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n993), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1010), .B1(new_n1001), .B2(new_n1011), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n905), .A2(new_n1013), .A3(new_n907), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n971), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n990), .A2(new_n992), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1012), .A2(new_n977), .A3(new_n1014), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1017), .A2(new_n1023), .A3(new_n954), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT43), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1017), .A2(new_n1023), .A3(new_n1026), .A4(new_n954), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT44), .B1(new_n1028), .B2(KEYINPUT109), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1030), .B(new_n1031), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1029), .A2(new_n1032), .ZN(G397));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n1034));
  INV_X1    g609(.A(G1966), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G1384), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n497), .B2(new_n502), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n495), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n475), .ZN(new_n1042));
  INV_X1    g617(.A(G137), .ZN(new_n1043));
  OAI211_X1 g618(.A(G40), .B(new_n480), .C1(new_n482), .C2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT116), .B(new_n1037), .C1(new_n497), .C2(new_n502), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1384), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT45), .B1(new_n926), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1035), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n472), .A2(new_n478), .A3(G40), .A4(new_n480), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n497), .B2(new_n502), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n926), .A2(new_n1054), .A3(new_n1048), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1050), .A2(G168), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n1059));
  AND2_X1   g634(.A1(KEYINPUT120), .A2(G8), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1050), .A2(new_n1057), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(G8), .A3(G286), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1059), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1034), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(KEYINPUT121), .A3(new_n1063), .A4(new_n1061), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1066), .A2(new_n1072), .A3(new_n1069), .ZN(new_n1073));
  INV_X1    g648(.A(G1976), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n578), .A2(new_n1074), .A3(new_n580), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1075), .A2(KEYINPUT114), .A3(new_n1076), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n926), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n577), .A2(new_n1074), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1079), .A2(new_n1080), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT49), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n832), .A2(new_n835), .A3(G1981), .ZN(new_n1087));
  INV_X1    g662(.A(G1981), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n590), .B2(new_n582), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n582), .ZN(new_n1091));
  OAI21_X1  g666(.A(G1981), .B1(new_n835), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1092), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1090), .A2(new_n1093), .A3(G8), .A4(new_n1081), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT52), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1085), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G8), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G166), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT55), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1051), .B1(new_n1052), .B2(new_n1036), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n926), .A2(new_n1037), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n841), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n926), .A2(new_n1048), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT50), .ZN(new_n1107));
  INV_X1    g682(.A(G2090), .ZN(new_n1108));
  INV_X1    g683(.A(new_n502), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1384), .B1(new_n922), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1051), .B1(new_n1110), .B2(new_n1054), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1105), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1100), .B(new_n1101), .C1(new_n1113), .C2(new_n1097), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1097), .B1(new_n1105), .B2(new_n1112), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT115), .B1(new_n1115), .B2(new_n1099), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1105), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(G2090), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1099), .B(G8), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1096), .A2(new_n1114), .A3(new_n1116), .A4(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1102), .A2(new_n443), .A3(new_n1103), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1122), .A2(new_n1123), .B1(new_n1118), .B2(new_n741), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(G2078), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OR3_X1    g701(.A1(new_n1047), .A2(new_n1049), .A3(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1121), .A2(G301), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1071), .A2(new_n1073), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1956), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1054), .B1(new_n926), .B2(new_n1048), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1045), .B1(new_n1052), .B2(KEYINPUT50), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1102), .A2(new_n1103), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT57), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n964), .A2(new_n1138), .A3(new_n564), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1134), .A2(new_n1136), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1134), .A2(new_n1137), .A3(new_n1139), .A4(new_n1136), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(new_n609), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1118), .A2(new_n736), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1081), .A2(G2067), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT117), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n736), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1149), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1140), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT60), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1144), .A2(new_n1146), .A3(KEYINPUT117), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1150), .B1(new_n1149), .B2(new_n1145), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1154), .A2(new_n610), .A3(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT60), .B(new_n609), .C1(new_n1147), .C2(new_n1151), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1142), .B2(new_n1140), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1052), .A2(new_n1036), .ZN(new_n1164));
  INV_X1    g739(.A(G1996), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1103), .A2(new_n1164), .A3(new_n1165), .A4(new_n1045), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1102), .A2(KEYINPUT118), .A3(new_n1165), .A4(new_n1103), .ZN(new_n1169));
  XOR2_X1   g744(.A(KEYINPUT58), .B(G1341), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1081), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n554), .ZN(new_n1173));
  XOR2_X1   g748(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1172), .A2(KEYINPUT119), .A3(KEYINPUT59), .A4(new_n554), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(KEYINPUT61), .A3(new_n1141), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1163), .A2(new_n1175), .A3(new_n1176), .A4(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1153), .B1(new_n1161), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT54), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n475), .B1(new_n1041), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n471), .A2(KEYINPUT122), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1044), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT123), .B1(new_n1049), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n502), .A2(KEYINPUT105), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n499), .A2(new_n501), .A3(new_n923), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(G1384), .B1(new_n1193), .B2(new_n922), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1190), .B(new_n1187), .C1(new_n1194), .C2(KEYINPUT45), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1126), .B1(new_n926), .B2(new_n1037), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1189), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n1124), .A2(new_n1197), .A3(G301), .ZN(new_n1198));
  AOI21_X1  g773(.A(G301), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1183), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g777(.A(KEYINPUT124), .B(new_n1183), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1124), .A2(new_n1127), .A3(G301), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(KEYINPUT54), .ZN(new_n1206));
  AOI21_X1  g781(.A(G301), .B1(new_n1124), .B2(new_n1197), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1121), .A2(new_n1208), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1182), .A2(new_n1070), .A3(new_n1204), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1096), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1212));
  NOR2_X1   g787(.A1(G288), .A2(G1976), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1087), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI22_X1  g789(.A1(new_n1211), .A2(new_n1120), .B1(new_n1214), .B2(new_n1082), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT63), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1062), .A2(G8), .A3(G168), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1216), .B1(new_n1121), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(G8), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1216), .B1(new_n1219), .B2(new_n1100), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1217), .ZN(new_n1221));
  NAND4_X1  g796(.A1(new_n1220), .A2(new_n1096), .A3(new_n1120), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1215), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1130), .A2(new_n1210), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1049), .A2(new_n1045), .ZN(new_n1225));
  NOR3_X1   g800(.A1(new_n1225), .A2(new_n765), .A3(new_n1165), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1226), .B(KEYINPUT111), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1225), .A2(G1996), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n765), .ZN(new_n1229));
  AND2_X1   g804(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g805(.A(new_n803), .B(new_n805), .ZN(new_n1231));
  INV_X1    g806(.A(new_n1225), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1233), .A2(KEYINPUT112), .ZN(new_n1234));
  INV_X1    g809(.A(KEYINPUT112), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1231), .A2(new_n1235), .A3(new_n1232), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g812(.A(new_n870), .ZN(new_n1238));
  AND2_X1   g813(.A1(new_n1238), .A2(new_n872), .ZN(new_n1239));
  NOR2_X1   g814(.A1(new_n1238), .A2(new_n872), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1232), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  XOR2_X1   g816(.A(new_n597), .B(G1986), .Z(new_n1242));
  NAND2_X1  g817(.A1(new_n1242), .A2(new_n1232), .ZN(new_n1243));
  NAND4_X1  g818(.A1(new_n1230), .A2(new_n1237), .A3(new_n1241), .A4(new_n1243), .ZN(new_n1244));
  INV_X1    g819(.A(KEYINPUT113), .ZN(new_n1245));
  XNOR2_X1  g820(.A(new_n1244), .B(new_n1245), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1224), .A2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g822(.A1(new_n1237), .A2(new_n1239), .A3(new_n1227), .A4(new_n1229), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n803), .A2(new_n805), .ZN(new_n1249));
  AOI21_X1  g824(.A(new_n1225), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g825(.A(new_n1250), .ZN(new_n1251));
  NOR3_X1   g826(.A1(new_n1225), .A2(G1986), .A3(G290), .ZN(new_n1252));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1253));
  XNOR2_X1  g828(.A(new_n1252), .B(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g829(.A(new_n1254), .B(KEYINPUT48), .ZN(new_n1255));
  NAND4_X1  g830(.A1(new_n1255), .A2(new_n1237), .A3(new_n1230), .A4(new_n1241), .ZN(new_n1256));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1257));
  INV_X1    g832(.A(KEYINPUT46), .ZN(new_n1258));
  XNOR2_X1  g833(.A(new_n1228), .B(new_n1258), .ZN(new_n1259));
  OAI21_X1  g834(.A(new_n1232), .B1(new_n1231), .B2(new_n941), .ZN(new_n1260));
  NAND2_X1  g835(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  XOR2_X1   g836(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1262));
  AND2_X1   g837(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g838(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1264));
  OR2_X1    g839(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g840(.A1(new_n1251), .A2(new_n1256), .A3(new_n1257), .A4(new_n1265), .ZN(new_n1266));
  NAND3_X1  g841(.A1(new_n1230), .A2(new_n1237), .A3(new_n1241), .ZN(new_n1267));
  INV_X1    g842(.A(KEYINPUT48), .ZN(new_n1268));
  XNOR2_X1  g843(.A(new_n1254), .B(new_n1268), .ZN(new_n1269));
  OAI22_X1  g844(.A1(new_n1267), .A2(new_n1269), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1270));
  OAI21_X1  g845(.A(KEYINPUT127), .B1(new_n1270), .B2(new_n1250), .ZN(new_n1271));
  NAND2_X1  g846(.A1(new_n1266), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g847(.A1(new_n1247), .A2(new_n1272), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g848(.A1(G227), .A2(new_n463), .ZN(new_n1275));
  AND3_X1   g849(.A1(new_n706), .A2(new_n661), .A3(new_n1275), .ZN(new_n1276));
  AND3_X1   g850(.A1(new_n1276), .A2(new_n957), .A3(new_n1028), .ZN(G308));
  NAND3_X1  g851(.A1(new_n1276), .A2(new_n957), .A3(new_n1028), .ZN(G225));
endmodule


