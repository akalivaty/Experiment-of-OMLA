//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n204));
  NAND2_X1  g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(KEYINPUT15), .B2(new_n203), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT86), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n210), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n204), .B1(new_n218), .B2(new_n205), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n202), .B1(new_n220), .B2(KEYINPUT87), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n218), .A2(new_n205), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n222), .A2(new_n204), .B1(new_n206), .B2(new_n213), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT87), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT17), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G22gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G15gat), .ZN(new_n228));
  INV_X1    g027(.A(G15gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G22gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT88), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(G15gat), .B(G22gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(KEYINPUT16), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n234), .B1(new_n233), .B2(new_n237), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT89), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n239), .B2(new_n240), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n233), .A2(new_n237), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G8gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT89), .A3(new_n238), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT90), .B1(new_n249), .B2(new_n223), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT90), .ZN(new_n251));
  AOI211_X1 g050(.A(new_n251), .B(new_n220), .C1(new_n245), .C2(new_n248), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n242), .B(new_n243), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT91), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n243), .B(KEYINPUT13), .Z(new_n257));
  NAND3_X1  g056(.A1(new_n245), .A2(new_n248), .A3(new_n220), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT92), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n250), .A2(new_n252), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n249), .A2(new_n223), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n251), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n249), .A2(KEYINPUT90), .A3(new_n223), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n255), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n265), .A2(new_n243), .A3(new_n242), .A4(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n256), .A2(new_n261), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G141gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G197gat), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT11), .B(G169gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT12), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n256), .A2(new_n261), .A3(new_n267), .A4(new_n273), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT24), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(G183gat), .B2(G190gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT23), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT25), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT64), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT65), .B(G190gat), .ZN(new_n304));
  INV_X1    g103(.A(G183gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n290), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(KEYINPUT25), .A3(new_n297), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n301), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT27), .B(G183gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT28), .Z(new_n312));
  INV_X1    g111(.A(KEYINPUT26), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n292), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT66), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n315), .B(new_n294), .C1(new_n313), .C2(new_n292), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n286), .A3(new_n316), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n309), .A2(KEYINPUT72), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT72), .B1(new_n309), .B2(new_n317), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n283), .B(new_n285), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT22), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n321), .A2(KEYINPUT69), .B1(G211gat), .B2(G218gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(KEYINPUT69), .B2(new_n321), .ZN(new_n323));
  XNOR2_X1  g122(.A(G197gat), .B(G204gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(G211gat), .B(G218gat), .Z(new_n326));
  INV_X1    g125(.A(KEYINPUT70), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n325), .B(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT71), .ZN(new_n330));
  INV_X1    g129(.A(new_n318), .ZN(new_n331));
  INV_X1    g130(.A(new_n319), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n284), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n309), .A2(new_n317), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT73), .B1(new_n336), .B2(new_n284), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n320), .B(new_n330), .C1(new_n333), .C2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n329), .B(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n309), .A2(new_n285), .A3(new_n317), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n318), .A2(new_n319), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n284), .A2(new_n335), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n340), .B(new_n341), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n282), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT74), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G155gat), .B(G162gat), .ZN(new_n352));
  XOR2_X1   g151(.A(G141gat), .B(G148gat), .Z(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(KEYINPUT75), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n355));
  AND2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n357), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G127gat), .B(G134gat), .Z(new_n361));
  XNOR2_X1  g160(.A(G113gat), .B(G120gat), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n361), .A2(KEYINPUT1), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G127gat), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n364), .A2(G134gat), .ZN(new_n365));
  MUX2_X1   g164(.A(new_n365), .B(new_n361), .S(KEYINPUT67), .Z(new_n366));
  AOI21_X1  g165(.A(KEYINPUT1), .B1(new_n362), .B2(KEYINPUT68), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(KEYINPUT68), .B2(new_n362), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n363), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n360), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n369), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n358), .A2(new_n359), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n373), .A3(KEYINPUT77), .ZN(new_n374));
  OR3_X1    g173(.A1(new_n360), .A2(KEYINPUT77), .A3(new_n369), .ZN(new_n375));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT5), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n360), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT4), .B1(new_n360), .B2(new_n369), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n369), .B1(new_n360), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT76), .B1(new_n372), .B2(KEYINPUT3), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n386));
  AOI211_X1 g185(.A(new_n386), .B(new_n383), .C1(new_n358), .C2(new_n359), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n384), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(new_n388), .A3(new_n376), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n379), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G1gat), .B(G29gat), .Z(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n382), .A2(new_n388), .A3(KEYINPUT5), .A4(new_n376), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n390), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n395), .B1(new_n390), .B2(new_n396), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n398), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n338), .A2(new_n344), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(new_n281), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(KEYINPUT30), .B2(new_n345), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n351), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  INV_X1    g207(.A(G50gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G22gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n325), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n328), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n325), .B1(new_n327), .B2(new_n326), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n335), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT3), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT81), .B(new_n335), .C1(new_n415), .C2(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n372), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n335), .B1(new_n372), .B2(KEYINPUT3), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n330), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n413), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n335), .B1(new_n414), .B2(new_n326), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n326), .B2(new_n414), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n372), .B1(new_n427), .B2(KEYINPUT3), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n413), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n425), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n360), .B1(new_n419), .B2(new_n420), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT29), .B1(new_n360), .B2(new_n383), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n340), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(G228gat), .B(G233gat), .C1(new_n434), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n433), .B1(new_n437), .B2(new_n429), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n412), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n431), .B1(new_n425), .B2(new_n430), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n429), .A3(new_n433), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n411), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n334), .A2(new_n369), .ZN(new_n446));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n309), .A2(new_n371), .A3(new_n317), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n450), .A2(KEYINPUT32), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(G15gat), .B(G43gat), .Z(new_n454));
  XNOR2_X1  g253(.A(G71gat), .B(G99gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT34), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n446), .A2(new_n449), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(new_n447), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n458), .A3(new_n447), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n456), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n450), .B2(new_n452), .ZN(new_n465));
  INV_X1    g264(.A(new_n462), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(new_n460), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n451), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n463), .A2(new_n467), .A3(new_n451), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(KEYINPUT36), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT36), .ZN(new_n472));
  INV_X1    g271(.A(new_n470), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n468), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n407), .A2(new_n445), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n381), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n360), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n371), .B1(KEYINPUT3), .B2(new_n372), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n386), .B1(new_n360), .B2(new_n383), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n372), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n377), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n377), .B1(new_n374), .B2(new_n375), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n485), .A2(KEYINPUT84), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n382), .A2(new_n388), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n377), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n485), .B2(KEYINPUT84), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n484), .A2(new_n486), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n487), .B2(new_n377), .ZN(new_n493));
  AOI211_X1 g292(.A(KEYINPUT83), .B(new_n376), .C1(new_n382), .C2(new_n388), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n395), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT40), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT85), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n397), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n489), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n395), .B1(new_n501), .B2(new_n490), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n502), .B2(new_n492), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n345), .A2(new_n349), .ZN(new_n505));
  AOI211_X1 g304(.A(KEYINPUT74), .B(new_n282), .C1(new_n338), .C2(new_n344), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT30), .ZN(new_n507));
  INV_X1    g306(.A(new_n405), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n346), .B2(new_n348), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n281), .B1(new_n404), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n338), .A2(KEYINPUT37), .A3(new_n344), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT38), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n402), .A2(new_n401), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n399), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n505), .A2(new_n506), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n320), .B1(new_n333), .B2(new_n337), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n340), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n511), .B1(new_n521), .B2(new_n330), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT38), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n515), .A2(new_n517), .A3(new_n518), .A4(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n443), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n475), .A2(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n443), .A2(new_n473), .A3(new_n468), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT35), .B1(new_n407), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n507), .A2(new_n509), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT35), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n403), .A4(new_n529), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n278), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G183gat), .B(G211gat), .Z(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G127gat), .B(G155gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT96), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT9), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G64gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(G57gat), .ZN(new_n546));
  INV_X1    g345(.A(G57gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(G64gat), .ZN(new_n548));
  OAI211_X1 g347(.A(KEYINPUT94), .B(new_n544), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G71gat), .B(G78gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(KEYINPUT93), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(G64gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n545), .A2(G57gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n553), .A2(new_n554), .B1(new_n543), .B2(new_n542), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(new_n555), .B2(KEYINPUT94), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n552), .B(new_n544), .C1(new_n546), .C2(new_n548), .ZN(new_n557));
  INV_X1    g356(.A(new_n550), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n551), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT95), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n562), .B(new_n551), .C1(new_n556), .C2(new_n559), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(G231gat), .B(G233gat), .C1(new_n564), .C2(KEYINPUT21), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n541), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n541), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n538), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n572), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n574), .A2(new_n537), .A3(new_n570), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n248), .B(new_n245), .C1(new_n565), .C2(new_n566), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(new_n575), .B2(new_n573), .ZN(new_n582));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT7), .ZN(new_n586));
  XNOR2_X1  g385(.A(G99gat), .B(G106gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(KEYINPUT8), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n587), .B1(new_n586), .B2(new_n591), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n223), .A2(new_n594), .B1(KEYINPUT41), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT98), .ZN(new_n598));
  INV_X1    g397(.A(new_n594), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n226), .B2(new_n599), .ZN(new_n600));
  AOI211_X1 g399(.A(KEYINPUT98), .B(new_n594), .C1(new_n221), .C2(new_n225), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(KEYINPUT99), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n584), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT97), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(KEYINPUT99), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND3_X1  g410(.A1(new_n602), .A2(new_n605), .A3(new_n584), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n607), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n611), .ZN(new_n614));
  INV_X1    g413(.A(new_n612), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(new_n606), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n580), .A2(new_n582), .A3(new_n613), .A4(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n561), .A2(new_n563), .A3(new_n599), .ZN(new_n619));
  INV_X1    g418(.A(new_n593), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n592), .B1(new_n620), .B2(KEYINPUT100), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n593), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n623), .A3(new_n560), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n618), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  AOI211_X1 g427(.A(KEYINPUT101), .B(new_n626), .C1(new_n619), .C2(new_n624), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n619), .A2(new_n631), .A3(new_n624), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n564), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n626), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  NAND3_X1  g437(.A1(new_n630), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n634), .B2(new_n626), .ZN(new_n641));
  AOI211_X1 g440(.A(KEYINPUT102), .B(new_n627), .C1(new_n632), .C2(new_n633), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n630), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n644));
  INV_X1    g443(.A(new_n638), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n643), .B2(new_n645), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n639), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n617), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n536), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n403), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n232), .ZN(G1324gat));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  OAI21_X1  g452(.A(G8gat), .B1(new_n650), .B2(new_n532), .ZN(new_n654));
  INV_X1    g453(.A(new_n532), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  NAND4_X1  g455(.A1(new_n536), .A2(new_n655), .A3(new_n649), .A4(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n653), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n658), .A2(KEYINPUT104), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT104), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(G1325gat));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n471), .A2(new_n474), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n664), .B1(new_n471), .B2(new_n474), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(G15gat), .B1(new_n650), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n473), .A2(new_n468), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n229), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n650), .B2(new_n670), .ZN(G1326gat));
  INV_X1    g470(.A(new_n445), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n650), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT43), .B(G22gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NAND2_X1  g474(.A1(new_n580), .A2(new_n582), .ZN(new_n676));
  INV_X1    g475(.A(new_n639), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n625), .A2(new_n627), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT101), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n625), .A2(new_n618), .A3(new_n627), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n635), .A2(KEYINPUT102), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n634), .A2(new_n640), .A3(new_n626), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT103), .B1(new_n684), .B2(new_n638), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n677), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n676), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n616), .A2(new_n613), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n536), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n208), .A3(new_n517), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n528), .A2(new_n535), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n688), .A2(new_n278), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n407), .A2(new_n445), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n667), .A2(new_n527), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n690), .B1(new_n700), .B2(new_n535), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n697), .B(new_n698), .C1(new_n701), .C2(KEYINPUT44), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(KEYINPUT106), .A3(new_n403), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT106), .B1(new_n702), .B2(new_n403), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G29gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n694), .B1(new_n703), .B2(new_n705), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n532), .A2(G36gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n692), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n536), .A2(new_n691), .ZN(new_n711));
  INV_X1    g510(.A(new_n709), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT107), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n707), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n710), .A2(new_n707), .A3(new_n713), .ZN(new_n717));
  OAI21_X1  g516(.A(G36gat), .B1(new_n702), .B2(new_n532), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n718), .ZN(G1329gat));
  OAI21_X1  g518(.A(G43gat), .B1(new_n702), .B2(new_n667), .ZN(new_n720));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n692), .A2(new_n721), .A3(new_n669), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1330gat));
  NAND2_X1  g524(.A1(new_n445), .A2(new_n409), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n692), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n727), .B2(new_n692), .ZN(new_n729));
  OAI21_X1  g528(.A(G50gat), .B1(new_n702), .B2(new_n526), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(KEYINPUT48), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G50gat), .B1(new_n702), .B2(new_n672), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g533(.A1(new_n700), .A2(new_n535), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n617), .A2(new_n277), .A3(new_n687), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n517), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G57gat), .ZN(G1332gat));
  INV_X1    g538(.A(KEYINPUT49), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n655), .B1(new_n740), .B2(new_n545), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT110), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n545), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n667), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n737), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n737), .A2(KEYINPUT111), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n669), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n746), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n752), .B2(new_n754), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(G1334gat));
  NAND2_X1  g557(.A1(new_n737), .A2(new_n445), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n676), .A2(new_n278), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n701), .A2(KEYINPUT51), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT51), .B1(new_n701), .B2(new_n762), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(new_n687), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n589), .A3(new_n517), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n761), .A2(new_n687), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n697), .B(new_n768), .C1(new_n701), .C2(KEYINPUT44), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n403), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(G1336gat));
  NOR2_X1   g570(.A1(new_n532), .A2(G92gat), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n648), .B(new_n772), .C1(new_n763), .C2(new_n764), .ZN(new_n773));
  OAI21_X1  g572(.A(G92gat), .B1(new_n769), .B2(new_n532), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n773), .B(new_n774), .C1(new_n776), .C2(KEYINPUT52), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n769), .B2(new_n667), .ZN(new_n782));
  INV_X1    g581(.A(G99gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n669), .A2(new_n783), .A3(new_n648), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n765), .B2(new_n784), .ZN(G1338gat));
  NOR2_X1   g584(.A1(new_n526), .A2(G106gat), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n648), .B(new_n786), .C1(new_n763), .C2(new_n764), .ZN(new_n787));
  OAI21_X1  g586(.A(G106gat), .B1(new_n769), .B2(new_n526), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n769), .A2(new_n672), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n766), .A2(new_n786), .B1(new_n791), .B2(G106gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n792), .B2(new_n789), .ZN(G1339gat));
  NAND2_X1  g592(.A1(new_n649), .A2(new_n278), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT114), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n649), .A2(new_n796), .A3(new_n278), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n682), .A2(new_n799), .A3(new_n683), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n632), .A2(new_n627), .A3(new_n633), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n635), .A2(KEYINPUT54), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n645), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n645), .A4(new_n802), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n639), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n259), .A2(new_n260), .A3(new_n257), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n243), .B1(new_n265), .B2(new_n242), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n272), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n276), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n809), .A2(new_n689), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n648), .A2(new_n814), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n277), .A2(new_n805), .A3(new_n639), .A4(new_n807), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n689), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT115), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n676), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n798), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n517), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n655), .A3(new_n530), .ZN(new_n827));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n277), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n655), .A2(new_n403), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n669), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n825), .A2(new_n831), .A3(new_n672), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n831), .B1(new_n825), .B2(new_n672), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT117), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n837), .B(new_n830), .C1(new_n833), .C2(new_n834), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n277), .A2(G113gat), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n828), .B1(new_n839), .B2(new_n840), .ZN(G1340gat));
  AOI21_X1  g640(.A(G120gat), .B1(new_n827), .B2(new_n648), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n648), .A2(G120gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n839), .B2(new_n843), .ZN(G1341gat));
  NAND3_X1  g643(.A1(new_n836), .A2(new_n824), .A3(new_n838), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G127gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n364), .A3(new_n824), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1342gat));
  NAND3_X1  g647(.A1(new_n836), .A2(new_n689), .A3(new_n838), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G134gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n532), .A2(new_n689), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT118), .ZN(new_n852));
  NOR4_X1   g651(.A1(new_n826), .A2(G134gat), .A3(new_n530), .A4(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT56), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n850), .A2(new_n854), .ZN(G1343gat));
  AND2_X1   g654(.A1(new_n829), .A2(new_n667), .ZN(new_n856));
  INV_X1    g655(.A(G141gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n278), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n687), .A2(KEYINPUT119), .A3(new_n813), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n648), .B2(new_n814), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT120), .B1(new_n806), .B2(new_n808), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n805), .A2(new_n864), .A3(new_n639), .A4(new_n807), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n277), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n689), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n676), .B1(new_n867), .B2(new_n816), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n798), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n672), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AND4_X1   g674(.A1(new_n277), .A2(new_n805), .A3(new_n639), .A4(new_n807), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n685), .A2(new_n686), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n813), .B1(new_n877), .B2(new_n639), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n820), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n690), .A3(new_n822), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n824), .B1(new_n880), .B2(new_n815), .ZN(new_n881));
  INV_X1    g680(.A(new_n797), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n796), .B1(new_n649), .B2(new_n278), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n443), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n870), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n872), .B2(new_n873), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n856), .B(new_n858), .C1(new_n875), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n889));
  NOR2_X1   g688(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n825), .A2(new_n517), .ZN(new_n891));
  INV_X1    g690(.A(new_n667), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n526), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n891), .A2(new_n277), .A3(new_n532), .A4(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n890), .B1(new_n894), .B2(new_n857), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n888), .A2(new_n889), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n889), .B1(new_n888), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(G1344gat));
  NAND3_X1  g697(.A1(new_n891), .A2(new_n532), .A3(new_n893), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n687), .A2(G148gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT123), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G148gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n856), .ZN(new_n905));
  AOI211_X1 g704(.A(new_n870), .B(new_n672), .C1(new_n868), .C2(new_n798), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n906), .A2(KEYINPUT121), .B1(new_n870), .B2(new_n885), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n907), .B2(new_n874), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n904), .B1(new_n908), .B2(new_n648), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n868), .A2(new_n794), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n445), .A2(new_n870), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI22_X1  g711(.A1(KEYINPUT57), .A2(new_n885), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n648), .A3(new_n856), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n903), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n902), .B1(new_n909), .B2(new_n915), .ZN(G1345gat));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n899), .A2(new_n917), .A3(new_n676), .ZN(new_n918));
  INV_X1    g717(.A(G155gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n899), .B2(new_n676), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n908), .A2(G155gat), .A3(new_n824), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n689), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G162gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n852), .A2(G162gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n891), .A2(new_n893), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1347gat));
  AND2_X1   g727(.A1(new_n825), .A2(new_n403), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n655), .A3(new_n529), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n277), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n655), .A2(new_n403), .A3(new_n669), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n825), .A2(new_n672), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT116), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n935), .B2(new_n832), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n277), .A2(G169gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(G1348gat));
  AOI21_X1  g737(.A(G176gat), .B1(new_n931), .B2(new_n648), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n648), .A2(G176gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n936), .B2(new_n940), .ZN(G1349gat));
  NAND3_X1  g740(.A1(new_n931), .A2(new_n310), .A3(new_n824), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n305), .B1(new_n936), .B2(new_n824), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT60), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n936), .A2(new_n824), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n946), .B(new_n942), .C1(new_n947), .C2(new_n305), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n304), .A3(new_n689), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n936), .A2(new_n689), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n951), .A2(new_n952), .A3(G190gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n951), .B2(G190gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(G1351gat));
  NOR3_X1   g754(.A1(new_n892), .A2(new_n532), .A3(new_n526), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n929), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n277), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n870), .B1(new_n825), .B2(new_n443), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n911), .B1(new_n868), .B2(new_n794), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n667), .A2(new_n403), .A3(new_n655), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n277), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  NOR2_X1   g764(.A1(new_n687), .A2(G204gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n929), .A2(new_n956), .A3(new_n966), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(G204gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n971), .B1(new_n963), .B2(new_n648), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT125), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(new_n972), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n974), .A2(new_n975), .A3(new_n969), .A4(new_n968), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n976), .ZN(G1353gat));
  INV_X1    g776(.A(G211gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n958), .A2(new_n978), .A3(new_n824), .ZN(new_n979));
  NOR4_X1   g778(.A1(new_n960), .A2(new_n961), .A3(new_n676), .A4(new_n962), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n885), .A2(KEYINPUT57), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n910), .A2(new_n912), .ZN(new_n984));
  INV_X1    g783(.A(new_n962), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n983), .A2(new_n984), .A3(new_n824), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT126), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n913), .A2(new_n981), .A3(new_n824), .A4(new_n985), .ZN(new_n989));
  AND4_X1   g788(.A1(KEYINPUT63), .A2(new_n987), .A3(new_n989), .A4(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n979), .B1(new_n988), .B2(new_n990), .ZN(G1354gat));
  NAND3_X1  g790(.A1(new_n913), .A2(new_n689), .A3(new_n985), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G218gat), .ZN(new_n993));
  OR3_X1    g792(.A1(new_n957), .A2(G218gat), .A3(new_n690), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(G1355gat));
endmodule


