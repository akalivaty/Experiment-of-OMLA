//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1321,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n201), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n203), .A2(G50), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT66), .Z(new_n229));
  AND2_X1   g0029(.A1(KEYINPUT65), .A2(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(KEYINPUT65), .A2(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n215), .A2(new_n227), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n222), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NAND3_X1  g0054(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT71), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n257), .A2(new_n209), .A3(G13), .A4(G20), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT70), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT70), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n262), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n233), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n209), .B2(G20), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n265), .A2(new_n269), .B1(new_n259), .B2(new_n268), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G58), .A2(G68), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT77), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT77), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G58), .A3(G68), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(new_n203), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n275), .A2(G20), .B1(G159), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n278), .A2(new_n279), .A3(G20), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT7), .ZN(new_n281));
  OAI21_X1  g0081(.A(G68), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT65), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n210), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT65), .A2(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n286), .A2(new_n291), .A3(KEYINPUT7), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n277), .B(KEYINPUT16), .C1(new_n282), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n264), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT7), .B1(new_n286), .B2(new_n291), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n278), .A2(new_n279), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(new_n281), .A3(new_n210), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(G68), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT16), .B1(new_n298), .B2(new_n277), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n270), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  INV_X1    g0101(.A(new_n233), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n303), .A2(G1), .A3(G13), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n305), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n307), .B1(new_n222), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G226), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n289), .B2(new_n290), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(G1698), .B1(G33), .B2(G87), .ZN(new_n313));
  INV_X1    g0113(.A(G1698), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT69), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT69), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G1698), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n315), .B(new_n317), .C1(new_n278), .C2(new_n279), .ZN(new_n318));
  INV_X1    g0118(.A(G223), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT78), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT69), .B(G1698), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT78), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n291), .A2(new_n321), .A3(new_n322), .A4(G223), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n313), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n310), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n326), .A2(G200), .ZN(new_n327));
  AOI211_X1 g0127(.A(G190), .B(new_n310), .C1(new_n324), .C2(new_n325), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n300), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT17), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  AOI211_X1 g0134(.A(new_n334), .B(new_n310), .C1(new_n324), .C2(new_n325), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n300), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT18), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n298), .A2(new_n277), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(new_n264), .A3(new_n293), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n326), .A2(G200), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n341), .B(new_n270), .C1(new_n342), .C2(new_n328), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT18), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n300), .B(new_n346), .C1(new_n333), .C2(new_n335), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n331), .A2(new_n337), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n261), .A2(new_n233), .A3(new_n263), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n256), .A2(new_n258), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n209), .A2(G20), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n350), .A2(new_n351), .A3(G68), .A4(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT12), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n259), .B2(new_n202), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n351), .A2(KEYINPUT12), .A3(G68), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n357), .A2(KEYINPUT76), .ZN(new_n358));
  OAI211_X1 g0158(.A(G232), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  OAI21_X1  g0160(.A(G226), .B1(new_n278), .B2(new_n279), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n315), .A2(new_n317), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n359), .B(new_n360), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n325), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  INV_X1    g0165(.A(new_n309), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(G238), .B1(new_n304), .B2(new_n306), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n365), .B1(new_n364), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g0169(.A(G200), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n276), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n284), .A2(G33), .A3(new_n285), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n206), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n264), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT11), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(KEYINPUT11), .A3(new_n264), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(KEYINPUT76), .B2(new_n357), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n364), .A2(new_n367), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT13), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(G190), .A3(new_n382), .ZN(new_n383));
  AND4_X1   g0183(.A1(new_n358), .A2(new_n370), .A3(new_n379), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n379), .A2(new_n358), .ZN(new_n385));
  OAI21_X1  g0185(.A(G169), .B1(new_n368), .B2(new_n369), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT14), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n381), .A2(G179), .A3(new_n382), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT14), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n389), .B(G169), .C1(new_n368), .C2(new_n369), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n384), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT73), .B1(new_n351), .B2(G77), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT73), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n256), .A2(new_n394), .A3(new_n206), .A4(new_n258), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n276), .B1(new_n266), .B2(new_n267), .ZN(new_n397));
  OAI21_X1  g0197(.A(G77), .B1(new_n230), .B2(new_n231), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g0199(.A(KEYINPUT15), .B(G87), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n372), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n264), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n206), .B1(new_n209), .B2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n350), .A2(new_n351), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n396), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n314), .B1(new_n289), .B2(new_n290), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(G238), .B1(new_n296), .B2(G107), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n291), .A2(new_n321), .A3(G232), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n308), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G244), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n307), .B1(new_n413), .B2(new_n309), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(G190), .A3(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n396), .A2(new_n402), .A3(KEYINPUT74), .A4(new_n404), .ZN(new_n417));
  OAI21_X1  g0217(.A(G200), .B1(new_n411), .B2(new_n414), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n407), .A2(new_n416), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n411), .A2(G179), .A3(new_n414), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n412), .A2(new_n415), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n332), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n407), .A2(new_n417), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n349), .A2(new_n392), .A3(new_n419), .A4(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n291), .B1(new_n319), .B2(new_n314), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(G222), .B2(new_n321), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n325), .B1(new_n291), .B2(G77), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n307), .B1(new_n311), .B2(new_n309), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G179), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n332), .B2(new_n429), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n205), .A2(new_n210), .ZN(new_n432));
  INV_X1    g0232(.A(G150), .ZN(new_n433));
  INV_X1    g0233(.A(new_n276), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n268), .A2(new_n372), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n264), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n350), .A2(new_n351), .A3(G50), .A4(new_n352), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  INV_X1    g0238(.A(G50), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n259), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n437), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n436), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n431), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(KEYINPUT9), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT9), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n436), .B(new_n446), .C1(new_n442), .C2(new_n441), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT10), .ZN(new_n449));
  INV_X1    g0249(.A(G190), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT75), .B1(new_n429), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(G200), .B2(new_n429), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n448), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n449), .B1(new_n448), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n444), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n209), .A2(G33), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n350), .A2(new_n351), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n259), .A2(KEYINPUT25), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT25), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n351), .B2(G107), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n458), .A2(G107), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n291), .A2(new_n232), .A3(G87), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT22), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT22), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n291), .A2(new_n232), .A3(new_n468), .A4(G87), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT23), .A2(G107), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(G20), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT23), .A2(G107), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n286), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n465), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n465), .A3(new_n475), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n464), .B1(new_n479), .B2(new_n264), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT88), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G294), .ZN(new_n482));
  INV_X1    g0282(.A(G294), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(KEYINPUT88), .ZN(new_n484));
  OAI21_X1  g0284(.A(G33), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(G257), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n486), .C1(new_n318), .C2(new_n219), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n325), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT5), .B(G41), .ZN(new_n489));
  INV_X1    g0289(.A(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G1), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n489), .A2(new_n491), .B1(new_n302), .B2(new_n303), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G264), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n489), .A2(G274), .A3(new_n308), .A4(new_n491), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n488), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT89), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n487), .A2(new_n325), .B1(G264), .B2(new_n492), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT89), .B1(new_n498), .B2(new_n494), .ZN(new_n499));
  OAI211_X1 g0299(.A(KEYINPUT91), .B(new_n450), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G200), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n495), .A2(new_n496), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n498), .A2(KEYINPUT89), .A3(new_n494), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT91), .B1(new_n506), .B2(new_n450), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n480), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n504), .A2(G169), .A3(new_n505), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n498), .A2(G179), .A3(new_n494), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT90), .B1(new_n511), .B2(new_n480), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n479), .A2(new_n264), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n463), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n509), .A2(new_n510), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT90), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n508), .A2(new_n512), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n289), .A2(G303), .A3(new_n290), .ZN(new_n519));
  OAI211_X1 g0319(.A(G264), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n520), .C1(new_n318), .C2(new_n224), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n325), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n209), .A2(G45), .ZN(new_n523));
  AND2_X1   g0323(.A1(KEYINPUT5), .A2(G41), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT5), .A2(G41), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n523), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n492), .A2(G270), .B1(new_n528), .B2(new_n304), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n522), .A2(new_n529), .A3(G190), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n491), .B1(new_n524), .B2(new_n526), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G270), .A3(new_n308), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n494), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n325), .B2(new_n521), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n530), .B1(new_n534), .B2(new_n501), .ZN(new_n535));
  AND2_X1   g0335(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n210), .A2(G116), .ZN(new_n539));
  INV_X1    g0339(.A(G283), .ZN(new_n540));
  MUX2_X1   g0340(.A(new_n223), .B(new_n540), .S(G33), .Z(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(new_n232), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n538), .B1(new_n542), .B2(new_n264), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n288), .A2(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G283), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n284), .A2(new_n544), .A3(new_n285), .A4(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n539), .ZN(new_n547));
  AND4_X1   g0347(.A1(new_n264), .A2(new_n538), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n537), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n350), .A2(new_n351), .A3(G116), .A4(new_n456), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT85), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n351), .B2(G116), .ZN(new_n552));
  INV_X1    g0352(.A(G116), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n256), .A2(KEYINPUT85), .A3(new_n553), .A4(new_n258), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n535), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n332), .B1(new_n522), .B2(new_n529), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT21), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT87), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n558), .A2(KEYINPUT21), .B1(new_n534), .B2(G179), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n264), .A2(new_n546), .A3(new_n547), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(KEYINPUT86), .B2(KEYINPUT20), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n542), .A2(new_n264), .A3(new_n538), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n562), .B1(new_n566), .B2(new_n537), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n560), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  AOI211_X1 g0369(.A(new_n569), .B(new_n332), .C1(new_n522), .C2(new_n529), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n522), .A2(new_n529), .A3(G179), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n556), .B(KEYINPUT87), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  AOI211_X1 g0373(.A(new_n557), .B(new_n559), .C1(new_n568), .C2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT83), .ZN(new_n575));
  INV_X1    g0375(.A(new_n400), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n458), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n372), .B2(new_n223), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n218), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n360), .A2(new_n578), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n286), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n291), .A2(new_n232), .A3(G68), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n579), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n264), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT83), .B1(new_n457), .B2(new_n400), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n259), .A2(new_n400), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n577), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n325), .A2(new_n219), .A3(new_n491), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n308), .A2(G274), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT82), .B1(new_n591), .B2(new_n523), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT82), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n304), .A2(new_n593), .A3(new_n491), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n590), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G116), .ZN(new_n596));
  OAI211_X1 g0396(.A(G244), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n318), .C2(new_n217), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n325), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n600), .A2(new_n334), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n332), .B1(new_n595), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n589), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT84), .B1(new_n600), .B2(new_n450), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n350), .A2(new_n351), .A3(G87), .A4(new_n456), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n586), .A2(new_n588), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT84), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n595), .A2(new_n599), .A3(new_n607), .A4(G190), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n600), .A2(G200), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n604), .A2(new_n606), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT79), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT6), .ZN(new_n614));
  AND2_X1   g0414(.A1(G97), .A2(G107), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n580), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n459), .A2(KEYINPUT6), .A3(G97), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n232), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n434), .A2(new_n206), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n613), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n619), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n459), .A2(KEYINPUT6), .A3(G97), .ZN(new_n622));
  XNOR2_X1  g0422(.A(G97), .B(G107), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n623), .B2(new_n614), .ZN(new_n624));
  OAI211_X1 g0424(.A(KEYINPUT79), .B(new_n621), .C1(new_n624), .C2(new_n232), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n295), .A2(G107), .A3(new_n297), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n620), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n264), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n457), .A2(G97), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n351), .A2(new_n223), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT4), .ZN(new_n633));
  OAI21_X1  g0433(.A(G244), .B1(new_n278), .B2(new_n279), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(new_n362), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n291), .A2(new_n321), .A3(KEYINPUT4), .A4(G244), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n408), .A2(G250), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .A4(new_n545), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n325), .ZN(new_n639));
  INV_X1    g0439(.A(new_n494), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n531), .A2(G257), .A3(new_n308), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT80), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n531), .A2(KEYINPUT80), .A3(G257), .A4(new_n308), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n639), .A2(new_n645), .A3(new_n334), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n639), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n332), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n632), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n627), .A2(new_n264), .B1(new_n629), .B2(new_n630), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n639), .A2(new_n645), .A3(new_n450), .ZN(new_n651));
  AOI21_X1  g0451(.A(G200), .B1(new_n639), .B2(new_n645), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT81), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n649), .A2(KEYINPUT81), .A3(new_n653), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n574), .B(new_n612), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  NOR4_X1   g0457(.A1(new_n425), .A2(new_n455), .A3(new_n518), .A4(new_n657), .ZN(G372));
  AND2_X1   g0458(.A1(new_n331), .A2(new_n345), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n390), .A2(new_n388), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n381), .A2(new_n382), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n389), .B1(new_n661), .B2(G169), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n385), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n384), .B2(new_n424), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n337), .A2(new_n347), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n453), .A2(new_n454), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n667), .A2(new_n668), .B1(new_n443), .B2(new_n431), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT92), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n425), .A2(new_n455), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n649), .A2(new_n653), .A3(new_n603), .A4(new_n610), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n511), .A2(new_n480), .ZN(new_n674));
  INV_X1    g0474(.A(new_n559), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n567), .B2(new_n561), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n508), .B(new_n673), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n611), .B2(new_n649), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n632), .A2(new_n646), .A3(new_n648), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(KEYINPUT26), .A3(new_n603), .A4(new_n610), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n601), .A2(new_n602), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n679), .A2(new_n681), .B1(new_n682), .B2(new_n589), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n671), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n670), .A2(new_n685), .ZN(G369));
  NAND2_X1  g0486(.A1(new_n209), .A2(G13), .ZN(new_n687));
  OR3_X1    g0487(.A1(new_n286), .A2(KEYINPUT27), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT27), .B1(new_n286), .B2(new_n687), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n574), .B1(new_n567), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n676), .A2(new_n556), .A3(new_n692), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n514), .A2(new_n692), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n508), .A2(new_n512), .A3(new_n517), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n674), .A2(new_n692), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n511), .A2(new_n480), .A3(new_n692), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n568), .A2(new_n573), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT93), .B(new_n693), .C1(new_n705), .C2(new_n559), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT93), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n559), .B1(new_n568), .B2(new_n573), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n692), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n704), .B1(new_n702), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n703), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n213), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n581), .A2(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n229), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n715), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n692), .B1(new_n677), .B2(new_n683), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n512), .A2(new_n517), .A3(new_n708), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n450), .B1(new_n497), .B2(new_n499), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT91), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n502), .A3(new_n500), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n672), .B1(new_n727), .B2(new_n480), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n679), .A2(new_n681), .A3(KEYINPUT96), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT96), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n612), .A2(new_n731), .A3(KEYINPUT26), .A4(new_n680), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n603), .A3(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(KEYINPUT29), .B(new_n693), .C1(new_n729), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n722), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n657), .A2(new_n518), .A3(new_n692), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n498), .A2(new_n599), .A3(new_n595), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n737), .A2(new_n647), .A3(new_n571), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT95), .B1(new_n738), .B2(KEYINPUT30), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT95), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n572), .A2(new_n498), .A3(new_n599), .A4(new_n595), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n740), .B(new_n741), .C1(new_n742), .C2(new_n647), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n738), .A2(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n522), .A2(new_n529), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n600), .A2(new_n745), .A3(new_n334), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT94), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT94), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n600), .A2(new_n745), .A3(new_n748), .A4(new_n334), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n747), .A2(new_n495), .A3(new_n647), .A4(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n739), .A2(new_n743), .A3(new_n744), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n692), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n741), .B1(new_n742), .B2(new_n647), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(new_n744), .A3(new_n750), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n693), .A2(new_n753), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(G330), .B1(new_n736), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n735), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n720), .B1(new_n762), .B2(G1), .ZN(G364));
  AND2_X1   g0563(.A1(new_n232), .A2(G13), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G45), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G1), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n714), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n213), .A2(new_n291), .ZN(new_n768));
  INV_X1    g0568(.A(G355), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(new_n769), .B1(G116), .B2(new_n213), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n250), .A2(G45), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n713), .A2(new_n291), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n229), .B2(new_n490), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n770), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n233), .B1(G20), .B2(new_n332), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n767), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n232), .A2(new_n334), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n450), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n785), .A2(new_n786), .B1(new_n789), .B2(G322), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT98), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n501), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n286), .A2(new_n450), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G179), .A2(G200), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n286), .A2(new_n450), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G329), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n540), .A2(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n792), .A2(G20), .A3(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G190), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n783), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n296), .B1(new_n798), .B2(new_n799), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n482), .A2(new_n484), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n232), .B1(new_n334), .B2(new_n787), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n797), .B(new_n803), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G326), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n784), .A2(new_n450), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT97), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n791), .B(new_n807), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n785), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT32), .ZN(new_n813));
  INV_X1    g0613(.A(G159), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n795), .A2(new_n814), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n812), .A2(new_n202), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n813), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n805), .A2(new_n223), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n801), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G77), .A2(new_n820), .B1(new_n789), .B2(G58), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n291), .B1(new_n218), .B2(new_n799), .C1(new_n793), .C2(new_n459), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G50), .B2(new_n809), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n817), .A2(new_n819), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n811), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n782), .B1(new_n825), .B2(new_n779), .ZN(new_n826));
  INV_X1    g0626(.A(new_n778), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n696), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n767), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n697), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n696), .A2(G330), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT99), .Z(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  OAI211_X1 g0634(.A(new_n397), .B(new_n398), .C1(new_n400), .C2(new_n372), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n265), .A2(new_n403), .B1(new_n835), .B2(new_n264), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT74), .B1(new_n836), .B2(new_n396), .ZN(new_n837));
  INV_X1    g0637(.A(new_n417), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n692), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n419), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n424), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT100), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n422), .A2(new_n423), .A3(new_n693), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n839), .A2(new_n419), .B1(new_n423), .B2(new_n422), .ZN(new_n845));
  INV_X1    g0645(.A(new_n843), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT100), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n721), .B(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n767), .B1(new_n849), .B2(new_n760), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n760), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n779), .A2(new_n776), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n829), .B1(new_n206), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n296), .B1(new_n799), .B2(new_n459), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n854), .B(new_n818), .C1(new_n809), .C2(G303), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n540), .B2(new_n812), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n788), .A2(new_n483), .B1(new_n802), .B2(new_n795), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n801), .A2(new_n553), .B1(new_n218), .B2(new_n793), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G159), .A2(new_n820), .B1(new_n789), .B2(G143), .ZN(new_n860));
  INV_X1    g0660(.A(G137), .ZN(new_n861));
  INV_X1    g0661(.A(new_n809), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n860), .B1(new_n812), .B2(new_n433), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT34), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n291), .B1(new_n439), .B2(new_n799), .C1(new_n805), .C2(new_n201), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n202), .A2(new_n793), .B1(new_n795), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n859), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n779), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n853), .B1(new_n869), .B2(new_n870), .C1(new_n848), .C2(new_n777), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n851), .A2(new_n871), .ZN(G384));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n343), .A2(new_n336), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  INV_X1    g0676(.A(new_n690), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n300), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n343), .A2(new_n336), .A3(new_n876), .A4(new_n878), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT104), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n343), .A2(new_n336), .A3(new_n878), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n879), .A2(new_n881), .B1(KEYINPUT37), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n878), .B1(new_n659), .B2(new_n666), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n873), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n232), .A2(new_n296), .A3(new_n281), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n886), .B(G68), .C1(new_n281), .C2(new_n280), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT16), .B1(new_n887), .B2(new_n277), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n270), .B1(new_n294), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n877), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n348), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n880), .B(new_n875), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n889), .B1(new_n333), .B2(new_n335), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n343), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n891), .B1(new_n895), .B2(KEYINPUT103), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT103), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n343), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n876), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT38), .B(new_n892), .C1(new_n893), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n379), .A2(new_n370), .A3(new_n383), .A4(new_n358), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n385), .A2(new_n692), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n663), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n903), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n384), .B2(new_n391), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT102), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT102), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n392), .A2(new_n908), .A3(new_n903), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n848), .A3(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n508), .A2(new_n512), .A3(new_n517), .ZN(new_n911));
  INV_X1    g0711(.A(new_n654), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n611), .B1(new_n912), .B2(new_n655), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n911), .A2(new_n574), .A3(new_n913), .A4(new_n693), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT31), .B1(new_n751), .B2(new_n692), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n910), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n901), .A2(new_n918), .A3(KEYINPUT40), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT105), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n885), .B2(new_n900), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT105), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n918), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n895), .A2(KEYINPUT103), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n898), .A3(new_n890), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .B1(new_n879), .B2(new_n881), .ZN(new_n928));
  INV_X1    g0728(.A(new_n892), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n873), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n900), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n918), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n921), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n914), .A2(new_n917), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n671), .ZN(new_n936));
  OAI21_X1  g0736(.A(G330), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n934), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n901), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n391), .A2(new_n385), .A3(new_n693), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n930), .A2(KEYINPUT39), .A3(new_n900), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n846), .B1(new_n721), .B2(new_n848), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n907), .A2(new_n909), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n931), .A3(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n944), .B(new_n949), .C1(new_n666), .C2(new_n877), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n722), .A2(new_n671), .A3(new_n734), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n670), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n950), .B(new_n952), .Z(new_n953));
  OAI22_X1  g0753(.A1(new_n938), .A2(new_n953), .B1(new_n209), .B2(new_n764), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n938), .ZN(new_n955));
  INV_X1    g0755(.A(new_n624), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT35), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT35), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n957), .A2(new_n958), .A3(G116), .A4(new_n234), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT36), .Z(new_n960));
  NAND4_X1  g0760(.A1(new_n229), .A2(G77), .A3(new_n274), .A4(new_n272), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n202), .A2(G50), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT101), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n209), .B(G13), .C1(new_n961), .C2(new_n963), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n955), .A2(new_n960), .A3(new_n964), .ZN(G367));
  OR2_X1    g0765(.A1(new_n793), .A2(new_n206), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n861), .B2(new_n795), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n291), .B1(new_n201), .B2(new_n799), .C1(new_n801), .C2(new_n439), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(G159), .C2(new_n785), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n806), .A2(G68), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n433), .B2(new_n788), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT111), .ZN(new_n972));
  INV_X1    g0772(.A(G143), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n969), .B(new_n972), .C1(new_n973), .C2(new_n810), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n810), .A2(new_n802), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n540), .A2(new_n801), .B1(new_n788), .B2(new_n798), .ZN(new_n976));
  INV_X1    g0776(.A(new_n795), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n976), .B1(G317), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n785), .A2(new_n804), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n805), .A2(new_n459), .B1(new_n793), .B2(new_n223), .ZN(new_n980));
  INV_X1    g0780(.A(new_n799), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n981), .A2(KEYINPUT46), .A3(G116), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT46), .B1(new_n981), .B2(G116), .ZN(new_n983));
  NOR4_X1   g0783(.A1(new_n980), .A2(new_n982), .A3(new_n983), .A4(new_n291), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n978), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n974), .B1(new_n975), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n779), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n606), .A2(new_n693), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n612), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n603), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(new_n778), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n772), .A2(new_n244), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n781), .B1(new_n713), .B2(new_n576), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n829), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n988), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT110), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n990), .A2(new_n991), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT43), .Z(new_n999));
  OAI211_X1 g0799(.A(new_n649), .B(new_n653), .C1(new_n650), .C2(new_n693), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n680), .A2(new_n692), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n702), .A2(new_n710), .A3(new_n1002), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n512), .A2(new_n517), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n649), .B1(new_n1004), .B2(new_n1000), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1003), .A2(KEYINPUT42), .B1(new_n693), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT106), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n700), .A2(new_n701), .B1(new_n706), .B2(new_n709), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT42), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n1009), .A3(new_n1002), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1007), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1012));
  OAI211_X1 g0812(.A(KEYINPUT107), .B(new_n999), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT106), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT107), .B1(new_n1020), .B2(new_n999), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1002), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1019), .A2(new_n1021), .B1(new_n703), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n999), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT107), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n703), .A2(new_n1022), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1026), .A2(new_n1027), .A3(new_n1018), .A4(new_n1013), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n711), .A2(new_n1002), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n711), .A2(KEYINPUT45), .A3(new_n1002), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n711), .B2(new_n1002), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1022), .B1(KEYINPUT108), .B2(KEYINPUT44), .C1(new_n1008), .C2(new_n704), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n703), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n702), .A2(new_n710), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(new_n697), .A3(KEYINPUT109), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n697), .B1(KEYINPUT109), .B2(new_n1044), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1046), .A2(new_n1047), .B1(new_n702), .B2(new_n710), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1047), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n702), .A2(new_n710), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n1050), .A3(new_n1045), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n761), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1035), .A2(new_n1040), .A3(new_n703), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1043), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n762), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n714), .B(KEYINPUT41), .Z(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n766), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n997), .B1(new_n1030), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n766), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1062), .A2(new_n1029), .A3(KEYINPUT110), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n996), .B1(new_n1061), .B2(new_n1063), .ZN(G387));
  NAND3_X1  g0864(.A1(new_n700), .A2(new_n701), .A3(new_n778), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n768), .A2(new_n716), .B1(G107), .B2(new_n213), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n241), .A2(new_n490), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n716), .ZN(new_n1068));
  AOI211_X1 g0868(.A(G45), .B(new_n1068), .C1(G68), .C2(G77), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n268), .A2(G50), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT50), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n773), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1066), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n767), .B1(new_n1073), .B2(new_n781), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n805), .A2(new_n400), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n801), .A2(new_n202), .B1(new_n433), .B2(new_n795), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(G50), .C2(new_n789), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n291), .B1(new_n206), .B2(new_n799), .C1(new_n793), .C2(new_n223), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n268), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n785), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1077), .B(new_n1080), .C1(new_n814), .C2(new_n862), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n291), .B1(new_n977), .B2(G326), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G303), .A2(new_n820), .B1(new_n789), .B2(G317), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT112), .Z(new_n1084));
  INV_X1    g0884(.A(G322), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1084), .B1(new_n802), .B2(new_n812), .C1(new_n810), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n806), .A2(G283), .B1(new_n981), .B2(new_n804), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT49), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1082), .B1(new_n553), .B2(new_n793), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1081), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1074), .B1(new_n1095), .B2(new_n779), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1065), .A2(new_n1096), .B1(new_n1097), .B2(new_n766), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n762), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n714), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1097), .A2(new_n762), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(G393));
  NAND3_X1  g0902(.A1(new_n1043), .A2(new_n766), .A3(new_n1053), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n780), .B1(new_n223), .B2(new_n213), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n772), .B2(new_n253), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n809), .A2(G150), .B1(new_n789), .B2(G159), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT51), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n805), .A2(new_n206), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n1079), .B2(new_n820), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n973), .B2(new_n795), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n296), .B1(new_n981), .B2(G68), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n218), .B2(new_n793), .C1(new_n812), .C2(new_n439), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1107), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(KEYINPUT113), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n809), .A2(G317), .B1(new_n789), .B2(G311), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT52), .Z(new_n1117));
  OAI22_X1  g0917(.A1(new_n805), .A2(new_n553), .B1(new_n795), .B2(new_n1085), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G294), .B2(new_n820), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n296), .B1(new_n540), .B2(new_n799), .C1(new_n793), .C2(new_n459), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G303), .B2(new_n785), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1114), .A2(KEYINPUT113), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1115), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n829), .B(new_n1105), .C1(new_n1124), .C2(new_n779), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n827), .B2(new_n1002), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1103), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1053), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n703), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1099), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(new_n714), .A3(new_n1054), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT114), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT114), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1130), .A2(new_n1133), .A3(new_n714), .A4(new_n1054), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1127), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(G390));
  OAI21_X1  g0936(.A(new_n941), .B1(new_n945), .B2(new_n947), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n943), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT39), .B1(new_n885), .B2(new_n900), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n693), .B(new_n848), .C1(new_n729), .C2(new_n733), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n843), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n948), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n941), .A3(new_n901), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n907), .A2(new_n848), .A3(new_n909), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n754), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(G330), .C1(new_n736), .C2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT116), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n918), .A2(KEYINPUT116), .A3(G330), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT115), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(G330), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n848), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n752), .A2(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1153), .B(new_n1154), .C1(new_n914), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n948), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1140), .B(new_n1144), .C1(new_n1152), .C2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT115), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n946), .A2(new_n948), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1161), .A2(new_n941), .B1(new_n940), .B2(new_n943), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n901), .A2(new_n941), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n948), .B2(new_n1142), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1160), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1158), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT117), .ZN(new_n1167));
  OAI211_X1 g0967(.A(G330), .B(new_n848), .C1(new_n736), .C2(new_n759), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n947), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1150), .A2(new_n1169), .A3(new_n1151), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n946), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1142), .B1(new_n1156), .B2(new_n948), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n935), .A2(G330), .A3(new_n848), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n947), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n935), .A2(G330), .A3(new_n671), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n670), .A2(new_n951), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1167), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1170), .A2(new_n946), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1181), .A2(KEYINPUT117), .A3(new_n1178), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1166), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1176), .A2(new_n1167), .A3(new_n1179), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT117), .B1(new_n1181), .B2(new_n1178), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1158), .A2(new_n1165), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1183), .A2(new_n714), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n776), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n788), .A2(new_n553), .B1(new_n483), .B2(new_n795), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1108), .B(new_n1190), .C1(G97), .C2(new_n820), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n296), .B1(new_n218), .B2(new_n799), .C1(new_n793), .C2(new_n202), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G107), .B2(new_n785), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(new_n540), .C2(new_n862), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n981), .A2(G150), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT53), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT54), .B(G143), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1196), .B1(new_n820), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n806), .A2(G159), .ZN(new_n1200));
  INV_X1    g1000(.A(G125), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n439), .A2(new_n793), .B1(new_n795), .B2(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n296), .B(new_n1202), .C1(G132), .C2(new_n789), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G128), .A2(new_n809), .B1(new_n785), .B2(G137), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n870), .B1(new_n1194), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n829), .B(new_n1206), .C1(new_n268), .C2(new_n852), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1166), .A2(new_n766), .B1(new_n1189), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1188), .A2(new_n1208), .ZN(G378));
  NOR2_X1   g1009(.A1(new_n793), .A2(new_n201), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G283), .B2(new_n977), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n785), .A2(G97), .ZN(new_n1212));
  INV_X1    g1012(.A(G41), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n296), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n981), .B2(G77), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n970), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G116), .B2(new_n809), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n820), .A2(new_n576), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n789), .A2(G107), .ZN(new_n1219));
  AND4_X1   g1019(.A1(new_n1211), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1220), .A2(KEYINPUT58), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(KEYINPUT58), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1214), .B(new_n439), .C1(G33), .C2(G41), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n806), .A2(G150), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n981), .A2(new_n1198), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(G128), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1227), .B1(new_n788), .B2(new_n1228), .C1(new_n861), .C2(new_n801), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1201), .A2(new_n862), .B1(new_n812), .B2(new_n866), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n288), .B(new_n1213), .C1(new_n793), .C2(new_n814), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G124), .B2(new_n977), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n870), .B1(new_n1224), .B2(new_n1237), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n829), .B(new_n1238), .C1(new_n439), .C2(new_n852), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n443), .A2(new_n877), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n455), .A2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n444), .B(new_n1240), .C1(new_n453), .C2(new_n454), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT118), .ZN(new_n1245));
  XOR2_X1   g1045(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1246));
  INV_X1    g1046(.A(KEYINPUT118), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1242), .A2(new_n1247), .A3(new_n1243), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1246), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1239), .B1(new_n1251), .B2(new_n777), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n922), .A2(new_n923), .A3(new_n918), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n923), .B1(new_n922), .B2(new_n918), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n933), .B(G330), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1251), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT119), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n950), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n925), .A2(new_n1251), .A3(G330), .A4(new_n933), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1259), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1252), .B1(new_n1263), .B2(new_n1059), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1257), .A2(new_n950), .A3(new_n1260), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n950), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT57), .ZN(new_n1268));
  OR3_X1    g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1178), .B1(new_n1270), .B2(new_n1166), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n714), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1183), .A2(new_n1179), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT57), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1265), .B1(new_n1272), .B2(new_n1275), .ZN(G375));
  AOI21_X1  g1076(.A(new_n829), .B1(new_n202), .B2(new_n852), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n291), .B1(new_n799), .B2(new_n814), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1210), .B(new_n1278), .C1(new_n809), .C2(G132), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n812), .B2(new_n1197), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n805), .A2(new_n439), .B1(new_n795), .B2(new_n1228), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n861), .A2(new_n788), .B1(new_n801), .B2(new_n433), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n291), .B1(new_n981), .B2(G97), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n966), .B(new_n1284), .C1(new_n862), .C2(new_n483), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1075), .B1(G303), .B2(new_n977), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n1286), .B1(new_n459), .B2(new_n801), .C1(new_n540), .C2(new_n788), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1285), .B(new_n1287), .C1(G116), .C2(new_n785), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1288), .A2(KEYINPUT120), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(KEYINPUT120), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1283), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1291), .A2(KEYINPUT121), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n779), .B1(new_n1291), .B2(KEYINPUT121), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n1277), .B1(new_n777), .B2(new_n948), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1181), .B2(new_n1059), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1171), .A2(new_n1178), .A3(new_n1175), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1184), .A2(new_n1185), .A3(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1298), .B2(new_n1056), .ZN(G381));
  INV_X1    g1099(.A(new_n996), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1030), .A2(new_n1060), .A3(new_n997), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT110), .B1(new_n1062), .B2(new_n1029), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1300), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(G393), .A2(G396), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1305), .A2(G381), .A3(G384), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1303), .A2(new_n1135), .A3(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT122), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT122), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n715), .B1(new_n1273), .B2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1268), .B1(new_n1271), .B2(new_n1263), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1264), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(G378), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1309), .A2(new_n1311), .A3(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(KEYINPUT123), .ZN(G407));
  INV_X1    g1120(.A(G213), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1318), .B2(new_n691), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1319), .A2(KEYINPUT123), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT123), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1317), .B1(new_n1308), .B2(KEYINPUT122), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1325), .B2(new_n1311), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1322), .B1(new_n1323), .B2(new_n1326), .ZN(G409));
  OR2_X1    g1127(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1298), .A2(KEYINPUT60), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT60), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1297), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n714), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1296), .B(new_n1328), .C1(new_n1329), .C2(new_n1332), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(G384), .B(KEYINPUT124), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1332), .B1(new_n1298), .B2(KEYINPUT60), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1334), .B1(new_n1335), .B2(new_n1295), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n691), .A2(G213), .A3(G2897), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1333), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1333), .B2(new_n1336), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n691), .A2(G213), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1273), .A2(new_n1274), .A3(new_n1057), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1252), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1343), .B1(new_n1344), .B2(new_n766), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1342), .A2(new_n1188), .A3(new_n1208), .A4(new_n1345), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1341), .B(new_n1346), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1347));
  AOI21_X1  g1147(.A(KEYINPUT61), .B1(new_n1340), .B2(new_n1347), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1333), .A2(new_n1336), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1349), .ZN(new_n1350));
  OAI21_X1  g1150(.A(KEYINPUT62), .B1(new_n1347), .B2(new_n1350), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1346), .A2(new_n1341), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G375), .A2(G378), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT62), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1352), .A2(new_n1353), .A3(new_n1354), .A4(new_n1349), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1348), .A2(new_n1351), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G393), .A2(G396), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  NOR3_X1   g1158(.A1(new_n1358), .A2(new_n1304), .A3(KEYINPUT125), .ZN(new_n1359));
  OAI211_X1 g1159(.A(new_n996), .B(new_n1135), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1360));
  OAI21_X1  g1160(.A(KEYINPUT125), .B1(new_n1358), .B2(new_n1304), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1135), .B1(new_n1363), .B2(new_n996), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1359), .B1(new_n1362), .B2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1361), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1366), .B1(new_n1303), .B2(new_n1135), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(G387), .A2(G390), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1359), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1367), .A2(new_n1368), .A3(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1365), .A2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1356), .A2(new_n1371), .ZN(new_n1372));
  NOR3_X1   g1172(.A1(new_n1362), .A2(new_n1359), .A3(new_n1364), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1369), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT63), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1376), .B1(new_n1347), .B2(new_n1350), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1352), .A2(new_n1353), .A3(KEYINPUT63), .A4(new_n1349), .ZN(new_n1378));
  NAND4_X1  g1178(.A1(new_n1375), .A2(new_n1348), .A3(new_n1377), .A4(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1372), .A2(new_n1379), .ZN(G405));
  NAND2_X1  g1180(.A1(new_n1349), .A2(KEYINPUT126), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1381), .A2(new_n1353), .A3(new_n1317), .ZN(new_n1382));
  INV_X1    g1182(.A(new_n1382), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1381), .B1(new_n1317), .B2(new_n1353), .ZN(new_n1384));
  OAI21_X1  g1184(.A(new_n1371), .B1(new_n1383), .B2(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1353), .A2(new_n1317), .ZN(new_n1386));
  AND2_X1   g1186(.A1(new_n1349), .A2(KEYINPUT126), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1386), .A2(new_n1387), .ZN(new_n1388));
  NAND4_X1  g1188(.A1(new_n1388), .A2(new_n1365), .A3(new_n1370), .A4(new_n1382), .ZN(new_n1389));
  AND2_X1   g1189(.A1(new_n1385), .A2(new_n1389), .ZN(G402));
endmodule


