//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n462), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT70), .B1(new_n462), .B2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(G137), .A3(new_n475), .ZN(new_n476));
  OAI22_X1  g051(.A1(new_n465), .A2(new_n466), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G125), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n474), .A2(new_n475), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n470), .A2(G2104), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(new_n472), .A3(G125), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n479), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n474), .A2(new_n475), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(KEYINPUT68), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n477), .B1(new_n484), .B2(new_n489), .ZN(G160));
  OAI221_X1 g065(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n483), .C2(G112), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n473), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n473), .A2(new_n483), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G124), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n491), .B(new_n493), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n462), .A2(G114), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n507), .A2(new_n502), .A3(KEYINPUT71), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n500), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n474), .A2(G138), .A3(new_n475), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT4), .B1(new_n473), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n483), .A2(new_n481), .A3(new_n512), .A4(G138), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(G164));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n515), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n524), .A2(new_n525), .B1(new_n523), .B2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(new_n519), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G88), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(G62), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n517), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(KEYINPUT73), .B1(new_n530), .B2(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G166));
  AND2_X1   g113(.A1(new_n526), .A2(new_n527), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n520), .A2(G51), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n540), .A2(new_n545), .ZN(G168));
  AOI22_X1  g121(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n517), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n520), .A2(G52), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n528), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(G171));
  AOI22_X1  g127(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n517), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n527), .A2(G543), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT74), .B(G43), .Z(new_n557));
  OAI22_X1  g132(.A1(new_n528), .A2(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n520), .A2(new_n566), .A3(G53), .ZN(new_n567));
  AND2_X1   g142(.A1(KEYINPUT6), .A2(G651), .ZN(new_n568));
  NOR2_X1   g143(.A1(KEYINPUT6), .A2(G651), .ZN(new_n569));
  OAI211_X1 g144(.A(G53), .B(G543), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n526), .A2(G91), .A3(new_n527), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n526), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n572), .B(new_n573), .C1(new_n574), .C2(new_n517), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n539), .A2(G87), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  INV_X1    g155(.A(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n556), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n520), .A2(KEYINPUT76), .A3(G49), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n579), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n523), .A2(G543), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n515), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n589));
  AOI21_X1  g164(.A(KEYINPUT72), .B1(new_n515), .B2(KEYINPUT5), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(KEYINPUT77), .A3(G651), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n539), .A2(G86), .B1(G48), .B2(new_n520), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G305));
  XNOR2_X1  g174(.A(KEYINPUT78), .B(G85), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n539), .A2(new_n600), .B1(G47), .B2(new_n520), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n517), .B2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n528), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n605), .A2(new_n608), .B1(G54), .B2(new_n520), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  INV_X1    g185(.A(G79), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n591), .A2(new_n610), .B1(new_n611), .B2(new_n515), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI221_X1 g189(.A(KEYINPUT79), .B1(new_n611), .B2(new_n515), .C1(new_n591), .C2(new_n610), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n614), .A2(G651), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n604), .B1(new_n618), .B2(G868), .ZN(G321));
  XNOR2_X1  g194(.A(G321), .B(KEYINPUT80), .ZN(G284));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  INV_X1    g196(.A(G299), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(G868), .B2(new_n622), .ZN(G280));
  XOR2_X1   g198(.A(G280), .B(KEYINPUT81), .Z(G297));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n618), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g205(.A(new_n464), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n462), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(new_n481), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT82), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n494), .A2(G123), .ZN(new_n640));
  OAI221_X1 g215(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n483), .C2(G111), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n492), .A2(G135), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT83), .Z(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n645), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n665), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n636), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n668), .B2(new_n664), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(G2096), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n683), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n685), .B(new_n688), .C1(new_n680), .C2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT88), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  MUX2_X1   g272(.A(G23), .B(G288), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT89), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT33), .B(G1976), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G16), .A2(G22), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G166), .B2(G16), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G6), .B(G305), .S(G16), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n701), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT34), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  MUX2_X1   g287(.A(G24), .B(G290), .S(G16), .Z(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(G1986), .Z(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G25), .ZN(new_n716));
  OAI221_X1 g291(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n483), .C2(G107), .ZN(new_n717));
  INV_X1    g292(.A(G119), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n495), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G131), .B2(new_n492), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n716), .B1(new_n720), .B2(new_n715), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n711), .A2(new_n712), .A3(new_n714), .A4(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G20), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n727), .B(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n622), .B2(new_n728), .ZN(new_n731));
  INV_X1    g306(.A(G1956), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G4), .A2(G16), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n618), .B2(G16), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT90), .B(G1348), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n481), .A2(G127), .ZN(new_n738));
  INV_X1    g313(.A(G115), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n468), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n740), .A2(new_n488), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT92), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT25), .ZN(new_n743));
  NAND2_X1  g318(.A1(G103), .A2(G2104), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n488), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n483), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n745), .A2(new_n746), .B1(new_n492), .B2(G139), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n740), .A2(KEYINPUT92), .A3(new_n488), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n742), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G33), .B(new_n749), .S(G29), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n733), .B(new_n737), .C1(new_n751), .C2(G2072), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n728), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n728), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(G1966), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT96), .Z(new_n756));
  AND2_X1   g331(.A1(new_n715), .A2(G32), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n492), .A2(G141), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT94), .Z(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  INV_X1    g336(.A(G105), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n465), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G129), .B2(new_n494), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n757), .B1(new_n765), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n715), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT91), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT28), .ZN(new_n772));
  OAI221_X1 g347(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n483), .C2(G116), .ZN(new_n773));
  INV_X1    g348(.A(G128), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n495), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G140), .B2(new_n492), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n772), .B1(new_n776), .B2(new_n715), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n756), .A2(new_n768), .A3(new_n769), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G171), .A2(new_n728), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G5), .B2(new_n728), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT24), .ZN(new_n785));
  INV_X1    g360(.A(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G160), .B2(new_n715), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n784), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G19), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n559), .B2(G16), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n644), .A2(new_n715), .B1(G1341), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(G1341), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n782), .B2(new_n783), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n754), .A2(G1966), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n790), .A2(new_n791), .ZN(new_n799));
  INV_X1    g374(.A(G28), .ZN(new_n800));
  OR3_X1    g375(.A1(new_n800), .A2(KEYINPUT95), .A3(KEYINPUT30), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT95), .B1(new_n800), .B2(KEYINPUT30), .ZN(new_n802));
  AOI21_X1  g377(.A(G29), .B1(new_n800), .B2(KEYINPUT30), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT31), .B(G11), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n798), .A2(new_n799), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n792), .A2(new_n795), .A3(new_n797), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n751), .A2(G2072), .ZN(new_n808));
  NOR2_X1   g383(.A1(G27), .A2(G29), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G164), .B2(G29), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n715), .A2(G35), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n715), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT29), .B(G2090), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n814), .B(new_n815), .Z(new_n816));
  NAND4_X1  g391(.A1(new_n807), .A2(new_n808), .A3(new_n812), .A4(new_n816), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n726), .A2(new_n752), .A3(new_n780), .A4(new_n817), .ZN(G311));
  OR4_X1    g393(.A1(new_n726), .A2(new_n752), .A3(new_n780), .A4(new_n817), .ZN(G150));
  NAND2_X1  g394(.A1(new_n618), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n517), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n520), .A2(G55), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n528), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n559), .A2(new_n827), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n554), .A2(new_n558), .B1(new_n823), .B2(new_n826), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n821), .B(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  INV_X1    g407(.A(G860), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n827), .A2(new_n833), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(G145));
  OR2_X1    g413(.A1(new_n749), .A2(KEYINPUT99), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n839), .A2(KEYINPUT100), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n749), .A2(KEYINPUT100), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n511), .A2(new_n513), .ZN(new_n843));
  INV_X1    g418(.A(new_n473), .ZN(new_n844));
  OAI21_X1  g419(.A(KEYINPUT71), .B1(new_n507), .B2(new_n502), .ZN(new_n845));
  OR2_X1    g420(.A1(G102), .A2(G2105), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n846), .A2(new_n505), .A3(new_n501), .A4(G2104), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n844), .A2(new_n499), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n765), .B(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n776), .B(KEYINPUT98), .Z(new_n851));
  AND2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n850), .A2(new_n851), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n851), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n840), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n494), .A2(G130), .ZN(new_n858));
  OAI221_X1 g433(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n483), .C2(G118), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n492), .A2(G142), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n635), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n720), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n854), .A2(new_n857), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n644), .B(new_n497), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G160), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n863), .B1(new_n854), .B2(new_n857), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(G37), .ZN(new_n870));
  INV_X1    g445(.A(new_n864), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n854), .A2(new_n857), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT101), .B1(new_n872), .B2(new_n863), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n871), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n870), .B1(new_n876), .B2(new_n866), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n868), .A2(new_n874), .ZN(new_n880));
  AOI211_X1 g455(.A(KEYINPUT101), .B(new_n863), .C1(new_n854), .C2(new_n857), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n864), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n866), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(KEYINPUT102), .A3(new_n870), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n879), .A2(KEYINPUT40), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT40), .B1(new_n879), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(G395));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n827), .B2(G868), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  XNOR2_X1  g466(.A(G166), .B(G290), .ZN(new_n892));
  XNOR2_X1  g467(.A(G305), .B(G288), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n892), .B(new_n893), .Z(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n894), .B2(KEYINPUT105), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n894), .B2(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(new_n895), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n617), .A2(new_n622), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n617), .A2(new_n622), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(KEYINPUT103), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n900), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n901), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n627), .B(new_n830), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n907), .A2(new_n901), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n899), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n899), .A2(new_n913), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(G868), .A3(new_n915), .ZN(new_n916));
  MUX2_X1   g491(.A(new_n889), .B(new_n890), .S(new_n916), .Z(G295));
  MUX2_X1   g492(.A(new_n889), .B(new_n890), .S(new_n916), .Z(G331));
  NAND2_X1  g493(.A1(new_n828), .A2(new_n829), .ZN(new_n919));
  NOR2_X1   g494(.A1(G301), .A2(KEYINPUT107), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G168), .B1(G301), .B2(KEYINPUT107), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n920), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n923), .ZN(new_n926));
  INV_X1    g501(.A(new_n924), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(new_n927), .B2(new_n921), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n906), .A3(new_n908), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(new_n928), .A3(new_n912), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n894), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  AOI21_X1  g509(.A(G37), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n894), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(new_n936), .A3(new_n931), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(KEYINPUT108), .A3(new_n894), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n905), .B1(new_n925), .B2(new_n928), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n894), .B1(new_n904), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n912), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n943), .B1(new_n944), .B2(new_n942), .ZN(new_n945));
  AND4_X1   g520(.A1(KEYINPUT43), .A2(new_n935), .A3(new_n938), .A4(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT44), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n935), .A2(new_n940), .A3(new_n938), .A4(new_n945), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n948), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n947), .B1(new_n953), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g529(.A(KEYINPUT121), .ZN(new_n955));
  INV_X1    g530(.A(G1966), .ZN(new_n956));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT45), .ZN(new_n958));
  OAI211_X1 g533(.A(G40), .B(G160), .C1(G164), .C2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT45), .B1(new_n849), .B2(new_n957), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT113), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n849), .A2(new_n957), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT50), .ZN(new_n964));
  INV_X1    g539(.A(new_n476), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n844), .A2(new_n965), .B1(new_n633), .B2(G101), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n482), .A2(new_n478), .A3(new_n483), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT68), .B1(new_n487), .B2(new_n488), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n966), .B(G40), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n843), .B2(new_n848), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n964), .A2(new_n970), .A3(new_n791), .A4(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n975), .B(new_n956), .C1(new_n959), .C2(new_n960), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n962), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT111), .B(G8), .ZN(new_n978));
  NOR2_X1   g553(.A1(G168), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n981));
  INV_X1    g556(.A(new_n979), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n976), .A2(new_n974), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n958), .B1(new_n843), .B2(new_n848), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n969), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(G164), .B2(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n975), .B1(new_n988), .B2(new_n956), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n981), .B(new_n982), .C1(new_n990), .C2(new_n978), .ZN(new_n991));
  OAI21_X1  g566(.A(G8), .B1(new_n983), .B2(new_n989), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n981), .B1(new_n992), .B2(new_n982), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT120), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n979), .B1(new_n977), .B2(G8), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n996), .A2(KEYINPUT120), .A3(new_n981), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n955), .B(new_n980), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT120), .B1(new_n996), .B2(new_n981), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n992), .A2(new_n982), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(new_n994), .A3(KEYINPUT51), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1002), .A3(new_n991), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n955), .B1(new_n1003), .B2(new_n980), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT62), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n980), .B1(new_n995), .B2(new_n997), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT121), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT62), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n998), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n969), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n1010));
  INV_X1    g585(.A(G2090), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n973), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT110), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n988), .A2(new_n704), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1010), .A2(new_n1015), .A3(new_n1011), .A4(new_n973), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n536), .A2(G8), .A3(new_n537), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1020), .A3(G8), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n970), .A2(new_n971), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n978), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n579), .A2(new_n584), .A3(G1976), .A4(new_n585), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1025), .B(new_n1026), .C1(new_n963), .C2(new_n969), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G305), .A2(G1981), .ZN(new_n1032));
  INV_X1    g607(.A(G1981), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n596), .A2(new_n1033), .A3(new_n597), .A4(new_n598), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1031), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(KEYINPUT49), .A3(new_n1034), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1030), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1018), .B(KEYINPUT55), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1014), .A2(new_n1012), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n978), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1021), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1021), .A2(new_n1042), .A3(KEYINPUT124), .A4(new_n1039), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(G40), .B(G160), .C1(new_n971), .C2(new_n972), .ZN(new_n1048));
  INV_X1    g623(.A(new_n973), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n783), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n959), .A2(new_n960), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT122), .B1(new_n1051), .B2(new_n811), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n985), .A2(new_n987), .A3(KEYINPUT122), .A4(new_n811), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT53), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT123), .B(new_n1050), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n988), .B2(G2078), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n988), .B2(G2078), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n1053), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT123), .B1(new_n1061), .B2(new_n1050), .ZN(new_n1062));
  OAI21_X1  g637(.A(G171), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1047), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1005), .A2(new_n1009), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT63), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n977), .A2(G168), .A3(new_n1025), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1043), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1066), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1017), .A2(G8), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1040), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1071), .A3(new_n1021), .A4(new_n1039), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1034), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G288), .A2(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1039), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1077), .A2(new_n1031), .B1(new_n1078), .B2(new_n1021), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1073), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(G301), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n811), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n1086), .B(new_n477), .C1(new_n488), .C2(new_n487), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n987), .B(new_n1087), .C1(G164), .C2(new_n958), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1057), .A2(new_n1050), .A3(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1089), .A2(KEYINPUT125), .ZN(new_n1090));
  AOI21_X1  g665(.A(G301), .B1(new_n1089), .B2(KEYINPUT125), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1085), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1089), .A2(G171), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(KEYINPUT54), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1084), .A2(new_n1092), .B1(new_n1063), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n572), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(G65), .B(new_n588), .C1(new_n589), .C2(new_n590), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G78), .A2(G543), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G651), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n567), .A2(new_n571), .A3(KEYINPUT114), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1097), .A2(new_n1101), .A3(new_n573), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT115), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g684(.A1(G91), .A2(new_n539), .B1(new_n1100), .B2(G651), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1110), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n572), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(G299), .B2(new_n1104), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1956), .B1(new_n1010), .B2(new_n973), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1116), .B(G2072), .Z(new_n1117));
  AND3_X1   g692(.A1(new_n985), .A2(new_n987), .A3(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1109), .B(new_n1114), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1103), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1107), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1114), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n732), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n985), .A2(new_n987), .A3(new_n1117), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1348), .B1(new_n1010), .B2(new_n973), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n970), .A2(new_n778), .A3(new_n971), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n618), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1119), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1119), .A2(new_n1125), .A3(KEYINPUT61), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT61), .B1(new_n1119), .B2(new_n1125), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1049), .A2(new_n1048), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n617), .B(new_n1128), .C1(new_n1135), .C2(G1348), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1132), .A2(new_n1133), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT58), .B(G1341), .Z(new_n1140));
  NAND3_X1  g715(.A1(new_n1022), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n963), .B2(new_n969), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT118), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1141), .B(new_n1143), .C1(G1996), .C2(new_n988), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1145));
  AND3_X1   g720(.A1(new_n1144), .A2(new_n559), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1144), .B2(new_n559), .ZN(new_n1147));
  NOR4_X1   g722(.A1(new_n1127), .A2(new_n1129), .A3(KEYINPUT60), .A4(new_n617), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1131), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1095), .A2(new_n1150), .A3(new_n1047), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1007), .A2(new_n998), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1083), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1065), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n987), .A2(new_n969), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n765), .B(G1996), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n776), .B(G2067), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n720), .A2(new_n722), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n720), .A2(new_n722), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(G290), .B(G1986), .Z(new_n1165));
  AOI21_X1  g740(.A(new_n1156), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1154), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1156), .A2(G1996), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT46), .Z(new_n1170));
  OAI21_X1  g745(.A(new_n1155), .B1(new_n1159), .B2(new_n765), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT47), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1164), .A2(new_n1156), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1156), .A2(G1986), .A3(G290), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT48), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1161), .B(KEYINPUT126), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1160), .A2(new_n1178), .B1(new_n778), .B2(new_n776), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1175), .A2(new_n1177), .B1(new_n1156), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1174), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1168), .A2(KEYINPUT127), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1166), .B1(new_n1065), .B2(new_n1153), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1181), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1182), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g762(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1189));
  AND3_X1   g763(.A1(new_n884), .A2(KEYINPUT102), .A3(new_n870), .ZN(new_n1190));
  AOI21_X1  g764(.A(KEYINPUT102), .B1(new_n884), .B2(new_n870), .ZN(new_n1191));
  OAI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g766(.A1(new_n953), .A2(new_n1192), .ZN(G308));
  OAI221_X1 g767(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .C1(new_n951), .C2(new_n952), .ZN(G225));
endmodule


