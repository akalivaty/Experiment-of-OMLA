

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G2104), .A2(n527), .ZN(n879) );
  XNOR2_X1 U554 ( .A(n529), .B(KEYINPUT64), .ZN(n718) );
  NOR2_X1 U555 ( .A1(n633), .A2(n922), .ZN(n644) );
  NAND2_X1 U556 ( .A1(G8), .A2(n669), .ZN(n708) );
  XOR2_X1 U557 ( .A(n536), .B(KEYINPUT66), .Z(n518) );
  NOR2_X2 U558 ( .A1(G164), .A2(G1384), .ZN(n732) );
  NOR2_X2 U559 ( .A1(n528), .A2(G2105), .ZN(n529) );
  BUF_X1 U560 ( .A(n878), .Z(n519) );
  NOR2_X1 U561 ( .A1(n528), .A2(n527), .ZN(n878) );
  XNOR2_X1 U562 ( .A(n622), .B(KEYINPUT94), .ZN(n633) );
  NOR2_X1 U563 ( .A1(n669), .A2(n970), .ZN(n619) );
  BUF_X1 U564 ( .A(n718), .Z(n719) );
  BUF_X1 U565 ( .A(n713), .Z(n714) );
  INV_X1 U566 ( .A(KEYINPUT97), .ZN(n605) );
  NOR2_X1 U567 ( .A1(G168), .A2(n609), .ZN(n611) );
  AND2_X1 U568 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U569 ( .A1(n537), .A2(n518), .ZN(n520) );
  NOR2_X1 U570 ( .A1(n708), .A2(n688), .ZN(n521) );
  INV_X1 U571 ( .A(KEYINPUT31), .ZN(n615) );
  INV_X1 U572 ( .A(n930), .ZN(n691) );
  NOR2_X1 U573 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U574 ( .A1(G543), .A2(G651), .ZN(n795) );
  INV_X1 U575 ( .A(G2104), .ZN(n528) );
  INV_X1 U576 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n519), .A2(G114), .ZN(n526) );
  XNOR2_X1 U578 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n523) );
  NOR2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X1 U580 ( .A(n523), .B(n522), .ZN(n713) );
  NAND2_X1 U581 ( .A1(n713), .A2(G138), .ZN(n524) );
  XOR2_X1 U582 ( .A(KEYINPUT85), .B(n524), .Z(n525) );
  NAND2_X1 U583 ( .A1(n526), .A2(n525), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n879), .A2(G126), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G102), .A2(n718), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U587 ( .A1(n533), .A2(n532), .ZN(G164) );
  NAND2_X1 U588 ( .A1(G137), .A2(n713), .ZN(n535) );
  NAND2_X1 U589 ( .A1(G125), .A2(n879), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X1 U591 ( .A1(G113), .A2(n878), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n718), .A2(G101), .ZN(n538) );
  XNOR2_X1 U593 ( .A(n538), .B(KEYINPUT65), .ZN(n539) );
  XNOR2_X1 U594 ( .A(KEYINPUT23), .B(n539), .ZN(n540) );
  AND2_X2 U595 ( .A1(n520), .A2(n540), .ZN(G160) );
  INV_X1 U596 ( .A(G651), .ZN(n546) );
  NOR2_X1 U597 ( .A1(G543), .A2(n546), .ZN(n541) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n541), .Z(n791) );
  NAND2_X1 U599 ( .A1(G64), .A2(n791), .ZN(n542) );
  XNOR2_X1 U600 ( .A(n542), .B(KEYINPUT68), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT0), .B(G543), .Z(n584) );
  NOR2_X2 U602 ( .A1(n584), .A2(G651), .ZN(n792) );
  NAND2_X1 U603 ( .A1(G52), .A2(n792), .ZN(n543) );
  XOR2_X1 U604 ( .A(KEYINPUT69), .B(n543), .Z(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n551) );
  NAND2_X1 U606 ( .A1(G90), .A2(n795), .ZN(n548) );
  NOR2_X1 U607 ( .A1(n584), .A2(n546), .ZN(n796) );
  NAND2_X1 U608 ( .A1(G77), .A2(n796), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U611 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U612 ( .A1(G63), .A2(n791), .ZN(n553) );
  NAND2_X1 U613 ( .A1(G51), .A2(n792), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U615 ( .A(KEYINPUT6), .B(n554), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n795), .A2(G89), .ZN(n555) );
  XNOR2_X1 U617 ( .A(KEYINPUT4), .B(n555), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n796), .A2(G76), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT75), .B(n556), .Z(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U621 ( .A(n559), .B(KEYINPUT5), .Z(n560) );
  NOR2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT76), .B(n562), .Z(n563) );
  XNOR2_X1 U624 ( .A(KEYINPUT7), .B(n563), .ZN(G168) );
  NAND2_X1 U625 ( .A1(G91), .A2(n795), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G78), .A2(n796), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n571) );
  NAND2_X1 U628 ( .A1(n792), .A2(G53), .ZN(n566) );
  XNOR2_X1 U629 ( .A(n566), .B(KEYINPUT70), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G65), .A2(n791), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT71), .B(n569), .Z(n570) );
  NOR2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT72), .B(n572), .Z(G299) );
  NAND2_X1 U635 ( .A1(G88), .A2(n795), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT82), .B(n573), .Z(n580) );
  NAND2_X1 U637 ( .A1(G62), .A2(n791), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G50), .A2(n792), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT81), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G75), .A2(n796), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U643 ( .A1(n580), .A2(n579), .ZN(G166) );
  INV_X1 U644 ( .A(G166), .ZN(G303) );
  XOR2_X1 U645 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U646 ( .A1(G49), .A2(n792), .ZN(n582) );
  NAND2_X1 U647 ( .A1(G74), .A2(G651), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U649 ( .A1(n791), .A2(n583), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n584), .A2(G87), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U652 ( .A1(G61), .A2(n791), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G86), .A2(n795), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n796), .A2(G73), .ZN(n589) );
  XOR2_X1 U656 ( .A(KEYINPUT2), .B(n589), .Z(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n792), .A2(G48), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(G305) );
  NAND2_X1 U660 ( .A1(G85), .A2(n795), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G72), .A2(n796), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G60), .A2(n791), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G47), .A2(n792), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n597), .A2(n596), .ZN(n598) );
  OR2_X1 U666 ( .A1(n599), .A2(n598), .ZN(G290) );
  NAND2_X1 U667 ( .A1(G160), .A2(G40), .ZN(n731) );
  INV_X1 U668 ( .A(n731), .ZN(n600) );
  NAND2_X2 U669 ( .A1(n732), .A2(n600), .ZN(n669) );
  NOR2_X1 U670 ( .A1(G2084), .A2(n669), .ZN(n604) );
  NAND2_X1 U671 ( .A1(G8), .A2(n604), .ZN(n668) );
  NOR2_X1 U672 ( .A1(G1966), .A2(n708), .ZN(n666) );
  XOR2_X1 U673 ( .A(KEYINPUT25), .B(G2078), .Z(n974) );
  NOR2_X1 U674 ( .A1(n974), .A2(n669), .ZN(n602) );
  AND2_X1 U675 ( .A1(n732), .A2(n600), .ZN(n653) );
  XOR2_X1 U676 ( .A(G1961), .B(KEYINPUT91), .Z(n945) );
  NOR2_X1 U677 ( .A1(n653), .A2(n945), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U679 ( .A(KEYINPUT92), .B(n603), .Z(n617) );
  OR2_X1 U680 ( .A1(G171), .A2(n617), .ZN(n613) );
  NOR2_X1 U681 ( .A1(n666), .A2(n604), .ZN(n606) );
  XNOR2_X1 U682 ( .A(n606), .B(n605), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n607), .A2(G8), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n608), .B(KEYINPUT30), .ZN(n609) );
  INV_X1 U685 ( .A(KEYINPUT98), .ZN(n610) );
  XNOR2_X1 U686 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(KEYINPUT99), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n616), .B(n615), .ZN(n677) );
  NAND2_X1 U690 ( .A1(G171), .A2(n617), .ZN(n664) );
  INV_X1 U691 ( .A(G1996), .ZN(n970) );
  XNOR2_X1 U692 ( .A(KEYINPUT26), .B(KEYINPUT93), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n619), .B(n618), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n669), .A2(G1341), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G56), .A2(n791), .ZN(n623) );
  XOR2_X1 U697 ( .A(KEYINPUT14), .B(n623), .Z(n630) );
  NAND2_X1 U698 ( .A1(G81), .A2(n795), .ZN(n624) );
  XOR2_X1 U699 ( .A(KEYINPUT73), .B(n624), .Z(n625) );
  XNOR2_X1 U700 ( .A(n625), .B(KEYINPUT12), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G68), .A2(n796), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U703 ( .A(KEYINPUT13), .B(n628), .Z(n629) );
  NOR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n792), .A2(G43), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n922) );
  NAND2_X1 U707 ( .A1(G79), .A2(n796), .ZN(n635) );
  NAND2_X1 U708 ( .A1(G54), .A2(n792), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U710 ( .A(KEYINPUT74), .B(n636), .ZN(n640) );
  NAND2_X1 U711 ( .A1(G66), .A2(n791), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G92), .A2(n795), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U715 ( .A(KEYINPUT15), .B(n641), .Z(n918) );
  NOR2_X1 U716 ( .A1(n644), .A2(n918), .ZN(n643) );
  INV_X1 U717 ( .A(KEYINPUT96), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n643), .B(n642), .ZN(n651) );
  NAND2_X1 U719 ( .A1(n644), .A2(n918), .ZN(n649) );
  INV_X1 U720 ( .A(G1348), .ZN(n919) );
  NOR2_X1 U721 ( .A1(n653), .A2(n919), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n645), .B(KEYINPUT95), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n653), .A2(G2067), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U727 ( .A1(n653), .A2(G2072), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(KEYINPUT27), .ZN(n655) );
  INV_X1 U729 ( .A(G1956), .ZN(n950) );
  NOR2_X1 U730 ( .A1(n950), .A2(n653), .ZN(n654) );
  NOR2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n658) );
  INV_X1 U732 ( .A(G299), .ZN(n771) );
  NAND2_X1 U733 ( .A1(n658), .A2(n771), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n657), .A2(n656), .ZN(n661) );
  NOR2_X1 U735 ( .A1(n658), .A2(n771), .ZN(n659) );
  XOR2_X1 U736 ( .A(n659), .B(KEYINPUT28), .Z(n660) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U738 ( .A(KEYINPUT29), .B(n662), .Z(n663) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n675) );
  AND2_X1 U740 ( .A1(n677), .A2(n675), .ZN(n665) );
  NOR2_X1 U741 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n684) );
  INV_X1 U743 ( .A(G8), .ZN(n674) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n708), .ZN(n671) );
  NOR2_X1 U745 ( .A1(G2090), .A2(n669), .ZN(n670) );
  NOR2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n672), .A2(G303), .ZN(n673) );
  OR2_X1 U748 ( .A1(n674), .A2(n673), .ZN(n678) );
  AND2_X1 U749 ( .A1(n675), .A2(n678), .ZN(n676) );
  NAND2_X1 U750 ( .A1(n677), .A2(n676), .ZN(n681) );
  INV_X1 U751 ( .A(n678), .ZN(n679) );
  OR2_X1 U752 ( .A1(n679), .A2(G286), .ZN(n680) );
  NAND2_X1 U753 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n682), .B(KEYINPUT32), .ZN(n683) );
  NAND2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n700) );
  NOR2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U758 ( .A1(n687), .A2(n685), .ZN(n931) );
  NAND2_X1 U759 ( .A1(n700), .A2(n931), .ZN(n686) );
  XNOR2_X1 U760 ( .A(n686), .B(KEYINPUT100), .ZN(n694) );
  XOR2_X1 U761 ( .A(G1981), .B(G305), .Z(n937) );
  INV_X1 U762 ( .A(n937), .ZN(n689) );
  NAND2_X1 U763 ( .A1(n687), .A2(KEYINPUT33), .ZN(n688) );
  NOR2_X1 U764 ( .A1(n689), .A2(n521), .ZN(n695) );
  INV_X1 U765 ( .A(n695), .ZN(n690) );
  OR2_X1 U766 ( .A1(n708), .A2(n690), .ZN(n692) );
  NAND2_X1 U767 ( .A1(G1976), .A2(G288), .ZN(n930) );
  AND2_X1 U768 ( .A1(n695), .A2(KEYINPUT33), .ZN(n696) );
  NOR2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n704) );
  NOR2_X1 U770 ( .A1(G2090), .A2(G303), .ZN(n698) );
  NAND2_X1 U771 ( .A1(G8), .A2(n698), .ZN(n699) );
  NAND2_X1 U772 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U773 ( .A1(n708), .A2(n701), .ZN(n702) );
  XOR2_X1 U774 ( .A(KEYINPUT101), .B(n702), .Z(n703) );
  NAND2_X1 U775 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U776 ( .A(n705), .B(KEYINPUT102), .ZN(n710) );
  NOR2_X1 U777 ( .A1(G1981), .A2(G305), .ZN(n706) );
  XOR2_X1 U778 ( .A(n706), .B(KEYINPUT24), .Z(n707) );
  NOR2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n747) );
  NAND2_X1 U781 ( .A1(G107), .A2(n519), .ZN(n712) );
  NAND2_X1 U782 ( .A1(G119), .A2(n879), .ZN(n711) );
  NAND2_X1 U783 ( .A1(n712), .A2(n711), .ZN(n717) );
  NAND2_X1 U784 ( .A1(G131), .A2(n714), .ZN(n715) );
  XNOR2_X1 U785 ( .A(KEYINPUT89), .B(n715), .ZN(n716) );
  NOR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U787 ( .A1(G95), .A2(n719), .ZN(n720) );
  NAND2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n890) );
  AND2_X1 U789 ( .A1(n890), .A2(G1991), .ZN(n730) );
  NAND2_X1 U790 ( .A1(G117), .A2(n519), .ZN(n723) );
  NAND2_X1 U791 ( .A1(G129), .A2(n879), .ZN(n722) );
  NAND2_X1 U792 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U793 ( .A1(n719), .A2(G105), .ZN(n724) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n724), .Z(n725) );
  NOR2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U796 ( .A1(n714), .A2(G141), .ZN(n727) );
  NAND2_X1 U797 ( .A1(n728), .A2(n727), .ZN(n875) );
  AND2_X1 U798 ( .A1(n875), .A2(G1996), .ZN(n729) );
  NOR2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n1009) );
  NOR2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n761) );
  INV_X1 U801 ( .A(n761), .ZN(n733) );
  NOR2_X1 U802 ( .A1(n1009), .A2(n733), .ZN(n753) );
  XOR2_X1 U803 ( .A(KEYINPUT90), .B(n753), .Z(n745) );
  NAND2_X1 U804 ( .A1(n714), .A2(G140), .ZN(n734) );
  XOR2_X1 U805 ( .A(KEYINPUT87), .B(n734), .Z(n736) );
  NAND2_X1 U806 ( .A1(G104), .A2(n719), .ZN(n735) );
  NAND2_X1 U807 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U808 ( .A(KEYINPUT34), .B(n737), .ZN(n742) );
  NAND2_X1 U809 ( .A1(G116), .A2(n519), .ZN(n739) );
  NAND2_X1 U810 ( .A1(G128), .A2(n879), .ZN(n738) );
  NAND2_X1 U811 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U812 ( .A(KEYINPUT35), .B(n740), .Z(n741) );
  NOR2_X1 U813 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U814 ( .A(KEYINPUT36), .B(n743), .ZN(n893) );
  XNOR2_X1 U815 ( .A(G2067), .B(KEYINPUT37), .ZN(n759) );
  NOR2_X1 U816 ( .A1(n893), .A2(n759), .ZN(n1001) );
  NAND2_X1 U817 ( .A1(n1001), .A2(n761), .ZN(n744) );
  XNOR2_X1 U818 ( .A(n744), .B(KEYINPUT88), .ZN(n757) );
  NAND2_X1 U819 ( .A1(n745), .A2(n757), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n750) );
  XNOR2_X1 U821 ( .A(G1986), .B(KEYINPUT86), .ZN(n748) );
  XNOR2_X1 U822 ( .A(n748), .B(G290), .ZN(n924) );
  NAND2_X1 U823 ( .A1(n924), .A2(n761), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n750), .A2(n749), .ZN(n764) );
  NOR2_X1 U825 ( .A1(G1996), .A2(n875), .ZN(n1004) );
  NOR2_X1 U826 ( .A1(G1986), .A2(G290), .ZN(n751) );
  NOR2_X1 U827 ( .A1(G1991), .A2(n890), .ZN(n996) );
  NOR2_X1 U828 ( .A1(n751), .A2(n996), .ZN(n752) );
  NOR2_X1 U829 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n1004), .A2(n754), .ZN(n755) );
  XOR2_X1 U831 ( .A(n755), .B(KEYINPUT103), .Z(n756) );
  XNOR2_X1 U832 ( .A(KEYINPUT39), .B(n756), .ZN(n758) );
  NAND2_X1 U833 ( .A1(n758), .A2(n757), .ZN(n760) );
  NAND2_X1 U834 ( .A1(n893), .A2(n759), .ZN(n1011) );
  NAND2_X1 U835 ( .A1(n760), .A2(n1011), .ZN(n762) );
  NAND2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n764), .A2(n763), .ZN(n766) );
  XNOR2_X1 U838 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n765) );
  XNOR2_X1 U839 ( .A(n766), .B(n765), .ZN(G329) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U841 ( .A(G57), .ZN(G237) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U843 ( .A(n767), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U844 ( .A(G223), .ZN(n830) );
  NAND2_X1 U845 ( .A1(n830), .A2(G567), .ZN(n768) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n768), .Z(G234) );
  INV_X1 U847 ( .A(G860), .ZN(n775) );
  OR2_X1 U848 ( .A1(n922), .A2(n775), .ZN(G153) );
  INV_X1 U849 ( .A(G171), .ZN(G301) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n770) );
  OR2_X1 U851 ( .A1(n918), .A2(G868), .ZN(n769) );
  NAND2_X1 U852 ( .A1(n770), .A2(n769), .ZN(G284) );
  INV_X1 U853 ( .A(G868), .ZN(n813) );
  NAND2_X1 U854 ( .A1(n771), .A2(n813), .ZN(n772) );
  XNOR2_X1 U855 ( .A(n772), .B(KEYINPUT77), .ZN(n774) );
  NOR2_X1 U856 ( .A1(G286), .A2(n813), .ZN(n773) );
  NOR2_X1 U857 ( .A1(n774), .A2(n773), .ZN(G297) );
  NAND2_X1 U858 ( .A1(n775), .A2(G559), .ZN(n776) );
  NAND2_X1 U859 ( .A1(n776), .A2(n918), .ZN(n777) );
  XNOR2_X1 U860 ( .A(n777), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U861 ( .A1(G868), .A2(n922), .ZN(n778) );
  XNOR2_X1 U862 ( .A(KEYINPUT78), .B(n778), .ZN(n781) );
  NAND2_X1 U863 ( .A1(G868), .A2(n918), .ZN(n779) );
  NOR2_X1 U864 ( .A1(G559), .A2(n779), .ZN(n780) );
  NOR2_X1 U865 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U866 ( .A1(G123), .A2(n879), .ZN(n782) );
  XNOR2_X1 U867 ( .A(n782), .B(KEYINPUT18), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n519), .A2(G111), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U870 ( .A1(G135), .A2(n714), .ZN(n786) );
  NAND2_X1 U871 ( .A1(G99), .A2(n719), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n995) );
  XNOR2_X1 U874 ( .A(n995), .B(G2096), .ZN(n790) );
  INV_X1 U875 ( .A(G2100), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(G156) );
  NAND2_X1 U877 ( .A1(G67), .A2(n791), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G55), .A2(n792), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n800) );
  NAND2_X1 U880 ( .A1(G93), .A2(n795), .ZN(n798) );
  NAND2_X1 U881 ( .A1(G80), .A2(n796), .ZN(n797) );
  NAND2_X1 U882 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U883 ( .A1(n800), .A2(n799), .ZN(n812) );
  NAND2_X1 U884 ( .A1(G559), .A2(n918), .ZN(n801) );
  XOR2_X1 U885 ( .A(n922), .B(n801), .Z(n810) );
  XNOR2_X1 U886 ( .A(KEYINPUT79), .B(n810), .ZN(n802) );
  NOR2_X1 U887 ( .A1(G860), .A2(n802), .ZN(n803) );
  XNOR2_X1 U888 ( .A(n812), .B(n803), .ZN(n804) );
  XNOR2_X1 U889 ( .A(n804), .B(KEYINPUT80), .ZN(G145) );
  XNOR2_X1 U890 ( .A(KEYINPUT19), .B(G305), .ZN(n805) );
  XNOR2_X1 U891 ( .A(n805), .B(G288), .ZN(n806) );
  XNOR2_X1 U892 ( .A(n812), .B(n806), .ZN(n808) );
  XNOR2_X1 U893 ( .A(G290), .B(G299), .ZN(n807) );
  XNOR2_X1 U894 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U895 ( .A(n809), .B(G303), .ZN(n896) );
  XNOR2_X1 U896 ( .A(n810), .B(n896), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n811), .A2(G868), .ZN(n815) );
  NAND2_X1 U898 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U899 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U900 ( .A(KEYINPUT83), .B(n816), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n817) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n817), .Z(n818) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n818), .ZN(n819) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n819), .ZN(n820) );
  NAND2_X1 U905 ( .A1(n820), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U907 ( .A1(G132), .A2(G82), .ZN(n821) );
  XNOR2_X1 U908 ( .A(n821), .B(KEYINPUT22), .ZN(n822) );
  XNOR2_X1 U909 ( .A(n822), .B(KEYINPUT84), .ZN(n823) );
  NOR2_X1 U910 ( .A1(G218), .A2(n823), .ZN(n824) );
  NAND2_X1 U911 ( .A1(G96), .A2(n824), .ZN(n834) );
  NAND2_X1 U912 ( .A1(n834), .A2(G2106), .ZN(n828) );
  NAND2_X1 U913 ( .A1(G120), .A2(G108), .ZN(n825) );
  NOR2_X1 U914 ( .A1(G237), .A2(n825), .ZN(n826) );
  NAND2_X1 U915 ( .A1(G69), .A2(n826), .ZN(n835) );
  NAND2_X1 U916 ( .A1(n835), .A2(G567), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n836) );
  NAND2_X1 U918 ( .A1(G483), .A2(G661), .ZN(n829) );
  NOR2_X1 U919 ( .A1(n836), .A2(n829), .ZN(n833) );
  NAND2_X1 U920 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U923 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U926 ( .A(G108), .B(KEYINPUT112), .Z(G238) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G82), .ZN(G220) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n836), .ZN(G319) );
  XNOR2_X1 U934 ( .A(G1996), .B(KEYINPUT41), .ZN(n846) );
  XOR2_X1 U935 ( .A(G1956), .B(G1966), .Z(n838) );
  XNOR2_X1 U936 ( .A(G1991), .B(G1986), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U938 ( .A(G1961), .B(G1971), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1981), .B(G1976), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U942 ( .A(KEYINPUT106), .B(G2474), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(G229) );
  XOR2_X1 U945 ( .A(G2100), .B(G2096), .Z(n848) );
  XNOR2_X1 U946 ( .A(KEYINPUT42), .B(G2678), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U948 ( .A(KEYINPUT43), .B(G2090), .Z(n850) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U951 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U952 ( .A(G2078), .B(G2084), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(G227) );
  NAND2_X1 U954 ( .A1(G124), .A2(n879), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n519), .A2(G112), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G136), .A2(n714), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G100), .A2(n719), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U961 ( .A1(n861), .A2(n860), .ZN(G162) );
  NAND2_X1 U962 ( .A1(G142), .A2(n714), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G106), .A2(n719), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT45), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G118), .A2(n519), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G130), .A2(n879), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U969 ( .A(KEYINPUT107), .B(n867), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n870), .B(G162), .ZN(n874) );
  XOR2_X1 U972 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n872) );
  XNOR2_X1 U973 ( .A(n995), .B(KEYINPUT48), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U975 ( .A(n874), .B(n873), .Z(n877) );
  XOR2_X1 U976 ( .A(G164), .B(n875), .Z(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n889) );
  NAND2_X1 U978 ( .A1(G115), .A2(n519), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G127), .A2(n879), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(KEYINPUT47), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G103), .A2(n719), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n887) );
  NAND2_X1 U984 ( .A1(n714), .A2(G139), .ZN(n885) );
  XOR2_X1 U985 ( .A(KEYINPUT108), .B(n885), .Z(n886) );
  NOR2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U987 ( .A(KEYINPUT109), .B(n888), .Z(n1014) );
  XOR2_X1 U988 ( .A(n889), .B(n1014), .Z(n892) );
  XOR2_X1 U989 ( .A(G160), .B(n890), .Z(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U992 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U993 ( .A(G286), .B(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(G171), .B(n918), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n922), .B(KEYINPUT111), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(G397) );
  XOR2_X1 U999 ( .A(G2454), .B(G2430), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G2451), .B(G2446), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n910) );
  XOR2_X1 U1002 ( .A(G2443), .B(G2427), .Z(n905) );
  XNOR2_X1 U1003 ( .A(G2438), .B(KEYINPUT105), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1005 ( .A(n906), .B(G2435), .Z(n908) );
  XNOR2_X1 U1006 ( .A(G1348), .B(G1341), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n911), .A2(G14), .ZN(n917) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n917), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G96), .ZN(G221) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  INV_X1 U1019 ( .A(n917), .ZN(G401) );
  XOR2_X1 U1020 ( .A(KEYINPUT56), .B(G16), .Z(n944) );
  XNOR2_X1 U1021 ( .A(G301), .B(G1961), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(G1341), .B(n922), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n929) );
  XOR2_X1 U1027 ( .A(G1956), .B(G299), .Z(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT123), .B(n927), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n936) );
  AND2_X1 U1030 ( .A1(G303), .A2(G1971), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT124), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(G1966), .B(G168), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1037 ( .A(KEYINPUT57), .B(n939), .Z(n940) );
  NOR2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1039 ( .A(KEYINPUT125), .B(n942), .Z(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n1029) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G21), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n945), .B(G5), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n959) );
  XOR2_X1 U1044 ( .A(KEYINPUT126), .B(G4), .Z(n949) );
  XNOR2_X1 U1045 ( .A(G1348), .B(KEYINPUT59), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n949), .B(n948), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(G20), .B(n950), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G1981), .B(G6), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(G1341), .B(G19), .ZN(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(KEYINPUT60), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(G1976), .B(G23), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n963) );
  XOR2_X1 U1058 ( .A(G1986), .B(G24), .Z(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(KEYINPUT58), .B(n964), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1062 ( .A(KEYINPUT61), .B(n967), .Z(n968) );
  NOR2_X1 U1063 ( .A1(G16), .A2(n968), .ZN(n994) );
  XOR2_X1 U1064 ( .A(G25), .B(G1991), .Z(n969) );
  NAND2_X1 U1065 ( .A1(n969), .A2(G28), .ZN(n973) );
  XOR2_X1 U1066 ( .A(KEYINPUT120), .B(n970), .Z(n971) );
  XNOR2_X1 U1067 ( .A(G32), .B(n971), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(n974), .B(G27), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G2067), .B(G26), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(G2072), .B(G33), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(KEYINPUT119), .B(n977), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(n982), .B(KEYINPUT53), .ZN(n985) );
  XOR2_X1 U1077 ( .A(G2084), .B(G34), .Z(n983) );
  XNOR2_X1 U1078 ( .A(KEYINPUT54), .B(n983), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(G35), .B(G2090), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1082 ( .A(KEYINPUT55), .B(n988), .Z(n989) );
  NOR2_X1 U1083 ( .A1(G29), .A2(n989), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(KEYINPUT121), .B(n990), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n991), .A2(G11), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(n992), .B(KEYINPUT122), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n1027) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1089 ( .A(KEYINPUT113), .B(n997), .Z(n999) );
  XNOR2_X1 U1090 ( .A(G160), .B(G2084), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1093 ( .A(KEYINPUT114), .B(n1002), .Z(n1007) );
  XOR2_X1 U1094 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(KEYINPUT51), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(n1010), .B(KEYINPUT115), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT116), .B(n1013), .ZN(n1021) );
  XNOR2_X1 U1102 ( .A(G2072), .B(n1014), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(G164), .B(G2078), .Z(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT117), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(n1018), .B(KEYINPUT118), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(n1019), .B(KEYINPUT50), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT52), .B(n1022), .ZN(n1024) );
  INV_X1 U1110 ( .A(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(G29), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1115 ( .A(KEYINPUT127), .B(n1030), .Z(n1031) );
  XNOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1031), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

