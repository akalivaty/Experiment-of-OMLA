//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246, new_n1247;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n460), .A2(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT71), .B(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT72), .B1(new_n465), .B2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n467), .A3(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n476), .A3(new_n466), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n479), .A2(new_n481), .A3(G137), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n473), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT73), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g060(.A(KEYINPUT73), .B(new_n473), .C1(new_n477), .C2(new_n482), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n471), .B1(new_n485), .B2(new_n486), .ZN(G160));
  NOR2_X1   g062(.A1(new_n477), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n464), .A2(G112), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n474), .A2(new_n476), .A3(new_n466), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n479), .A2(new_n481), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G124), .ZN(new_n496));
  OR3_X1    g071(.A1(new_n495), .A2(KEYINPUT74), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT74), .B1(new_n495), .B2(new_n496), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n492), .B1(new_n497), .B2(new_n498), .ZN(G162));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n466), .A2(new_n468), .A3(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n494), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(G126), .A2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT4), .A2(G138), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(new_n464), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n502), .B(new_n506), .C1(new_n477), .C2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n513), .B1(new_n518), .B2(KEYINPUT77), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT5), .B(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT77), .A3(G62), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(G651), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT75), .B1(new_n524), .B2(KEYINPUT76), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT6), .B1(new_n524), .B2(KEYINPUT75), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g102(.A(KEYINPUT75), .B(KEYINPUT6), .C1(new_n524), .C2(KEYINPUT76), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n527), .A2(G50), .A3(G543), .A4(new_n528), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n527), .A2(G88), .A3(new_n520), .A4(new_n528), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  AND2_X1   g109(.A1(new_n527), .A2(new_n528), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G51), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n535), .A2(new_n520), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT78), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n538), .A2(new_n540), .A3(new_n542), .A4(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n537), .A2(G52), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n539), .A2(G90), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n524), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND3_X1  g127(.A1(new_n535), .A2(G43), .A3(G543), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n527), .A2(G81), .A3(new_n520), .A4(new_n528), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n516), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND4_X1  g139(.A1(new_n527), .A2(G53), .A3(G543), .A4(new_n528), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n516), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n527), .A2(G91), .A3(new_n520), .A4(new_n528), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT79), .ZN(new_n574));
  NOR3_X1   g149(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n576), .A2(new_n577), .B1(G651), .B2(new_n569), .ZN(new_n578));
  INV_X1    g153(.A(new_n574), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT80), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n575), .A2(new_n580), .ZN(G299));
  NAND4_X1  g156(.A1(new_n527), .A2(G87), .A3(new_n520), .A4(new_n528), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n527), .A2(G49), .A3(G543), .A4(new_n528), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n582), .A2(new_n583), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n584), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT82), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(KEYINPUT82), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(G288));
  NAND4_X1  g167(.A1(new_n527), .A2(G86), .A3(new_n520), .A4(new_n528), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n527), .A2(G48), .A3(G543), .A4(new_n528), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n520), .B2(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n596), .B1(new_n599), .B2(new_n524), .ZN(new_n600));
  OAI21_X1  g175(.A(G61), .B1(new_n514), .B2(new_n515), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(new_n597), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n602), .A2(KEYINPUT83), .A3(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n595), .B1(new_n604), .B2(KEYINPUT84), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n600), .A2(new_n606), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n537), .A2(G47), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n539), .A2(G85), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n609), .B(new_n610), .C1(new_n524), .C2(new_n611), .ZN(G290));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  OR3_X1    g188(.A1(G171), .A2(KEYINPUT85), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT85), .B1(G171), .B2(new_n613), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(new_n524), .ZN(new_n617));
  INV_X1    g192(.A(G54), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n536), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n535), .A2(new_n520), .ZN(new_n622));
  INV_X1    g197(.A(G92), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n619), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n614), .B(new_n615), .C1(G868), .C2(new_n625), .ZN(G284));
  OAI211_X1 g201(.A(new_n614), .B(new_n615), .C1(G868), .C2(new_n625), .ZN(G321));
  NAND2_X1  g202(.A1(G299), .A2(new_n613), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n613), .B2(G168), .ZN(G280));
  XNOR2_X1  g204(.A(G280), .B(KEYINPUT86), .ZN(G297));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n625), .B1(new_n631), .B2(G860), .ZN(G148));
  INV_X1    g207(.A(new_n559), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(new_n613), .ZN(new_n634));
  INV_X1    g209(.A(new_n625), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n635), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n634), .B1(new_n636), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XOR2_X1   g213(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n639));
  NOR3_X1   g214(.A1(new_n465), .A2(new_n467), .A3(G2105), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n488), .A2(G135), .ZN(new_n645));
  OAI221_X1 g220(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n646));
  INV_X1    g221(.A(G123), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n495), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(G2096), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(G2096), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n644), .A2(new_n649), .A3(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT90), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT89), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT14), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G14), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n659), .A2(new_n665), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT17), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n673), .B(KEYINPUT92), .Z(new_n678));
  INV_X1    g253(.A(new_n672), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n680), .A2(new_n671), .ZN(new_n681));
  INV_X1    g256(.A(new_n678), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n672), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n671), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n676), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1971), .B(G1976), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n690), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT93), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n695), .B(new_n697), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(new_n693), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT20), .Z(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT94), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1981), .B(G1986), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT95), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n704), .B(new_n708), .ZN(G229));
  NAND2_X1  g284(.A1(G299), .A2(G16), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G20), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT23), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1956), .ZN(new_n715));
  INV_X1    g290(.A(G28), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT30), .ZN(new_n717));
  AOI21_X1  g292(.A(G29), .B1(new_n716), .B2(KEYINPUT30), .ZN(new_n718));
  OR2_X1    g293(.A1(KEYINPUT31), .A2(G11), .ZN(new_n719));
  NAND2_X1  g294(.A1(KEYINPUT31), .A2(G11), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n717), .A2(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(G164), .A2(G29), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G27), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2078), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n721), .B1(new_n722), .B2(new_n648), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(G301), .A2(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n711), .A2(G5), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n726), .B1(new_n730), .B2(G1961), .ZN(new_n731));
  INV_X1    g306(.A(G1341), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n559), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G16), .B2(G19), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT97), .B(KEYINPUT26), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G105), .B2(new_n472), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n488), .A2(G141), .ZN(new_n739));
  INV_X1    g314(.A(G129), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n495), .ZN(new_n741));
  MUX2_X1   g316(.A(G32), .B(new_n741), .S(G29), .Z(new_n742));
  XOR2_X1   g317(.A(KEYINPUT27), .B(G1996), .Z(new_n743));
  OAI221_X1 g318(.A(new_n731), .B1(new_n732), .B2(new_n734), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G34), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(G29), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G160), .B2(G29), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G2084), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n711), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n711), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n742), .A2(new_n743), .B1(new_n732), .B2(new_n734), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n722), .A2(G33), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n466), .A2(new_n468), .A3(G127), .ZN(new_n757));
  INV_X1    g332(.A(G115), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(new_n467), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n760));
  NAND2_X1  g335(.A1(G103), .A2(G2104), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n494), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n494), .A2(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n488), .A2(G139), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n756), .B1(new_n766), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2072), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n724), .A2(new_n725), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n748), .A2(G2084), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n769), .B(new_n770), .C1(new_n768), .C2(new_n767), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n744), .A2(new_n749), .A3(new_n755), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n722), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n722), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT29), .B(G2090), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n711), .A2(G4), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n625), .B2(new_n711), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n722), .A2(G26), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT28), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n488), .A2(G140), .ZN(new_n783));
  OAI221_X1 g358(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n784));
  INV_X1    g359(.A(G128), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n495), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n782), .B1(new_n787), .B2(new_n722), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(G2067), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(G2067), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G1961), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n789), .B(new_n791), .C1(new_n792), .C2(new_n729), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n772), .A2(new_n776), .A3(new_n780), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n711), .A2(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n711), .ZN(new_n796));
  INV_X1    g371(.A(G1971), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n711), .A2(G6), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G305), .B2(G16), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n798), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n711), .A2(G23), .ZN(new_n804));
  INV_X1    g379(.A(new_n589), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n711), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT33), .B(G1976), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n799), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n801), .ZN(new_n810));
  OR3_X1    g385(.A1(new_n803), .A2(new_n810), .A3(KEYINPUT34), .ZN(new_n811));
  OAI21_X1  g386(.A(KEYINPUT34), .B1(new_n803), .B2(new_n810), .ZN(new_n812));
  MUX2_X1   g387(.A(G24), .B(G290), .S(G16), .Z(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G1986), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n722), .A2(G25), .ZN(new_n815));
  OAI221_X1 g390(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n816));
  INV_X1    g391(.A(G119), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n495), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G131), .B2(new_n488), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n815), .B1(new_n819), .B2(new_n722), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n811), .A2(new_n812), .A3(new_n814), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n826));
  AOI211_X1 g401(.A(new_n715), .B(new_n794), .C1(new_n825), .C2(new_n826), .ZN(G311));
  INV_X1    g402(.A(G311), .ZN(G150));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  INV_X1    g404(.A(G80), .ZN(new_n830));
  INV_X1    g405(.A(G543), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n516), .A2(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI221_X1 g409(.A(KEYINPUT98), .B1(new_n830), .B2(new_n831), .C1(new_n516), .C2(new_n829), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(G651), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT99), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT99), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n834), .A2(new_n838), .A3(new_n835), .A4(G651), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n527), .A2(G55), .A3(G543), .A4(new_n528), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n527), .A2(G93), .A3(new_n520), .A4(new_n528), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n837), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n625), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n633), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n842), .B1(new_n836), .B2(KEYINPUT99), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n850), .A2(new_n559), .A3(new_n839), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n848), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT100), .Z(new_n856));
  INV_X1    g431(.A(G860), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n846), .B1(new_n856), .B2(new_n858), .ZN(G145));
  XNOR2_X1  g434(.A(new_n741), .B(new_n766), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n819), .B(new_n641), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n511), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n479), .A2(new_n481), .A3(new_n509), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n507), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n493), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n867), .A2(KEYINPUT101), .A3(new_n502), .A4(new_n506), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n787), .ZN(new_n870));
  OAI221_X1 g445(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n871));
  INV_X1    g446(.A(G130), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n495), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(G142), .B2(new_n488), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n870), .B(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n862), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n862), .A2(new_n875), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(G160), .B(new_n648), .Z(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(G162), .Z(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT102), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n878), .B2(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g461(.A(new_n635), .B1(new_n575), .B2(new_n580), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n572), .B1(new_n571), .B2(new_n574), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT80), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n625), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n636), .B(new_n852), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n891), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(KEYINPUT42), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n897), .B(new_n899), .C1(new_n901), .C2(KEYINPUT42), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(G290), .B(G303), .ZN(new_n906));
  XNOR2_X1  g481(.A(G305), .B(new_n805), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n901), .B2(KEYINPUT42), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n903), .A2(new_n910), .A3(new_n904), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n613), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n844), .A2(new_n613), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n914), .A2(KEYINPUT104), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n918));
  INV_X1    g493(.A(new_n913), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n910), .B1(new_n903), .B2(new_n904), .ZN(new_n920));
  OAI21_X1  g495(.A(G868), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n921), .B2(new_n915), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n917), .A2(new_n922), .ZN(G295));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n915), .ZN(G331));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n850), .A2(new_n559), .A3(new_n839), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n559), .B1(new_n850), .B2(new_n839), .ZN(new_n927));
  OAI21_X1  g502(.A(G171), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n849), .A2(G301), .A3(new_n851), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n928), .A2(G168), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G168), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n891), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n929), .ZN(new_n935));
  AOI21_X1  g510(.A(G301), .B1(new_n849), .B2(new_n851), .ZN(new_n936));
  OAI21_X1  g511(.A(G286), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n928), .A2(G168), .A3(new_n929), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(KEYINPUT106), .A3(new_n891), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n893), .A2(new_n894), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n939), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n895), .A2(KEYINPUT105), .A3(new_n938), .A4(new_n937), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n941), .A2(new_n944), .A3(new_n909), .A4(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n932), .B1(new_n943), .B2(new_n939), .ZN(new_n947));
  AOI21_X1  g522(.A(G37), .B1(new_n947), .B2(new_n908), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n948), .A3(KEYINPUT107), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(KEYINPUT43), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n954), .B2(new_n908), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n946), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n925), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n955), .B2(new_n946), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n946), .A2(new_n956), .A3(new_n948), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n958), .A2(new_n961), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT127), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n864), .A2(new_n964), .A3(new_n868), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n485), .A2(new_n486), .ZN(new_n968));
  INV_X1    g543(.A(new_n471), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(G40), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n741), .B(G1996), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n786), .B(G2067), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT108), .B(new_n971), .C1(new_n972), .C2(new_n973), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n819), .B(new_n821), .Z(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n971), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  NOR2_X1   g558(.A1(G290), .A2(G1986), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n971), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n605), .A2(new_n987), .A3(new_n988), .A4(new_n607), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT83), .B1(new_n602), .B2(G651), .ZN(new_n990));
  AOI211_X1 g565(.A(new_n596), .B(new_n524), .C1(new_n601), .C2(new_n597), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT84), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n595), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n607), .A3(new_n988), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT113), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n595), .A2(KEYINPUT114), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(new_n603), .A3(new_n600), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n595), .A2(KEYINPUT114), .ZN(new_n999));
  OAI21_X1  g574(.A(G1981), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  INV_X1    g579(.A(G40), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n1005), .B(new_n471), .C1(new_n485), .C2(new_n486), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n505), .B1(new_n866), .B2(new_n493), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1007), .B2(new_n502), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n1000), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n584), .A2(new_n587), .A3(G1976), .A4(new_n588), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(KEYINPUT112), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1009), .A2(new_n1014), .A3(new_n1018), .A4(new_n1015), .ZN(new_n1021));
  NOR2_X1   g596(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n590), .A2(new_n591), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1011), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1026));
  NAND3_X1  g601(.A1(new_n511), .A2(new_n964), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1008), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(new_n970), .ZN(new_n1030));
  INV_X1    g605(.A(G2090), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n864), .A2(KEYINPUT45), .A3(new_n964), .A4(new_n868), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(G160), .B(G40), .C1(new_n1008), .C2(KEYINPUT45), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n797), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1004), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n520), .A2(G62), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT77), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1039), .A2(new_n1040), .B1(G75), .B2(G543), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n524), .B1(new_n1041), .B2(new_n521), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT55), .B(G8), .C1(new_n1042), .C2(new_n531), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1038), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1037), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1025), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1009), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1003), .A2(new_n1010), .ZN(new_n1050));
  NOR2_X1   g625(.A1(G288), .A2(G1976), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1049), .B1(new_n1052), .B2(new_n996), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n511), .A2(new_n964), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT50), .ZN(new_n1056));
  INV_X1    g631(.A(G2084), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1006), .A2(new_n1056), .A3(new_n1057), .A4(new_n1027), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n966), .B(G1384), .C1(new_n1007), .C2(new_n502), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT45), .B1(new_n511), .B2(new_n964), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n970), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(G168), .B(new_n1058), .C1(new_n1061), .C2(G1966), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1055), .A2(new_n966), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1008), .A2(KEYINPUT45), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1006), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n752), .ZN(new_n1067));
  AOI21_X1  g642(.A(G168), .B1(new_n1067), .B2(new_n1058), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT51), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1062), .A2(new_n1070), .A3(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT62), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1033), .A2(new_n725), .A3(new_n1006), .A4(new_n1064), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1006), .A2(new_n1056), .A3(new_n1027), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1074), .A2(new_n1075), .B1(new_n1076), .B2(new_n792), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n970), .A2(new_n1060), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1075), .A2(G2078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1065), .ZN(new_n1080));
  AOI21_X1  g655(.A(G301), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1069), .A2(new_n1082), .A3(new_n1071), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1073), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n1000), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT49), .B1(new_n996), .B2(new_n1000), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1049), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1011), .A2(KEYINPUT116), .A3(new_n1024), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1004), .B(new_n1045), .C1(new_n1036), .C2(new_n1032), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1026), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1055), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n511), .A2(new_n1028), .A3(new_n964), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1006), .A2(new_n1094), .A3(new_n1031), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1004), .B1(new_n1036), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT115), .B1(new_n1097), .B2(new_n1046), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1971), .B1(new_n1078), .B2(new_n1033), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1096), .ZN(new_n1100));
  OAI21_X1  g675(.A(G8), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(new_n1102), .A3(new_n1045), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1092), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1090), .A2(new_n1091), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1054), .B1(new_n1084), .B2(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1037), .A2(new_n1046), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1067), .A2(new_n1058), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1108), .A2(new_n1004), .A3(G286), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1107), .A2(KEYINPUT63), .A3(new_n1047), .A4(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(new_n1025), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1090), .A2(new_n1091), .A3(new_n1104), .A4(new_n1109), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n779), .B1(new_n1029), .B2(new_n970), .ZN(new_n1116));
  INV_X1    g691(.A(G2067), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1006), .A2(new_n1117), .A3(new_n1008), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n625), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1119), .A2(new_n1120), .A3(new_n635), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(KEYINPUT60), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT123), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT58), .B(G1341), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(G1996), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1033), .A2(new_n1133), .A3(new_n1006), .A4(new_n1064), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n633), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1135), .B(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT56), .B(G2072), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1078), .A2(new_n1033), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(G1956), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1095), .B1(new_n1008), .B2(new_n1026), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT117), .B(new_n1141), .C1(new_n1142), .C2(new_n970), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1006), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT117), .B1(new_n1145), .B2(new_n1141), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1140), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT57), .B1(new_n566), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n571), .B2(new_n574), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT118), .B1(new_n576), .B2(new_n577), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n578), .B(new_n579), .C1(new_n1151), .C2(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1147), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1140), .B(new_n1153), .C1(new_n1144), .C2(new_n1146), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1138), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1141), .B1(new_n1142), .B2(new_n970), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1164), .A2(new_n1143), .B1(new_n1165), .B2(new_n1139), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1166), .A2(KEYINPUT121), .A3(new_n1153), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1154), .B1(new_n1166), .B2(KEYINPUT119), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT119), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1147), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1161), .B(new_n1167), .C1(new_n1168), .C2(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1119), .A2(new_n1120), .A3(new_n635), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n635), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1173));
  OAI22_X1  g748(.A1(new_n1172), .A2(new_n1173), .B1(new_n1120), .B2(new_n1119), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1128), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1129), .A2(new_n1159), .A3(new_n1171), .A4(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1127), .A2(new_n635), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1179), .B1(new_n1156), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1076), .A2(new_n792), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1183), .A2(G301), .A3(new_n1080), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT124), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n967), .A2(new_n1006), .A3(new_n1033), .A4(new_n1079), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1183), .A2(new_n1184), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(G171), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1077), .A2(new_n1190), .A3(G301), .A4(new_n1080), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1186), .A2(new_n1189), .A3(KEYINPUT54), .A4(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT54), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1077), .A2(G301), .A3(new_n1187), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1193), .B1(new_n1194), .B2(new_n1081), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1072), .A2(new_n1192), .A3(new_n1195), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1097), .A2(KEYINPUT115), .A3(new_n1046), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1102), .B1(new_n1101), .B2(new_n1045), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1047), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(KEYINPUT116), .B1(new_n1011), .B2(new_n1024), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AND3_X1   g776(.A1(new_n1196), .A2(new_n1091), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1182), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n986), .B1(new_n1115), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n971), .A2(new_n984), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT48), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n982), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n971), .B1(new_n741), .B2(new_n973), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT126), .Z(new_n1209));
  NAND2_X1  g784(.A1(new_n971), .A2(new_n1133), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT46), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1212), .A2(KEYINPUT47), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1212), .A2(KEYINPUT47), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1207), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n978), .A2(new_n821), .A3(new_n819), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n787), .A2(new_n1117), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(KEYINPUT125), .B1(new_n1218), .B2(new_n971), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g795(.A1(new_n1218), .A2(KEYINPUT125), .A3(new_n971), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n963), .B1(new_n1204), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(new_n986), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1226));
  INV_X1    g801(.A(new_n1111), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI22_X1  g803(.A1(new_n1050), .A2(new_n1051), .B1(new_n995), .B2(new_n989), .ZN(new_n1229));
  OAI22_X1  g804(.A1(new_n1229), .A2(new_n1049), .B1(new_n1025), .B2(new_n1047), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1083), .A2(new_n1081), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1082), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AND3_X1   g808(.A1(new_n1090), .A2(new_n1091), .A3(new_n1104), .ZN(new_n1234));
  AOI21_X1  g809(.A(new_n1230), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1228), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1196), .A2(new_n1201), .A3(new_n1091), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1237), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1238));
  OAI21_X1  g813(.A(new_n1225), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  NOR3_X1   g814(.A1(new_n1221), .A2(new_n1215), .A3(new_n1219), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1239), .A2(KEYINPUT127), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1224), .A2(new_n1241), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g817(.A(G319), .B1(new_n667), .B2(new_n668), .ZN(new_n1244));
  NOR3_X1   g818(.A1(G229), .A2(G227), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g819(.A1(new_n885), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g820(.A1(new_n959), .A2(new_n960), .ZN(new_n1247));
  NOR2_X1   g821(.A1(new_n1246), .A2(new_n1247), .ZN(G308));
  OR2_X1    g822(.A1(new_n1246), .A2(new_n1247), .ZN(G225));
endmodule


