//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT66), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n189), .B2(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .A4(new_n194), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n203), .B(new_n205), .C1(KEYINPUT1), .C2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n204), .A2(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(G143), .ZN(new_n210));
  OAI211_X1 g024(.A(G128), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n196), .A2(new_n201), .A3(new_n207), .A4(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n203), .A2(new_n205), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT0), .B(G128), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n198), .A2(new_n199), .A3(new_n194), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n217), .B1(new_n219), .B2(new_n201), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n212), .B1(new_n220), .B2(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n201), .ZN(new_n222));
  INV_X1    g036(.A(new_n217), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n222), .A2(KEYINPUT65), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n188), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G116), .ZN(new_n228));
  INV_X1    g042(.A(G116), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT67), .A3(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n229), .A2(G119), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT2), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT2), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G113), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT68), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n232), .B1(new_n228), .B2(new_n230), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(new_n238), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n241), .A2(new_n238), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n211), .A2(new_n207), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n248), .A2(KEYINPUT69), .A3(new_n201), .A4(new_n196), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n211), .A2(new_n201), .A3(new_n207), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n195), .A2(G131), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n222), .A2(new_n223), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n249), .A2(new_n253), .A3(KEYINPUT30), .A4(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n225), .A2(new_n247), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n245), .B1(new_n240), .B2(new_n243), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n249), .A2(new_n257), .A3(new_n253), .A4(new_n254), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(G210), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n261), .A3(G210), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n267), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n265), .B1(new_n269), .B2(new_n263), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(new_n268), .B2(new_n270), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n260), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n247), .B1(new_n221), .B2(new_n224), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(new_n258), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n247), .A2(new_n220), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT28), .B1(new_n279), .B2(new_n212), .ZN(new_n280));
  INV_X1    g094(.A(new_n274), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  OR3_X1    g096(.A1(new_n275), .A2(KEYINPUT29), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n249), .A2(new_n253), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n247), .B1(new_n285), .B2(new_n220), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n258), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n280), .B1(new_n287), .B2(KEYINPUT28), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n274), .A2(KEYINPUT29), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n187), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n281), .B1(new_n278), .B2(new_n280), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n258), .A2(new_n274), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT72), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n258), .A2(new_n297), .A3(new_n274), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT31), .B1(new_n299), .B2(new_n256), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n258), .A2(new_n297), .A3(new_n274), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n297), .B1(new_n258), .B2(new_n274), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n256), .B(KEYINPUT31), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n294), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n256), .B1(new_n301), .B2(new_n302), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT31), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n303), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT73), .A3(new_n294), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n293), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n314), .ZN(new_n316));
  AOI211_X1 g130(.A(KEYINPUT32), .B(new_n316), .C1(new_n307), .C2(new_n312), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n292), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G475), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G125), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT76), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT74), .B1(new_n321), .B2(G125), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(G125), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n325), .A2(new_n328), .B1(G125), .B2(new_n321), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT75), .B1(new_n334), .B2(KEYINPUT16), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n324), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n202), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(G143), .B1(new_n262), .B2(G214), .ZN(new_n340));
  OAI21_X1  g154(.A(G131), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n340), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n200), .A3(new_n338), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT17), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n345), .A2(KEYINPUT94), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n341), .A2(new_n344), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n345), .B2(KEYINPUT94), .ZN(new_n348));
  OAI211_X1 g162(.A(G146), .B(new_n324), .C1(new_n333), .C2(new_n335), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n337), .A2(new_n346), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n342), .A2(new_n338), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT18), .A2(G131), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G125), .B(G140), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n354), .A2(new_n202), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n334), .B2(new_n202), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n350), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G113), .B(G122), .ZN(new_n360));
  INV_X1    g174(.A(G104), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n350), .A2(new_n362), .A3(new_n358), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G902), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n319), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT96), .ZN(new_n369));
  INV_X1    g183(.A(G478), .ZN(new_n370));
  NOR2_X1   g184(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  INV_X1    g190(.A(G217), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n376), .A2(new_n377), .A3(G953), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n204), .A2(G128), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n206), .A2(G143), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(new_n189), .ZN(new_n382));
  XNOR2_X1  g196(.A(G116), .B(G122), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n229), .A2(KEYINPUT14), .A3(G122), .ZN(new_n386));
  INV_X1    g200(.A(new_n383), .ZN(new_n387));
  OAI211_X1 g201(.A(G107), .B(new_n386), .C1(new_n387), .C2(KEYINPUT14), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n379), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n380), .B1(new_n390), .B2(KEYINPUT13), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n379), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G134), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n383), .B(new_n384), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n381), .A2(new_n189), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n378), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n389), .A2(new_n397), .A3(new_n378), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n375), .B1(new_n401), .B2(new_n367), .ZN(new_n402));
  INV_X1    g216(.A(new_n400), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n367), .B(new_n375), .C1(new_n403), .C2(new_n398), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n369), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(G234), .A2(G237), .ZN(new_n407));
  INV_X1    g221(.A(G953), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(G952), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT21), .B(G898), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(G902), .A3(G953), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n403), .A2(new_n398), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n374), .B1(new_n414), .B2(G902), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT96), .A3(new_n404), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n406), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(G475), .A2(G902), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n329), .A2(new_n330), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT19), .ZN(new_n420));
  AND2_X1   g234(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n421));
  NOR2_X1   g235(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT91), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n354), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n354), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT91), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n420), .A2(new_n202), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT92), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n423), .A2(new_n354), .A3(new_n424), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n424), .B1(new_n423), .B2(new_n354), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n202), .A4(new_n420), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n341), .A2(new_n343), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n429), .A2(new_n349), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n358), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT93), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n363), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n365), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n438), .B1(new_n437), .B2(new_n363), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n418), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT20), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n444), .B(new_n418), .C1(new_n440), .C2(new_n441), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n368), .B(new_n417), .C1(new_n443), .C2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n217), .A2(G125), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n217), .A2(KEYINPUT85), .A3(G125), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(KEYINPUT86), .A3(new_n452), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n248), .A2(G125), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n408), .A2(G224), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n459), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n361), .A2(G107), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n384), .A2(KEYINPUT3), .A3(G104), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT3), .B1(new_n384), .B2(G104), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT4), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n467), .A3(G101), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(G101), .ZN(new_n469));
  INV_X1    g283(.A(G101), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n470), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(KEYINPUT4), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n247), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT80), .B1(new_n384), .B2(G104), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT80), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n361), .A3(G107), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n384), .A2(G104), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n471), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n234), .B1(new_n482), .B2(new_n232), .ZN(new_n483));
  INV_X1    g297(.A(new_n241), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n482), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n244), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n473), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT84), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT84), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n473), .A2(new_n490), .A3(new_n486), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G122), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n488), .A2(new_n489), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n473), .A2(new_n490), .A3(new_n486), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n490), .B1(new_n473), .B2(new_n486), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n495), .A2(new_n496), .A3(new_n492), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n473), .A2(new_n486), .A3(new_n492), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n462), .B(new_n494), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n460), .A2(KEYINPUT7), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n453), .B2(new_n457), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT88), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT7), .B1(new_n460), .B2(KEYINPUT89), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(KEYINPUT89), .B2(new_n460), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n455), .A2(new_n456), .A3(new_n458), .A4(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(new_n501), .C1(new_n453), .C2(new_n457), .ZN(new_n508));
  AND4_X1   g322(.A1(new_n498), .A2(new_n503), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n481), .B1(new_n244), .B2(new_n485), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n483), .B1(new_n484), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n244), .A2(new_n481), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n492), .B(KEYINPUT8), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(G902), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n500), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G210), .B1(G237), .B2(G902), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n500), .A2(new_n520), .A3(new_n522), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n448), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G221), .ZN(new_n527));
  INV_X1    g341(.A(new_n376), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(new_n367), .ZN(new_n529));
  XNOR2_X1  g343(.A(G110), .B(G140), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n408), .A2(G227), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT79), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n479), .A2(new_n471), .A3(new_n207), .A4(new_n211), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT10), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT10), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n248), .A2(new_n537), .A3(new_n471), .A4(new_n479), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n219), .A2(new_n201), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n472), .A2(new_n223), .A3(new_n468), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n211), .A2(new_n207), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n480), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n540), .B1(new_n544), .B2(new_n535), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT12), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n547), .B(new_n540), .C1(new_n544), .C2(new_n535), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n542), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT81), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT81), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n542), .B(new_n551), .C1(new_n546), .C2(new_n548), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n534), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n554), .A2(new_n555), .A3(new_n532), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n367), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G469), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n532), .B1(new_n554), .B2(new_n555), .ZN(new_n559));
  INV_X1    g373(.A(new_n532), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n542), .B(new_n560), .C1(new_n546), .C2(new_n548), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G469), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n367), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT82), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n559), .B2(new_n561), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT82), .A3(new_n563), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n529), .B1(new_n558), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n446), .A2(new_n526), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n408), .A2(G221), .A3(G234), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g389(.A(KEYINPUT23), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n227), .B2(G128), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n577), .B(new_n578), .C1(G119), .C2(new_n206), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G110), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT24), .B(G110), .Z(new_n581));
  XNOR2_X1  g395(.A(G119), .B(G128), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n337), .B2(new_n349), .ZN(new_n585));
  OAI22_X1  g399(.A1(new_n579), .A2(G110), .B1(new_n582), .B2(new_n581), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n349), .A2(new_n356), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT77), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n331), .A2(new_n332), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n334), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(G146), .B1(new_n592), .B2(new_n324), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n202), .B(new_n323), .C1(new_n590), .C2(new_n591), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n583), .B(new_n580), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT77), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n587), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n575), .B1(new_n589), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n575), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n595), .B2(new_n587), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n367), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT25), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT25), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n603), .B(new_n367), .C1(new_n598), .C2(new_n600), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n377), .B1(G234), .B2(new_n367), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n598), .A2(new_n600), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n605), .A2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT78), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  OR3_X1    g424(.A1(new_n607), .A2(KEYINPUT78), .A3(new_n609), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n318), .A2(new_n572), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  INV_X1    g429(.A(new_n312), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT73), .B1(new_n311), .B2(new_n294), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n314), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n307), .B2(new_n312), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n187), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n570), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n612), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT97), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n368), .B1(new_n443), .B2(new_n445), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n401), .A2(KEYINPUT33), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n378), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT98), .B1(new_n389), .B2(new_n397), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n629), .A2(new_n630), .B1(new_n400), .B2(KEYINPUT99), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n627), .B1(new_n632), .B2(KEYINPUT33), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n370), .A2(G902), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n414), .A2(G902), .ZN(new_n636));
  OAI22_X1  g450(.A1(new_n633), .A2(new_n635), .B1(G478), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n626), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n639), .A2(new_n526), .A3(new_n413), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n625), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND2_X1  g457(.A1(new_n406), .A2(new_n416), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n526), .A2(new_n626), .A3(new_n413), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n625), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n589), .A2(new_n597), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n649), .A2(KEYINPUT36), .A3(new_n599), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n599), .A2(KEYINPUT36), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n589), .B2(new_n597), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n608), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n606), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n654), .B(new_n618), .C1(new_n619), .C2(new_n187), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n572), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT37), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  NAND2_X1  g475(.A1(new_n618), .A2(KEYINPUT32), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n313), .A2(new_n293), .A3(new_n314), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n291), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n368), .ZN(new_n665));
  INV_X1    g479(.A(new_n445), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n437), .A2(new_n363), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT93), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n365), .A3(new_n439), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n444), .B1(new_n669), .B2(new_n418), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n665), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n644), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n409), .B(KEYINPUT101), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n673), .B1(G900), .B2(new_n412), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n671), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n570), .A3(new_n526), .A4(new_n654), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n664), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT102), .B(G128), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G30));
  XNOR2_X1  g494(.A(new_n674), .B(KEYINPUT39), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n570), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT104), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n287), .A2(new_n281), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n308), .ZN(new_n687));
  AOI21_X1  g501(.A(G902), .B1(new_n687), .B2(KEYINPUT103), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(KEYINPUT103), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G472), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n315), .B2(new_n317), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n524), .A2(new_n525), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT38), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT38), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n672), .A2(new_n448), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n671), .A2(new_n699), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n692), .A2(new_n698), .A3(new_n654), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n683), .A2(new_n684), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n685), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n204), .ZN(G45));
  NOR3_X1   g518(.A1(new_n626), .A2(new_n638), .A3(new_n675), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n570), .A3(new_n526), .A4(new_n654), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n664), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n202), .ZN(G48));
  INV_X1    g522(.A(new_n567), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n566), .A2(new_n568), .B1(G469), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  INV_X1    g525(.A(new_n529), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n709), .A2(G469), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n567), .A2(KEYINPUT82), .A3(new_n563), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT82), .B1(new_n567), .B2(new_n563), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n712), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT105), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n612), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n318), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n640), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT106), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n722), .B(new_n724), .ZN(G15));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n645), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  AND4_X1   g541(.A1(new_n526), .A2(new_n713), .A3(new_n654), .A4(new_n718), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n318), .A3(new_n446), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  OAI21_X1  g544(.A(new_n311), .B1(new_n274), .B2(new_n288), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n314), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n619), .B2(new_n187), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n612), .ZN(new_n734));
  INV_X1    g548(.A(new_n719), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n693), .A2(new_n671), .A3(new_n413), .A4(new_n699), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NAND2_X1  g552(.A1(new_n313), .A2(new_n367), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n739), .A2(G472), .B1(new_n314), .B2(new_n731), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n728), .A2(new_n705), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  NOR2_X1   g556(.A1(new_n664), .A2(new_n612), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n524), .A2(new_n447), .A3(new_n525), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n570), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n743), .A2(KEYINPUT42), .A3(new_n705), .A4(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n318), .A2(new_n746), .A3(new_n613), .A4(new_n705), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  AND3_X1   g566(.A1(new_n676), .A2(new_n570), .A3(new_n744), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n318), .A3(new_n613), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT107), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n753), .A2(new_n756), .A3(new_n318), .A4(new_n613), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  OAI211_X1 g573(.A(new_n665), .B(new_n637), .C1(new_n666), .C2(new_n670), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT43), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n626), .A2(new_n762), .A3(new_n637), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n620), .A2(new_n654), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n552), .ZN(new_n767));
  INV_X1    g581(.A(new_n535), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n479), .A2(new_n471), .B1(new_n207), .B2(new_n211), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n222), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n547), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n545), .A2(KEYINPUT12), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n551), .B1(new_n773), .B2(new_n542), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n533), .B1(new_n767), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n556), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(KEYINPUT45), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n553), .B2(new_n556), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n779), .A3(G469), .ZN(new_n780));
  NAND2_X1  g594(.A1(G469), .A2(G902), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n781), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n569), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n712), .A3(new_n681), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n766), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n764), .A2(new_n765), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n744), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  NAND4_X1  g605(.A1(new_n664), .A2(new_n612), .A3(new_n705), .A4(new_n744), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n786), .A2(new_n712), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n786), .B2(new_n712), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n792), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  AND3_X1   g613(.A1(new_n654), .A2(new_n526), .A3(new_n570), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n318), .B(new_n800), .C1(new_n676), .C2(new_n705), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n606), .A2(new_n653), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n570), .A3(KEYINPUT111), .A4(new_n674), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  AOI21_X1  g618(.A(G902), .B1(new_n775), .B2(new_n776), .ZN(new_n805));
  OAI22_X1  g619(.A1(new_n805), .A2(new_n563), .B1(new_n715), .B2(new_n716), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n712), .A3(new_n674), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n804), .B1(new_n807), .B2(new_n654), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n694), .A2(new_n700), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n691), .A2(new_n803), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n801), .A2(new_n810), .A3(new_n741), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n801), .A2(new_n810), .A3(new_n741), .A4(KEYINPUT52), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT113), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n813), .A2(new_n817), .A3(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n621), .A2(new_n640), .A3(new_n623), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n614), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n614), .B2(new_n820), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n415), .A2(new_n404), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n526), .A2(new_n626), .A3(new_n413), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n621), .A2(new_n825), .A3(new_n623), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n657), .B2(new_n658), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n822), .A2(new_n823), .A3(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n720), .B(new_n318), .C1(new_n645), .C2(new_n640), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n729), .A3(new_n737), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n755), .B2(new_n757), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n740), .A2(new_n705), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n626), .A2(new_n415), .A3(new_n404), .A4(new_n674), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n664), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n745), .A2(new_n802), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n747), .A2(new_n750), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n828), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n819), .A2(new_n837), .A3(KEYINPUT53), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n664), .B1(new_n677), .B2(new_n706), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n654), .A2(new_n713), .A3(new_n718), .A4(new_n526), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n832), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT52), .A4(new_n810), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n828), .A2(new_n831), .A3(new_n845), .A4(new_n836), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n813), .A2(KEYINPUT112), .A3(new_n814), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n839), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n838), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n851));
  INV_X1    g665(.A(new_n673), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n761), .A2(new_n852), .A3(new_n763), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT114), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n761), .A2(new_n763), .A3(new_n855), .A4(new_n852), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n744), .A2(new_n713), .A3(new_n718), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT116), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n861), .B(new_n858), .C1(new_n854), .C2(new_n856), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n743), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT118), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n865), .B(new_n743), .C1(new_n860), .C2(new_n862), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(KEYINPUT48), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT48), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n863), .A2(KEYINPUT118), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n733), .A2(new_n719), .A3(new_n612), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n447), .B1(new_n695), .B2(new_n697), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n857), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(KEYINPUT50), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n876), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n857), .A2(new_n872), .A3(new_n878), .A4(new_n873), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n612), .A2(new_n409), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n671), .A2(new_n637), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n692), .A2(new_n859), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n710), .A2(new_n529), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n795), .B2(new_n797), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n734), .A2(new_n744), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n856), .B2(new_n854), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n740), .A2(new_n654), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n860), .B2(new_n862), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n880), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n885), .A2(new_n887), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n883), .A2(new_n893), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n880), .A2(new_n891), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n692), .A2(new_n859), .A3(new_n881), .ZN(new_n898));
  INV_X1    g712(.A(new_n639), .ZN(new_n899));
  OAI211_X1 g713(.A(G952), .B(new_n408), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n857), .A2(new_n526), .A3(new_n872), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT117), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(KEYINPUT117), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n870), .A2(new_n871), .A3(new_n894), .A4(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n813), .A2(new_n817), .A3(new_n814), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n817), .B1(new_n813), .B2(new_n814), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n828), .A2(new_n831), .A3(new_n836), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n839), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n837), .A2(KEYINPUT53), .A3(new_n847), .A4(new_n845), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n894), .A2(new_n897), .A3(new_n904), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n867), .A2(new_n869), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT119), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n851), .A2(new_n906), .A3(new_n914), .A4(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(G952), .A2(G953), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n760), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n613), .A2(new_n712), .A3(new_n447), .A4(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(KEYINPUT109), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(KEYINPUT109), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n710), .B(KEYINPUT49), .Z(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n695), .B2(new_n697), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n923), .A2(new_n692), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT120), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n920), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(G75));
  NOR2_X1   g746(.A1(new_n408), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n367), .B1(new_n911), .B2(new_n913), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(G210), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n497), .A2(new_n499), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n489), .B2(new_n497), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n462), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT55), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n934), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n936), .B2(new_n941), .ZN(G51));
  INV_X1    g757(.A(new_n780), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT53), .B1(new_n819), .B2(new_n837), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n846), .A2(new_n839), .A3(new_n848), .ZN(new_n946));
  OAI211_X1 g760(.A(G902), .B(new_n944), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n781), .B(KEYINPUT57), .Z(new_n949));
  NOR3_X1   g763(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT54), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n948), .B1(new_n952), .B2(new_n562), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT121), .B1(new_n953), .B2(new_n933), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT121), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT54), .B1(new_n945), .B2(new_n946), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n914), .ZN(new_n957));
  AOI22_X1  g771(.A1(new_n957), .A2(new_n949), .B1(new_n559), .B2(new_n561), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n955), .B(new_n934), .C1(new_n958), .C2(new_n948), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n954), .A2(new_n959), .ZN(G54));
  NAND3_X1  g774(.A1(new_n935), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  INV_X1    g775(.A(new_n669), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n933), .ZN(G60));
  XOR2_X1   g779(.A(new_n633), .B(KEYINPUT122), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n851), .A2(new_n914), .ZN(new_n967));
  NAND2_X1  g781(.A1(G478), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT59), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n966), .A2(new_n969), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n933), .B(new_n970), .C1(new_n957), .C2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(new_n911), .A2(new_n913), .ZN(new_n973));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT60), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n607), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n973), .B(new_n975), .C1(new_n650), .C2(new_n652), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n934), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G66));
  INV_X1    g795(.A(new_n830), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n828), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n408), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT123), .Z(new_n985));
  AOI21_X1  g799(.A(new_n408), .B1(new_n411), .B2(G224), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT124), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT125), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n985), .A2(new_n990), .A3(new_n987), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(G898), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n938), .B1(new_n993), .B2(G953), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n992), .B(new_n994), .ZN(G69));
  NAND2_X1  g809(.A1(new_n225), .A2(new_n255), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n432), .A2(new_n420), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n996), .B(new_n997), .Z(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(G900), .B2(G953), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n743), .A2(new_n809), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n843), .B1(new_n787), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(new_n750), .B2(new_n747), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1002), .A2(new_n790), .A3(new_n758), .A4(new_n798), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n999), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n843), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n703), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT62), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n626), .A2(new_n824), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n899), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n743), .A2(new_n683), .A3(new_n744), .A4(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1009), .A2(new_n790), .A3(new_n798), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n408), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n998), .B(KEYINPUT126), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1006), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n408), .B1(G227), .B2(G900), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1016), .B(new_n1018), .ZN(G72));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT63), .Z(new_n1021));
  OAI21_X1  g835(.A(new_n1021), .B1(new_n1013), .B2(new_n983), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1022), .A2(new_n274), .A3(new_n259), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n308), .B1(new_n260), .B2(new_n274), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n850), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1021), .B1(new_n1003), .B2(new_n983), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n281), .A3(new_n260), .ZN(new_n1027));
  AND4_X1   g841(.A1(new_n934), .A2(new_n1023), .A3(new_n1025), .A4(new_n1027), .ZN(G57));
endmodule


