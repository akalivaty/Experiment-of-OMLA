

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752;

  NAND2_X1 U362 ( .A1(n340), .A2(n435), .ZN(n655) );
  AND2_X1 U363 ( .A1(n432), .A2(n433), .ZN(n340) );
  OR2_X2 U364 ( .A1(n631), .A2(G902), .ZN(n391) );
  XNOR2_X2 U365 ( .A(n431), .B(G122), .ZN(n471) );
  XNOR2_X2 U366 ( .A(G116), .B(G107), .ZN(n431) );
  XNOR2_X2 U367 ( .A(n342), .B(KEYINPUT4), .ZN(n737) );
  XNOR2_X2 U368 ( .A(KEYINPUT64), .B(KEYINPUT70), .ZN(n342) );
  XNOR2_X2 U369 ( .A(n344), .B(n345), .ZN(n546) );
  AND2_X1 U370 ( .A1(n367), .A2(n368), .ZN(n366) );
  XNOR2_X1 U371 ( .A(n364), .B(n427), .ZN(n583) );
  OR2_X1 U372 ( .A1(n612), .A2(n664), .ZN(n354) );
  OR2_X1 U373 ( .A1(n574), .A2(n353), .ZN(n435) );
  XNOR2_X1 U374 ( .A(n498), .B(n497), .ZN(n536) );
  XNOR2_X1 U375 ( .A(n380), .B(n564), .ZN(n574) );
  XNOR2_X1 U376 ( .A(n341), .B(KEYINPUT111), .ZN(n535) );
  AND2_X1 U377 ( .A1(n400), .A2(n399), .ZN(n398) );
  XNOR2_X1 U378 ( .A(n538), .B(KEYINPUT106), .ZN(n665) );
  AND2_X1 U379 ( .A1(n426), .A2(n425), .ZN(n424) );
  XNOR2_X1 U380 ( .A(n493), .B(KEYINPUT95), .ZN(n494) );
  XNOR2_X1 U381 ( .A(n527), .B(n526), .ZN(n649) );
  XNOR2_X1 U382 ( .A(n525), .B(n524), .ZN(n527) );
  NAND2_X1 U383 ( .A1(n548), .A2(n532), .ZN(n341) );
  XNOR2_X2 U384 ( .A(n682), .B(KEYINPUT91), .ZN(n548) );
  XNOR2_X2 U385 ( .A(n607), .B(KEYINPUT1), .ZN(n682) );
  NAND2_X1 U386 ( .A1(n398), .A2(n395), .ZN(n343) );
  NAND2_X1 U387 ( .A1(n398), .A2(n395), .ZN(n610) );
  NOR2_X1 U388 ( .A1(n638), .A2(n482), .ZN(n344) );
  XOR2_X1 U389 ( .A(n486), .B(n485), .Z(n345) );
  INV_X1 U390 ( .A(KEYINPUT76), .ZN(n412) );
  AND2_X1 U391 ( .A1(n372), .A2(n672), .ZN(n369) );
  NOR2_X1 U392 ( .A1(n750), .A2(n751), .ZN(n407) );
  XNOR2_X1 U393 ( .A(n447), .B(n446), .ZN(n738) );
  XNOR2_X1 U394 ( .A(n477), .B(G140), .ZN(n446) );
  XOR2_X1 U395 ( .A(G104), .B(G122), .Z(n452) );
  XNOR2_X1 U396 ( .A(KEYINPUT73), .B(G131), .ZN(n499) );
  NAND2_X1 U397 ( .A1(n676), .A2(KEYINPUT19), .ZN(n399) );
  NOR2_X1 U398 ( .A1(G237), .A2(G953), .ZN(n453) );
  NAND2_X1 U399 ( .A1(n578), .A2(n577), .ZN(n420) );
  INV_X1 U400 ( .A(KEYINPUT44), .ZN(n363) );
  INV_X1 U401 ( .A(KEYINPUT84), .ZN(n582) );
  NAND2_X2 U402 ( .A1(n424), .A2(n421), .ZN(n607) );
  XNOR2_X1 U403 ( .A(G128), .B(G119), .ZN(n512) );
  XOR2_X1 U404 ( .A(KEYINPUT23), .B(G110), .Z(n513) );
  XNOR2_X1 U405 ( .A(n740), .B(G146), .ZN(n526) );
  NAND2_X1 U406 ( .A1(n346), .A2(n357), .ZN(n741) );
  INV_X1 U407 ( .A(KEYINPUT2), .ZN(n379) );
  BUF_X1 U408 ( .A(n607), .Z(n402) );
  XNOR2_X1 U409 ( .A(KEYINPUT116), .B(KEYINPUT28), .ZN(n605) );
  XNOR2_X1 U410 ( .A(n392), .B(KEYINPUT39), .ZN(n626) );
  NOR2_X1 U411 ( .A1(n665), .A2(n602), .ZN(n544) );
  XNOR2_X1 U412 ( .A(n575), .B(KEYINPUT34), .ZN(n429) );
  NOR2_X1 U413 ( .A1(n361), .A2(n574), .ZN(n575) );
  BUF_X1 U414 ( .A(n546), .Z(n623) );
  XNOR2_X1 U415 ( .A(n459), .B(n458), .ZN(n620) );
  XNOR2_X1 U416 ( .A(n457), .B(n456), .ZN(n458) );
  INV_X1 U417 ( .A(G475), .ZN(n456) );
  XNOR2_X1 U418 ( .A(n520), .B(n519), .ZN(n404) );
  XNOR2_X1 U419 ( .A(KEYINPUT97), .B(KEYINPUT25), .ZN(n519) );
  XNOR2_X1 U420 ( .A(n465), .B(G478), .ZN(n616) );
  XNOR2_X1 U421 ( .A(n635), .B(KEYINPUT92), .ZN(n714) );
  OR2_X1 U422 ( .A1(n661), .A2(KEYINPUT47), .ZN(n612) );
  INV_X1 U423 ( .A(KEYINPUT102), .ZN(n394) );
  NAND2_X1 U424 ( .A1(n668), .A2(n665), .ZN(n672) );
  NOR2_X1 U425 ( .A1(n410), .A2(n598), .ZN(n673) );
  INV_X1 U426 ( .A(n672), .ZN(n410) );
  INV_X1 U427 ( .A(G237), .ZN(n483) );
  NAND2_X1 U428 ( .A1(n423), .A2(n484), .ZN(n422) );
  XNOR2_X1 U429 ( .A(n381), .B(G119), .ZN(n502) );
  XNOR2_X1 U430 ( .A(G113), .B(KEYINPUT3), .ZN(n381) );
  XNOR2_X1 U431 ( .A(G143), .B(G113), .ZN(n451) );
  XNOR2_X1 U432 ( .A(n499), .B(G137), .ZN(n500) );
  XNOR2_X1 U433 ( .A(n445), .B(G125), .ZN(n477) );
  INV_X1 U434 ( .A(G146), .ZN(n445) );
  XOR2_X1 U435 ( .A(KEYINPUT80), .B(KEYINPUT17), .Z(n475) );
  NAND2_X1 U436 ( .A1(G234), .A2(G237), .ZN(n488) );
  NOR2_X1 U437 ( .A1(n671), .A2(n598), .ZN(n678) );
  XNOR2_X1 U438 ( .A(n623), .B(n409), .ZN(n598) );
  INV_X1 U439 ( .A(KEYINPUT38), .ZN(n409) );
  NAND2_X1 U440 ( .A1(n397), .A2(n396), .ZN(n395) );
  NOR2_X1 U441 ( .A1(n676), .A2(KEYINPUT19), .ZN(n396) );
  NOR2_X1 U442 ( .A1(n594), .A2(KEYINPUT99), .ZN(n434) );
  INV_X1 U443 ( .A(KEYINPUT99), .ZN(n436) );
  NOR2_X1 U444 ( .A1(n671), .A2(n469), .ZN(n470) );
  XNOR2_X1 U445 ( .A(n502), .B(n441), .ZN(n505) );
  XNOR2_X1 U446 ( .A(n443), .B(n442), .ZN(n441) );
  XNOR2_X1 U447 ( .A(KEYINPUT100), .B(G116), .ZN(n443) );
  XNOR2_X1 U448 ( .A(KEYINPUT5), .B(KEYINPUT77), .ZN(n442) );
  XNOR2_X1 U449 ( .A(n737), .B(n360), .ZN(n506) );
  XNOR2_X1 U450 ( .A(n419), .B(KEYINPUT67), .ZN(n360) );
  XNOR2_X1 U451 ( .A(KEYINPUT68), .B(G101), .ZN(n419) );
  XNOR2_X1 U452 ( .A(n430), .B(n502), .ZN(n723) );
  XNOR2_X1 U453 ( .A(n471), .B(KEYINPUT16), .ZN(n430) );
  XNOR2_X1 U454 ( .A(n573), .B(n572), .ZN(n361) );
  XNOR2_X1 U455 ( .A(n563), .B(n562), .ZN(n437) );
  XNOR2_X1 U456 ( .A(n689), .B(KEYINPUT112), .ZN(n603) );
  XNOR2_X1 U457 ( .A(n566), .B(n418), .ZN(n625) );
  INV_X1 U458 ( .A(KEYINPUT107), .ZN(n418) );
  XNOR2_X1 U459 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U460 ( .A(n515), .B(n514), .ZN(n517) );
  XOR2_X1 U461 ( .A(n708), .B(n707), .Z(n709) );
  XNOR2_X1 U462 ( .A(n639), .B(n642), .ZN(n643) );
  NAND2_X1 U463 ( .A1(n375), .A2(n374), .ZN(n373) );
  NOR2_X1 U464 ( .A1(n741), .A2(n379), .ZN(n374) );
  AND2_X1 U465 ( .A1(n378), .A2(n377), .ZN(n376) );
  INV_X2 U466 ( .A(G953), .ZN(n742) );
  XNOR2_X1 U467 ( .A(n408), .B(KEYINPUT42), .ZN(n751) );
  XNOR2_X1 U468 ( .A(n597), .B(n596), .ZN(n750) );
  NOR2_X1 U469 ( .A1(n553), .A2(n623), .ZN(n547) );
  INV_X1 U470 ( .A(KEYINPUT35), .ZN(n427) );
  NAND2_X1 U471 ( .A1(n429), .A2(n356), .ZN(n364) );
  INV_X1 U472 ( .A(KEYINPUT32), .ZN(n388) );
  NOR2_X1 U473 ( .A1(n624), .A2(n623), .ZN(n662) );
  AND2_X1 U474 ( .A1(n613), .A2(n625), .ZN(n661) );
  XNOR2_X1 U475 ( .A(n371), .B(n370), .ZN(n567) );
  INV_X1 U476 ( .A(KEYINPUT109), .ZN(n370) );
  OR2_X1 U477 ( .A1(n536), .A2(n350), .ZN(n371) );
  XNOR2_X1 U478 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U479 ( .A(n717), .B(n716), .ZN(n405) );
  XNOR2_X1 U480 ( .A(n649), .B(n648), .ZN(n650) );
  OR2_X1 U481 ( .A1(n402), .A2(n681), .ZN(n593) );
  AND2_X1 U482 ( .A1(n385), .A2(n382), .ZN(n346) );
  OR2_X1 U483 ( .A1(n615), .A2(n614), .ZN(n347) );
  OR2_X1 U484 ( .A1(G902), .A2(n719), .ZN(n348) );
  XOR2_X1 U485 ( .A(n450), .B(n449), .Z(n349) );
  OR2_X1 U486 ( .A1(n537), .A2(n560), .ZN(n350) );
  AND2_X1 U487 ( .A1(n376), .A2(n373), .ZN(n351) );
  AND2_X1 U488 ( .A1(n667), .A2(KEYINPUT102), .ZN(n352) );
  OR2_X1 U489 ( .A1(n593), .A2(n436), .ZN(n353) );
  AND2_X1 U490 ( .A1(n435), .A2(n394), .ZN(n355) );
  AND2_X1 U491 ( .A1(n576), .A2(n428), .ZN(n356) );
  AND2_X1 U492 ( .A1(n670), .A2(n627), .ZN(n357) );
  NOR2_X1 U493 ( .A1(n679), .A2(n361), .ZN(n358) );
  XNOR2_X1 U494 ( .A(n518), .B(n738), .ZN(n719) );
  XNOR2_X1 U495 ( .A(n359), .B(n582), .ZN(n588) );
  NAND2_X1 U496 ( .A1(n580), .A2(n581), .ZN(n359) );
  AND2_X2 U497 ( .A1(n373), .A2(n482), .ZN(n362) );
  NAND2_X1 U498 ( .A1(n549), .A2(n548), .ZN(n440) );
  NOR2_X1 U499 ( .A1(n439), .A2(KEYINPUT48), .ZN(n387) );
  XNOR2_X2 U500 ( .A(n506), .B(n724), .ZN(n525) );
  NOR2_X1 U501 ( .A1(n699), .A2(n361), .ZN(n700) );
  AND2_X4 U502 ( .A1(n362), .A2(n376), .ZN(n715) );
  INV_X1 U503 ( .A(n583), .ZN(n749) );
  NAND2_X1 U504 ( .A1(n583), .A2(n363), .ZN(n584) );
  NAND2_X1 U505 ( .A1(n365), .A2(n567), .ZN(n569) );
  NAND2_X1 U506 ( .A1(n366), .A2(n369), .ZN(n365) );
  NAND2_X1 U507 ( .A1(n352), .A2(n655), .ZN(n367) );
  NAND2_X1 U508 ( .A1(n355), .A2(n340), .ZN(n368) );
  NAND2_X1 U509 ( .A1(n393), .A2(n394), .ZN(n372) );
  INV_X1 U510 ( .A(n728), .ZN(n375) );
  NAND2_X1 U511 ( .A1(n741), .A2(n379), .ZN(n377) );
  NAND2_X1 U512 ( .A1(n728), .A2(n379), .ZN(n378) );
  XNOR2_X2 U513 ( .A(n590), .B(n589), .ZN(n728) );
  AND2_X2 U514 ( .A1(n380), .A2(n496), .ZN(n498) );
  AND2_X1 U515 ( .A1(n380), .A2(n689), .ZN(n561) );
  XNOR2_X2 U516 ( .A(n401), .B(n495), .ZN(n380) );
  NAND2_X1 U517 ( .A1(n383), .A2(KEYINPUT48), .ZN(n382) );
  NAND2_X1 U518 ( .A1(n386), .A2(n384), .ZN(n383) );
  INV_X1 U519 ( .A(n439), .ZN(n384) );
  NAND2_X1 U520 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U521 ( .A(n407), .B(KEYINPUT46), .ZN(n386) );
  XNOR2_X2 U522 ( .A(n389), .B(n388), .ZN(n578) );
  NOR2_X2 U523 ( .A1(n536), .A2(n390), .ZN(n389) );
  NAND2_X1 U524 ( .A1(n535), .A2(n534), .ZN(n390) );
  NAND2_X1 U525 ( .A1(n603), .A2(n599), .ZN(n591) );
  XNOR2_X2 U526 ( .A(n391), .B(G472), .ZN(n689) );
  NAND2_X1 U527 ( .A1(n618), .A2(n595), .ZN(n392) );
  NOR2_X2 U528 ( .A1(n592), .A2(n593), .ZN(n618) );
  INV_X1 U529 ( .A(n667), .ZN(n393) );
  INV_X1 U530 ( .A(n546), .ZN(n397) );
  NAND2_X1 U531 ( .A1(n546), .A2(KEYINPUT19), .ZN(n400) );
  NAND2_X1 U532 ( .A1(n610), .A2(n494), .ZN(n401) );
  XNOR2_X1 U533 ( .A(n403), .B(n501), .ZN(n464) );
  XNOR2_X1 U534 ( .A(n471), .B(n460), .ZN(n403) );
  NOR2_X1 U535 ( .A1(n434), .A2(n689), .ZN(n433) );
  XNOR2_X2 U536 ( .A(n348), .B(n404), .ZN(n558) );
  XNOR2_X1 U537 ( .A(n413), .B(n412), .ZN(n411) );
  NAND2_X1 U538 ( .A1(n585), .A2(n583), .ZN(n579) );
  XNOR2_X2 U539 ( .A(n420), .B(KEYINPUT85), .ZN(n585) );
  NOR2_X1 U540 ( .A1(n405), .A2(n722), .ZN(G63) );
  XNOR2_X1 U541 ( .A(n406), .B(n349), .ZN(n708) );
  XNOR2_X1 U542 ( .A(n455), .B(n738), .ZN(n406) );
  NAND2_X1 U543 ( .A1(n415), .A2(n414), .ZN(n413) );
  AND2_X1 U544 ( .A1(n680), .A2(n609), .ZN(n408) );
  NAND2_X1 U545 ( .A1(n411), .A2(n440), .ZN(n439) );
  INV_X1 U546 ( .A(n662), .ZN(n414) );
  NAND2_X1 U547 ( .A1(n354), .A2(n347), .ZN(n415) );
  NOR2_X1 U548 ( .A1(n608), .A2(n416), .ZN(n613) );
  NOR2_X1 U549 ( .A1(n608), .A2(n402), .ZN(n609) );
  NAND2_X1 U550 ( .A1(n343), .A2(n417), .ZN(n416) );
  INV_X1 U551 ( .A(n402), .ZN(n417) );
  INV_X1 U552 ( .A(n625), .ZN(n668) );
  NAND2_X1 U553 ( .A1(n649), .A2(n529), .ZN(n426) );
  OR2_X1 U554 ( .A1(n649), .A2(n422), .ZN(n421) );
  INV_X1 U555 ( .A(n529), .ZN(n423) );
  NAND2_X1 U556 ( .A1(n529), .A2(G902), .ZN(n425) );
  INV_X1 U557 ( .A(n616), .ZN(n428) );
  NAND2_X1 U558 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U559 ( .A1(n574), .A2(n436), .ZN(n432) );
  XNOR2_X2 U560 ( .A(n438), .B(n437), .ZN(n667) );
  NAND2_X1 U561 ( .A1(n561), .A2(n690), .ZN(n438) );
  XNOR2_X1 U562 ( .A(n509), .B(n526), .ZN(n631) );
  XNOR2_X1 U563 ( .A(n606), .B(n605), .ZN(n608) );
  BUF_X1 U564 ( .A(n715), .Z(n718) );
  XOR2_X1 U565 ( .A(n452), .B(n451), .Z(n444) );
  INV_X1 U566 ( .A(KEYINPUT110), .ZN(n568) );
  INV_X1 U567 ( .A(n682), .ZN(n560) );
  INV_X1 U568 ( .A(KEYINPUT96), .ZN(n564) );
  XNOR2_X1 U569 ( .A(n444), .B(n454), .ZN(n455) );
  XNOR2_X1 U570 ( .A(n501), .B(n500), .ZN(n740) );
  INV_X1 U571 ( .A(KEYINPUT101), .ZN(n562) );
  INV_X1 U572 ( .A(KEYINPUT40), .ZN(n596) );
  XOR2_X1 U573 ( .A(KEYINPUT10), .B(KEYINPUT72), .Z(n447) );
  XOR2_X1 U574 ( .A(KEYINPUT103), .B(KEYINPUT12), .Z(n450) );
  INV_X1 U575 ( .A(n499), .ZN(n448) );
  XNOR2_X1 U576 ( .A(n448), .B(KEYINPUT11), .ZN(n449) );
  XNOR2_X1 U577 ( .A(n453), .B(KEYINPUT78), .ZN(n503) );
  NAND2_X1 U578 ( .A1(G214), .A2(n503), .ZN(n454) );
  NOR2_X1 U579 ( .A1(G902), .A2(n708), .ZN(n459) );
  XNOR2_X1 U580 ( .A(KEYINPUT13), .B(KEYINPUT104), .ZN(n457) );
  XOR2_X1 U581 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n460) );
  XNOR2_X2 U582 ( .A(G143), .B(G128), .ZN(n476) );
  XNOR2_X1 U583 ( .A(G134), .B(n476), .ZN(n501) );
  NAND2_X1 U584 ( .A1(n742), .A2(G234), .ZN(n462) );
  XNOR2_X1 U585 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n461) );
  XNOR2_X1 U586 ( .A(n462), .B(n461), .ZN(n511) );
  NAND2_X1 U587 ( .A1(n511), .A2(G217), .ZN(n463) );
  XOR2_X1 U588 ( .A(n464), .B(n463), .Z(n716) );
  NOR2_X1 U589 ( .A1(n716), .A2(G902), .ZN(n465) );
  NAND2_X1 U590 ( .A1(n620), .A2(n616), .ZN(n671) );
  XNOR2_X1 U591 ( .A(KEYINPUT15), .B(G902), .ZN(n628) );
  NAND2_X1 U592 ( .A1(n628), .A2(G234), .ZN(n467) );
  XNOR2_X1 U593 ( .A(KEYINPUT98), .B(KEYINPUT20), .ZN(n466) );
  XNOR2_X1 U594 ( .A(n467), .B(n466), .ZN(n510) );
  NAND2_X1 U595 ( .A1(n510), .A2(G221), .ZN(n468) );
  XOR2_X1 U596 ( .A(KEYINPUT21), .B(n468), .Z(n684) );
  INV_X1 U597 ( .A(n684), .ZN(n469) );
  XNOR2_X1 U598 ( .A(n470), .B(KEYINPUT108), .ZN(n496) );
  NAND2_X1 U599 ( .A1(G224), .A2(n742), .ZN(n473) );
  XNOR2_X1 U600 ( .A(KEYINPUT89), .B(KEYINPUT18), .ZN(n472) );
  XNOR2_X1 U601 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U602 ( .A(n475), .B(n474), .ZN(n479) );
  XNOR2_X1 U603 ( .A(n476), .B(n477), .ZN(n478) );
  XNOR2_X1 U604 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U605 ( .A(n723), .B(n480), .ZN(n481) );
  XNOR2_X1 U606 ( .A(G110), .B(G104), .ZN(n724) );
  XNOR2_X1 U607 ( .A(n481), .B(n525), .ZN(n638) );
  INV_X1 U608 ( .A(n628), .ZN(n482) );
  INV_X1 U609 ( .A(G902), .ZN(n484) );
  NAND2_X1 U610 ( .A1(n484), .A2(n483), .ZN(n487) );
  NAND2_X1 U611 ( .A1(n487), .A2(G210), .ZN(n486) );
  INV_X1 U612 ( .A(KEYINPUT93), .ZN(n485) );
  NAND2_X1 U613 ( .A1(n487), .A2(G214), .ZN(n599) );
  INV_X1 U614 ( .A(n599), .ZN(n676) );
  XNOR2_X1 U615 ( .A(n488), .B(KEYINPUT14), .ZN(n490) );
  NAND2_X1 U616 ( .A1(G952), .A2(n490), .ZN(n698) );
  NOR2_X1 U617 ( .A1(n698), .A2(G953), .ZN(n489) );
  XNOR2_X1 U618 ( .A(n489), .B(KEYINPUT94), .ZN(n541) );
  AND2_X1 U619 ( .A1(G953), .A2(n490), .ZN(n491) );
  NAND2_X1 U620 ( .A1(G902), .A2(n491), .ZN(n539) );
  NOR2_X1 U621 ( .A1(G898), .A2(n539), .ZN(n492) );
  NOR2_X1 U622 ( .A1(n541), .A2(n492), .ZN(n493) );
  INV_X1 U623 ( .A(KEYINPUT0), .ZN(n495) );
  XNOR2_X1 U624 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n497) );
  NAND2_X1 U625 ( .A1(n503), .A2(G210), .ZN(n504) );
  XNOR2_X1 U626 ( .A(n505), .B(n504), .ZN(n508) );
  INV_X1 U627 ( .A(n506), .ZN(n507) );
  XNOR2_X1 U628 ( .A(n508), .B(n507), .ZN(n509) );
  NAND2_X1 U629 ( .A1(G217), .A2(n510), .ZN(n520) );
  NAND2_X1 U630 ( .A1(n511), .A2(G221), .ZN(n515) );
  XNOR2_X1 U631 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U632 ( .A(G137), .B(KEYINPUT24), .Z(n516) );
  NOR2_X1 U633 ( .A1(n603), .A2(n558), .ZN(n530) );
  NAND2_X1 U634 ( .A1(n742), .A2(G227), .ZN(n521) );
  XNOR2_X1 U635 ( .A(n521), .B(G107), .ZN(n523) );
  XNOR2_X1 U636 ( .A(KEYINPUT79), .B(G140), .ZN(n522) );
  XNOR2_X1 U637 ( .A(n523), .B(n522), .ZN(n524) );
  INV_X1 U638 ( .A(KEYINPUT74), .ZN(n528) );
  XNOR2_X1 U639 ( .A(n528), .B(G469), .ZN(n529) );
  NAND2_X1 U640 ( .A1(n530), .A2(n682), .ZN(n531) );
  OR2_X1 U641 ( .A1(n536), .A2(n531), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G110), .ZN(G12) );
  INV_X1 U643 ( .A(n558), .ZN(n532) );
  XNOR2_X1 U644 ( .A(n689), .B(KEYINPUT6), .ZN(n570) );
  INV_X1 U645 ( .A(n570), .ZN(n533) );
  XNOR2_X1 U646 ( .A(n533), .B(KEYINPUT81), .ZN(n534) );
  XNOR2_X1 U647 ( .A(n578), .B(G119), .ZN(G21) );
  NAND2_X1 U648 ( .A1(n570), .A2(n558), .ZN(n537) );
  XNOR2_X1 U649 ( .A(n567), .B(G101), .ZN(G3) );
  XNOR2_X1 U650 ( .A(n620), .B(KEYINPUT105), .ZN(n565) );
  NAND2_X1 U651 ( .A1(n565), .A2(n616), .ZN(n538) );
  XOR2_X1 U652 ( .A(KEYINPUT113), .B(n539), .Z(n540) );
  NOR2_X1 U653 ( .A1(G900), .A2(n540), .ZN(n542) );
  NOR2_X1 U654 ( .A1(n542), .A2(n541), .ZN(n617) );
  NOR2_X1 U655 ( .A1(n617), .A2(n558), .ZN(n543) );
  NAND2_X1 U656 ( .A1(n543), .A2(n684), .ZN(n602) );
  NAND2_X1 U657 ( .A1(n544), .A2(n599), .ZN(n545) );
  OR2_X1 U658 ( .A1(n545), .A2(n570), .ZN(n553) );
  XNOR2_X1 U659 ( .A(n547), .B(KEYINPUT36), .ZN(n549) );
  XOR2_X1 U660 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n551) );
  XNOR2_X1 U661 ( .A(G125), .B(KEYINPUT37), .ZN(n550) );
  XNOR2_X1 U662 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U663 ( .A(n440), .B(n552), .Z(G27) );
  XOR2_X1 U664 ( .A(n553), .B(KEYINPUT114), .Z(n554) );
  AND2_X1 U665 ( .A1(n554), .A2(n682), .ZN(n556) );
  XNOR2_X1 U666 ( .A(KEYINPUT115), .B(KEYINPUT43), .ZN(n555) );
  XNOR2_X1 U667 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U668 ( .A1(n557), .A2(n623), .ZN(n627) );
  XNOR2_X1 U669 ( .A(n627), .B(G140), .ZN(G42) );
  INV_X1 U670 ( .A(KEYINPUT31), .ZN(n563) );
  NAND2_X1 U671 ( .A1(n684), .A2(n558), .ZN(n681) );
  INV_X1 U672 ( .A(n681), .ZN(n559) );
  NAND2_X1 U673 ( .A1(n560), .A2(n559), .ZN(n571) );
  INV_X1 U674 ( .A(n571), .ZN(n690) );
  NOR2_X1 U675 ( .A1(n565), .A2(n616), .ZN(n566) );
  XNOR2_X1 U676 ( .A(n569), .B(n568), .ZN(n581) );
  NOR2_X1 U677 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U678 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n572) );
  INV_X1 U679 ( .A(n620), .ZN(n576) );
  NAND2_X1 U680 ( .A1(n579), .A2(KEYINPUT44), .ZN(n580) );
  XNOR2_X1 U681 ( .A(KEYINPUT69), .B(n584), .ZN(n586) );
  NAND2_X1 U682 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U683 ( .A(KEYINPUT82), .B(KEYINPUT45), .Z(n589) );
  XNOR2_X1 U684 ( .A(KEYINPUT30), .B(n591), .ZN(n592) );
  INV_X1 U685 ( .A(n593), .ZN(n594) );
  NOR2_X1 U686 ( .A1(n598), .A2(n617), .ZN(n595) );
  INV_X1 U687 ( .A(n665), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n626), .A2(n611), .ZN(n597) );
  XOR2_X1 U689 ( .A(KEYINPUT41), .B(KEYINPUT117), .Z(n601) );
  NAND2_X1 U690 ( .A1(n678), .A2(n599), .ZN(n600) );
  XNOR2_X1 U691 ( .A(n601), .B(n600), .ZN(n680) );
  INV_X1 U692 ( .A(n602), .ZN(n604) );
  NAND2_X1 U693 ( .A1(n604), .A2(n603), .ZN(n606) );
  AND2_X1 U694 ( .A1(n613), .A2(n611), .ZN(n664) );
  INV_X1 U695 ( .A(n613), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n672), .A2(KEYINPUT47), .ZN(n614) );
  NOR2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n622) );
  INV_X1 U698 ( .A(n618), .ZN(n619) );
  NOR2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n670) );
  NAND2_X1 U702 ( .A1(n715), .A2(G472), .ZN(n633) );
  XNOR2_X1 U703 ( .A(KEYINPUT90), .B(KEYINPUT118), .ZN(n629) );
  XOR2_X1 U704 ( .A(n629), .B(KEYINPUT62), .Z(n630) );
  XNOR2_X1 U705 ( .A(n633), .B(n632), .ZN(n636) );
  INV_X1 U706 ( .A(G952), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n634), .A2(G953), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n636), .A2(n714), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n637), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U710 ( .A1(n715), .A2(G210), .ZN(n644) );
  BUF_X1 U711 ( .A(n638), .Z(n639) );
  XOR2_X1 U712 ( .A(KEYINPUT87), .B(KEYINPUT54), .Z(n641) );
  XNOR2_X1 U713 ( .A(KEYINPUT55), .B(KEYINPUT86), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n645), .A2(n714), .ZN(n647) );
  XNOR2_X1 U717 ( .A(KEYINPUT83), .B(KEYINPUT56), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(G51) );
  NAND2_X1 U719 ( .A1(n715), .A2(G469), .ZN(n651) );
  XNOR2_X1 U720 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U722 ( .A1(n652), .A2(n714), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n653), .B(KEYINPUT123), .ZN(G54) );
  NOR2_X1 U724 ( .A1(n665), .A2(n655), .ZN(n654) );
  XOR2_X1 U725 ( .A(G104), .B(n654), .Z(G6) );
  NOR2_X1 U726 ( .A1(n655), .A2(n668), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT119), .B(KEYINPUT26), .Z(n657) );
  XNOR2_X1 U728 ( .A(G107), .B(KEYINPUT27), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n659), .B(n658), .ZN(G9) );
  XNOR2_X1 U731 ( .A(G128), .B(KEYINPUT29), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(G30) );
  XOR2_X1 U733 ( .A(G143), .B(n662), .Z(n663) );
  XNOR2_X1 U734 ( .A(KEYINPUT120), .B(n663), .ZN(G45) );
  XOR2_X1 U735 ( .A(G146), .B(n664), .Z(G48) );
  NOR2_X1 U736 ( .A1(n665), .A2(n667), .ZN(n666) );
  XOR2_X1 U737 ( .A(G113), .B(n666), .Z(G15) );
  NOR2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U739 ( .A(G116), .B(n669), .Z(G18) );
  XNOR2_X1 U740 ( .A(G134), .B(n670), .ZN(G36) );
  INV_X1 U741 ( .A(n671), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  INV_X1 U745 ( .A(n680), .ZN(n699) );
  NAND2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U747 ( .A(n683), .B(KEYINPUT50), .ZN(n688) );
  NOR2_X1 U748 ( .A1(n684), .A2(n558), .ZN(n685) );
  XOR2_X1 U749 ( .A(KEYINPUT49), .B(n685), .Z(n686) );
  NOR2_X1 U750 ( .A1(n689), .A2(n686), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U752 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U754 ( .A(KEYINPUT51), .B(n693), .ZN(n694) );
  NOR2_X1 U755 ( .A1(n699), .A2(n694), .ZN(n695) );
  NOR2_X1 U756 ( .A1(n358), .A2(n695), .ZN(n696) );
  XNOR2_X1 U757 ( .A(n696), .B(KEYINPUT52), .ZN(n697) );
  NOR2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U760 ( .A1(n702), .A2(n742), .ZN(n703) );
  NOR2_X1 U761 ( .A1(n351), .A2(n703), .ZN(n704) );
  XNOR2_X1 U762 ( .A(n704), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U763 ( .A1(n715), .A2(G475), .ZN(n710) );
  XOR2_X1 U764 ( .A(KEYINPUT65), .B(KEYINPUT125), .Z(n706) );
  XNOR2_X1 U765 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n705) );
  XNOR2_X1 U766 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U767 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U768 ( .A1(n711), .A2(n714), .ZN(n713) );
  XOR2_X1 U769 ( .A(KEYINPUT60), .B(KEYINPUT66), .Z(n712) );
  XNOR2_X1 U770 ( .A(n713), .B(n712), .ZN(G60) );
  INV_X1 U771 ( .A(n714), .ZN(n722) );
  NAND2_X1 U772 ( .A1(n718), .A2(G478), .ZN(n717) );
  NAND2_X1 U773 ( .A1(n718), .A2(G217), .ZN(n720) );
  XNOR2_X1 U774 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U775 ( .A1(n722), .A2(n721), .ZN(G66) );
  XNOR2_X1 U776 ( .A(n723), .B(G101), .ZN(n725) );
  XNOR2_X1 U777 ( .A(n725), .B(n724), .ZN(n727) );
  NOR2_X1 U778 ( .A1(G898), .A2(n742), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n736) );
  NOR2_X1 U780 ( .A1(n728), .A2(G953), .ZN(n733) );
  INV_X1 U781 ( .A(G898), .ZN(n731) );
  NAND2_X1 U782 ( .A1(G953), .A2(G224), .ZN(n729) );
  XOR2_X1 U783 ( .A(KEYINPUT61), .B(n729), .Z(n730) );
  NOR2_X1 U784 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U785 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U786 ( .A(n734), .B(KEYINPUT126), .Z(n735) );
  XNOR2_X1 U787 ( .A(n736), .B(n735), .ZN(G69) );
  XNOR2_X1 U788 ( .A(n737), .B(n738), .ZN(n739) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n744), .B(n741), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n748) );
  XNOR2_X1 U792 ( .A(G227), .B(n744), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U794 ( .A1(G953), .A2(n746), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U796 ( .A(G122), .B(n749), .Z(G24) );
  XOR2_X1 U797 ( .A(G131), .B(n750), .Z(G33) );
  XNOR2_X1 U798 ( .A(G137), .B(KEYINPUT127), .ZN(n752) );
  XNOR2_X1 U799 ( .A(n752), .B(n751), .ZN(G39) );
endmodule

