

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763;

  INV_X2 U376 ( .A(G953), .ZN(n752) );
  AND2_X1 U377 ( .A1(n417), .A2(n416), .ZN(n415) );
  AND2_X1 U378 ( .A1(n722), .A2(n752), .ZN(n406) );
  NOR2_X1 U379 ( .A1(n644), .A2(KEYINPUT44), .ZN(n526) );
  NAND2_X1 U380 ( .A1(n415), .A2(n411), .ZN(n708) );
  NAND2_X1 U381 ( .A1(n414), .A2(n412), .ZN(n411) );
  XNOR2_X1 U382 ( .A(G146), .B(G125), .ZN(n475) );
  XNOR2_X1 U383 ( .A(G128), .B(G140), .ZN(n381) );
  XNOR2_X1 U384 ( .A(G110), .B(G119), .ZN(n382) );
  XNOR2_X1 U385 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n440) );
  XNOR2_X2 U386 ( .A(n489), .B(n488), .ZN(n591) );
  XNOR2_X2 U387 ( .A(n461), .B(n497), .ZN(n750) );
  XNOR2_X2 U388 ( .A(n512), .B(n472), .ZN(n461) );
  BUF_X2 U389 ( .A(n534), .Z(n354) );
  XNOR2_X1 U390 ( .A(n444), .B(n362), .ZN(n513) );
  XNOR2_X1 U391 ( .A(n363), .B(KEYINPUT8), .ZN(n362) );
  INV_X1 U392 ( .A(KEYINPUT80), .ZN(n363) );
  NAND2_X1 U393 ( .A1(n626), .A2(n625), .ZN(n751) );
  XNOR2_X1 U394 ( .A(n395), .B(n394), .ZN(n626) );
  INV_X1 U395 ( .A(KEYINPUT48), .ZN(n394) );
  XNOR2_X1 U396 ( .A(n368), .B(n367), .ZN(n480) );
  XNOR2_X1 U397 ( .A(G107), .B(G104), .ZN(n367) );
  XNOR2_X1 U398 ( .A(n426), .B(G110), .ZN(n368) );
  XNOR2_X1 U399 ( .A(G101), .B(KEYINPUT88), .ZN(n426) );
  INV_X1 U400 ( .A(KEYINPUT96), .ZN(n379) );
  INV_X1 U401 ( .A(KEYINPUT46), .ZN(n397) );
  XNOR2_X1 U402 ( .A(G902), .B(KEYINPUT87), .ZN(n435) );
  INV_X1 U403 ( .A(n738), .ZN(n387) );
  XOR2_X1 U404 ( .A(G140), .B(G131), .Z(n497) );
  NOR2_X1 U405 ( .A1(n731), .A2(G902), .ZN(n399) );
  XNOR2_X1 U406 ( .A(n371), .B(n370), .ZN(n479) );
  XNOR2_X1 U407 ( .A(G119), .B(G116), .ZN(n370) );
  XNOR2_X1 U408 ( .A(n451), .B(G113), .ZN(n371) );
  INV_X1 U409 ( .A(KEYINPUT3), .ZN(n451) );
  XNOR2_X1 U410 ( .A(n364), .B(n749), .ZN(n630) );
  XNOR2_X1 U411 ( .A(G107), .B(G116), .ZN(n517) );
  INV_X1 U412 ( .A(KEYINPUT9), .ZN(n516) );
  XNOR2_X1 U413 ( .A(n429), .B(n428), .ZN(n430) );
  INV_X1 U414 ( .A(G146), .ZN(n428) );
  XNOR2_X1 U415 ( .A(n735), .B(n481), .ZN(n664) );
  NAND2_X1 U416 ( .A1(n405), .A2(n404), .ZN(n403) );
  INV_X1 U417 ( .A(KEYINPUT78), .ZN(n402) );
  NAND2_X1 U418 ( .A1(n725), .A2(G217), .ZN(n422) );
  NOR2_X1 U419 ( .A1(n376), .A2(n705), .ZN(n375) );
  AND2_X1 U420 ( .A1(n642), .A2(n379), .ZN(n373) );
  OR2_X1 U421 ( .A1(n638), .A2(n635), .ZN(n544) );
  AND2_X1 U422 ( .A1(n424), .A2(n359), .ZN(n398) );
  XNOR2_X1 U423 ( .A(n607), .B(n397), .ZN(n396) );
  XNOR2_X1 U424 ( .A(n382), .B(n381), .ZN(n442) );
  XNOR2_X1 U425 ( .A(G122), .B(G143), .ZN(n503) );
  XNOR2_X1 U426 ( .A(KEYINPUT75), .B(KEYINPUT89), .ZN(n470) );
  XNOR2_X1 U427 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n474) );
  NAND2_X1 U428 ( .A1(G237), .A2(G234), .ZN(n490) );
  INV_X1 U429 ( .A(KEYINPUT45), .ZN(n568) );
  NAND2_X1 U430 ( .A1(n556), .A2(n393), .ZN(n703) );
  AND2_X1 U431 ( .A1(n466), .A2(n413), .ZN(n412) );
  INV_X1 U432 ( .A(G902), .ZN(n484) );
  XNOR2_X1 U433 ( .A(G146), .B(G131), .ZN(n453) );
  XOR2_X1 U434 ( .A(KEYINPUT94), .B(KEYINPUT72), .Z(n454) );
  XNOR2_X1 U435 ( .A(G137), .B(G101), .ZN(n456) );
  NAND2_X1 U436 ( .A1(n482), .A2(KEYINPUT2), .ZN(n383) );
  NAND2_X1 U437 ( .A1(n387), .A2(n385), .ZN(n384) );
  NOR2_X1 U438 ( .A1(n425), .A2(n629), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n392), .B(n391), .ZN(n717) );
  INV_X1 U440 ( .A(KEYINPUT41), .ZN(n391) );
  NOR2_X1 U441 ( .A1(n704), .A2(n703), .ZN(n392) );
  AND2_X1 U442 ( .A1(n578), .A2(n365), .ZN(n596) );
  NOR2_X1 U443 ( .A1(n605), .A2(n366), .ZN(n365) );
  XNOR2_X1 U444 ( .A(n447), .B(KEYINPUT25), .ZN(n448) );
  XNOR2_X1 U445 ( .A(n369), .B(n480), .ZN(n735) );
  XNOR2_X1 U446 ( .A(n479), .B(n356), .ZN(n369) );
  XNOR2_X1 U447 ( .A(n519), .B(n400), .ZN(n731) );
  XNOR2_X1 U448 ( .A(n512), .B(n518), .ZN(n400) );
  XNOR2_X1 U449 ( .A(n480), .B(n390), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n430), .B(n427), .ZN(n390) );
  NAND2_X1 U451 ( .A1(n687), .A2(n355), .ZN(n409) );
  INV_X1 U452 ( .A(KEYINPUT118), .ZN(n418) );
  XNOR2_X1 U453 ( .A(n422), .B(n421), .ZN(n420) );
  XNOR2_X1 U454 ( .A(n410), .B(G128), .ZN(n679) );
  INV_X1 U455 ( .A(KEYINPUT29), .ZN(n410) );
  XOR2_X1 U456 ( .A(n403), .B(n402), .Z(n355) );
  XOR2_X1 U457 ( .A(KEYINPUT16), .B(G122), .Z(n356) );
  OR2_X1 U458 ( .A1(n573), .A2(n494), .ZN(n357) );
  AND2_X2 U459 ( .A1(n687), .A2(n645), .ZN(n725) );
  XNOR2_X1 U460 ( .A(n399), .B(n520), .ZN(n556) );
  AND2_X1 U461 ( .A1(G221), .A2(n513), .ZN(n358) );
  AND2_X1 U462 ( .A1(n595), .A2(n684), .ZN(n359) );
  AND2_X1 U463 ( .A1(n354), .A2(n691), .ZN(n577) );
  AND2_X1 U464 ( .A1(n627), .A2(KEYINPUT2), .ZN(n360) );
  XNOR2_X1 U465 ( .A(n750), .B(n389), .ZN(n726) );
  XNOR2_X1 U466 ( .A(n435), .B(n434), .ZN(n629) );
  AND2_X1 U467 ( .A1(n631), .A2(G953), .ZN(n734) );
  NAND2_X1 U468 ( .A1(n628), .A2(n627), .ZN(n405) );
  NAND2_X1 U469 ( .A1(n384), .A2(n383), .ZN(n645) );
  XNOR2_X1 U470 ( .A(n591), .B(n401), .ZN(n608) );
  XNOR2_X2 U471 ( .A(n531), .B(n530), .ZN(n560) );
  XNOR2_X1 U472 ( .A(n550), .B(n433), .ZN(n532) );
  BUF_X1 U473 ( .A(n644), .Z(n361) );
  XNOR2_X1 U474 ( .A(n445), .B(n358), .ZN(n364) );
  NAND2_X1 U475 ( .A1(n420), .A2(n667), .ZN(n419) );
  NAND2_X1 U476 ( .A1(n398), .A2(n396), .ZN(n395) );
  INV_X1 U477 ( .A(n577), .ZN(n366) );
  XNOR2_X2 U478 ( .A(n431), .B(KEYINPUT68), .ZN(n472) );
  XNOR2_X2 U479 ( .A(n469), .B(G134), .ZN(n512) );
  XNOR2_X2 U480 ( .A(n372), .B(KEYINPUT0), .ZN(n554) );
  NAND2_X1 U481 ( .A1(n608), .A2(n357), .ZN(n372) );
  XNOR2_X1 U482 ( .A(n549), .B(n548), .ZN(n642) );
  NOR2_X1 U483 ( .A1(n374), .A2(n373), .ZN(n561) );
  NAND2_X1 U484 ( .A1(n377), .A2(n375), .ZN(n374) );
  AND2_X1 U485 ( .A1(n672), .A2(n379), .ZN(n376) );
  NAND2_X1 U486 ( .A1(n380), .A2(n378), .ZN(n377) );
  NOR2_X1 U487 ( .A1(n672), .A2(n379), .ZN(n378) );
  INV_X1 U488 ( .A(n642), .ZN(n380) );
  XNOR2_X2 U489 ( .A(n386), .B(KEYINPUT74), .ZN(n687) );
  NAND2_X1 U490 ( .A1(n628), .A2(n360), .ZN(n386) );
  XNOR2_X2 U491 ( .A(n569), .B(n568), .ZN(n628) );
  XNOR2_X2 U492 ( .A(n388), .B(KEYINPUT71), .ZN(n547) );
  NAND2_X1 U493 ( .A1(n532), .A2(n577), .ZN(n388) );
  XNOR2_X2 U494 ( .A(n432), .B(G469), .ZN(n550) );
  NAND2_X1 U495 ( .A1(n609), .A2(n717), .ZN(n606) );
  INV_X1 U496 ( .A(n557), .ZN(n393) );
  NAND2_X1 U497 ( .A1(n701), .A2(n700), .ZN(n704) );
  INV_X1 U498 ( .A(KEYINPUT19), .ZN(n401) );
  INV_X1 U499 ( .A(KEYINPUT2), .ZN(n404) );
  NAND2_X1 U500 ( .A1(n407), .A2(n406), .ZN(n723) );
  XNOR2_X1 U501 ( .A(n409), .B(n408), .ZN(n407) );
  INV_X1 U502 ( .A(KEYINPUT81), .ZN(n408) );
  INV_X1 U503 ( .A(n468), .ZN(n413) );
  INV_X1 U504 ( .A(n450), .ZN(n414) );
  NAND2_X1 U505 ( .A1(n588), .A2(n468), .ZN(n416) );
  NAND2_X1 U506 ( .A1(n450), .A2(n468), .ZN(n417) );
  NOR2_X2 U507 ( .A1(n708), .A2(n554), .ZN(n495) );
  XNOR2_X1 U508 ( .A(n419), .B(n418), .ZN(G66) );
  INV_X1 U509 ( .A(n630), .ZN(n421) );
  NOR2_X2 U510 ( .A1(n655), .A2(n654), .ZN(n659) );
  NOR2_X2 U511 ( .A1(n655), .A2(n646), .ZN(n650) );
  XNOR2_X1 U512 ( .A(n448), .B(n449), .ZN(n534) );
  BUF_X1 U513 ( .A(n708), .Z(n719) );
  AND2_X1 U514 ( .A1(n615), .A2(KEYINPUT47), .ZN(n423) );
  NOR2_X1 U515 ( .A1(n616), .A2(n423), .ZN(n424) );
  XOR2_X1 U516 ( .A(n751), .B(KEYINPUT73), .Z(n425) );
  INV_X1 U517 ( .A(KEYINPUT5), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U521 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U522 ( .A(G137), .B(KEYINPUT69), .ZN(n439) );
  INV_X1 U523 ( .A(n439), .ZN(n427) );
  NAND2_X1 U524 ( .A1(G227), .A2(n752), .ZN(n429) );
  XNOR2_X2 U525 ( .A(G143), .B(G128), .ZN(n469) );
  XNOR2_X2 U526 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n431) );
  NAND2_X1 U527 ( .A1(n726), .A2(n484), .ZN(n432) );
  XNOR2_X1 U528 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n433) );
  XOR2_X1 U529 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n437) );
  INV_X1 U530 ( .A(KEYINPUT15), .ZN(n434) );
  NAND2_X1 U531 ( .A1(G234), .A2(n629), .ZN(n436) );
  XNOR2_X1 U532 ( .A(n437), .B(n436), .ZN(n446) );
  AND2_X1 U533 ( .A1(n446), .A2(G221), .ZN(n438) );
  XNOR2_X1 U534 ( .A(n438), .B(KEYINPUT21), .ZN(n691) );
  XNOR2_X1 U535 ( .A(KEYINPUT10), .B(n475), .ZN(n496) );
  XNOR2_X1 U536 ( .A(n496), .B(n439), .ZN(n749) );
  XOR2_X1 U537 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n441) );
  XNOR2_X1 U538 ( .A(n441), .B(n440), .ZN(n443) );
  NAND2_X1 U539 ( .A1(G234), .A2(n752), .ZN(n444) );
  NOR2_X1 U540 ( .A1(n630), .A2(G902), .ZN(n449) );
  NAND2_X1 U541 ( .A1(n446), .A2(G217), .ZN(n447) );
  XNOR2_X1 U542 ( .A(n547), .B(KEYINPUT103), .ZN(n450) );
  NOR2_X1 U543 ( .A1(G953), .A2(G237), .ZN(n500) );
  NAND2_X1 U544 ( .A1(n500), .A2(G210), .ZN(n452) );
  XNOR2_X1 U545 ( .A(n479), .B(n452), .ZN(n460) );
  XNOR2_X1 U546 ( .A(n454), .B(n453), .ZN(n458) );
  XNOR2_X1 U547 ( .A(n460), .B(n459), .ZN(n463) );
  BUF_X1 U548 ( .A(n461), .Z(n462) );
  XNOR2_X1 U549 ( .A(n463), .B(n462), .ZN(n657) );
  NAND2_X1 U550 ( .A1(n657), .A2(n484), .ZN(n464) );
  XNOR2_X2 U551 ( .A(n464), .B(G472), .ZN(n574) );
  XNOR2_X1 U552 ( .A(KEYINPUT102), .B(KEYINPUT6), .ZN(n465) );
  XNOR2_X1 U553 ( .A(n574), .B(n465), .ZN(n588) );
  INV_X1 U554 ( .A(n588), .ZN(n466) );
  XOR2_X1 U555 ( .A(KEYINPUT33), .B(KEYINPUT104), .Z(n467) );
  XNOR2_X1 U556 ( .A(n467), .B(KEYINPUT86), .ZN(n468) );
  XNOR2_X1 U557 ( .A(n469), .B(n470), .ZN(n471) );
  XNOR2_X1 U558 ( .A(n472), .B(n471), .ZN(n478) );
  NAND2_X1 U559 ( .A1(n752), .A2(G224), .ZN(n473) );
  XNOR2_X1 U560 ( .A(n474), .B(n473), .ZN(n476) );
  XNOR2_X1 U561 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U562 ( .A(n478), .B(n477), .ZN(n481) );
  INV_X1 U563 ( .A(n629), .ZN(n482) );
  NOR2_X1 U564 ( .A1(n664), .A2(n482), .ZN(n486) );
  INV_X1 U565 ( .A(G237), .ZN(n483) );
  NAND2_X1 U566 ( .A1(n484), .A2(n483), .ZN(n487) );
  NAND2_X1 U567 ( .A1(n487), .A2(G210), .ZN(n485) );
  XNOR2_X1 U568 ( .A(n486), .B(n485), .ZN(n579) );
  NAND2_X1 U569 ( .A1(n487), .A2(G214), .ZN(n700) );
  NAND2_X1 U570 ( .A1(n579), .A2(n700), .ZN(n489) );
  INV_X1 U571 ( .A(KEYINPUT84), .ZN(n488) );
  XNOR2_X1 U572 ( .A(n490), .B(KEYINPUT14), .ZN(n491) );
  XNOR2_X1 U573 ( .A(KEYINPUT70), .B(n491), .ZN(n492) );
  NAND2_X1 U574 ( .A1(G952), .A2(n492), .ZN(n716) );
  NOR2_X1 U575 ( .A1(n716), .A2(G953), .ZN(n573) );
  NAND2_X1 U576 ( .A1(n492), .A2(G902), .ZN(n570) );
  NOR2_X1 U577 ( .A1(G898), .A2(n752), .ZN(n493) );
  XOR2_X1 U578 ( .A(KEYINPUT90), .B(n493), .Z(n736) );
  NOR2_X1 U579 ( .A1(n570), .A2(n736), .ZN(n494) );
  XNOR2_X1 U580 ( .A(n495), .B(KEYINPUT34), .ZN(n522) );
  XNOR2_X1 U581 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n510) );
  XNOR2_X1 U582 ( .A(n496), .B(G104), .ZN(n499) );
  XOR2_X1 U583 ( .A(n497), .B(G113), .Z(n498) );
  XNOR2_X1 U584 ( .A(n499), .B(n498), .ZN(n508) );
  XOR2_X1 U585 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n502) );
  NAND2_X1 U586 ( .A1(n500), .A2(G214), .ZN(n501) );
  XNOR2_X1 U587 ( .A(n502), .B(n501), .ZN(n506) );
  XOR2_X1 U588 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n504) );
  XNOR2_X1 U589 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U590 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U591 ( .A(n508), .B(n507), .ZN(n648) );
  NOR2_X1 U592 ( .A1(G902), .A2(n648), .ZN(n509) );
  XNOR2_X1 U593 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U594 ( .A(G475), .ZN(n646) );
  XNOR2_X1 U595 ( .A(n511), .B(n646), .ZN(n557) );
  XOR2_X1 U596 ( .A(G122), .B(KEYINPUT7), .Z(n515) );
  NAND2_X1 U597 ( .A1(G217), .A2(n513), .ZN(n514) );
  XNOR2_X1 U598 ( .A(n515), .B(n514), .ZN(n519) );
  XNOR2_X1 U599 ( .A(KEYINPUT100), .B(G478), .ZN(n520) );
  INV_X1 U600 ( .A(n556), .ZN(n527) );
  NAND2_X1 U601 ( .A1(n557), .A2(n527), .ZN(n580) );
  INV_X1 U602 ( .A(n580), .ZN(n521) );
  NAND2_X1 U603 ( .A1(n522), .A2(n521), .ZN(n524) );
  XNOR2_X1 U604 ( .A(KEYINPUT76), .B(KEYINPUT35), .ZN(n523) );
  XNOR2_X2 U605 ( .A(n524), .B(n523), .ZN(n644) );
  INV_X1 U606 ( .A(KEYINPUT67), .ZN(n525) );
  XNOR2_X1 U607 ( .A(n526), .B(n525), .ZN(n543) );
  INV_X1 U608 ( .A(n703), .ZN(n528) );
  NAND2_X1 U609 ( .A1(n528), .A2(n691), .ZN(n529) );
  OR2_X1 U610 ( .A1(n554), .A2(n529), .ZN(n531) );
  XNOR2_X1 U611 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n530) );
  BUF_X1 U612 ( .A(n532), .Z(n533) );
  INV_X1 U613 ( .A(n533), .ZN(n688) );
  INV_X1 U614 ( .A(n354), .ZN(n587) );
  AND2_X1 U615 ( .A1(n588), .A2(n587), .ZN(n535) );
  NAND2_X1 U616 ( .A1(n533), .A2(n535), .ZN(n536) );
  XNOR2_X1 U617 ( .A(n536), .B(KEYINPUT77), .ZN(n537) );
  NAND2_X1 U618 ( .A1(n560), .A2(n537), .ZN(n539) );
  INV_X1 U619 ( .A(KEYINPUT32), .ZN(n538) );
  XNOR2_X1 U620 ( .A(n539), .B(n538), .ZN(n638) );
  OR2_X1 U621 ( .A1(n574), .A2(n354), .ZN(n540) );
  NOR2_X1 U622 ( .A1(n533), .A2(n540), .ZN(n541) );
  AND2_X1 U623 ( .A1(n560), .A2(n541), .ZN(n635) );
  INV_X1 U624 ( .A(n544), .ZN(n542) );
  NAND2_X1 U625 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U626 ( .A1(n544), .A2(KEYINPUT44), .ZN(n545) );
  NAND2_X1 U627 ( .A1(n546), .A2(n545), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n644), .A2(KEYINPUT44), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n547), .A2(n574), .ZN(n696) );
  NOR2_X1 U630 ( .A1(n696), .A2(n554), .ZN(n549) );
  XNOR2_X1 U631 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n548) );
  BUF_X1 U632 ( .A(n550), .Z(n551) );
  NOR2_X1 U633 ( .A1(n574), .A2(n366), .ZN(n552) );
  NAND2_X1 U634 ( .A1(n551), .A2(n552), .ZN(n553) );
  NOR2_X1 U635 ( .A1(n554), .A2(n553), .ZN(n672) );
  OR2_X1 U636 ( .A1(n557), .A2(n556), .ZN(n641) );
  INV_X1 U637 ( .A(KEYINPUT101), .ZN(n555) );
  XNOR2_X1 U638 ( .A(n641), .B(n555), .ZN(n623) );
  NAND2_X1 U639 ( .A1(n557), .A2(n556), .ZN(n633) );
  AND2_X1 U640 ( .A1(n623), .A2(n633), .ZN(n705) );
  NAND2_X1 U641 ( .A1(n588), .A2(n354), .ZN(n558) );
  NOR2_X1 U642 ( .A1(n533), .A2(n558), .ZN(n559) );
  AND2_X1 U643 ( .A1(n560), .A2(n559), .ZN(n636) );
  NOR2_X1 U644 ( .A1(n561), .A2(n636), .ZN(n562) );
  NAND2_X1 U645 ( .A1(n563), .A2(n562), .ZN(n565) );
  INV_X1 U646 ( .A(KEYINPUT83), .ZN(n564) );
  XNOR2_X1 U647 ( .A(n565), .B(n564), .ZN(n566) );
  NOR2_X2 U648 ( .A1(n567), .A2(n566), .ZN(n569) );
  INV_X1 U649 ( .A(n551), .ZN(n605) );
  OR2_X1 U650 ( .A1(n752), .A2(n570), .ZN(n571) );
  NOR2_X1 U651 ( .A1(G900), .A2(n571), .ZN(n572) );
  NOR2_X1 U652 ( .A1(n573), .A2(n572), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n574), .A2(n700), .ZN(n575) );
  XNOR2_X1 U654 ( .A(KEYINPUT30), .B(n575), .ZN(n576) );
  NOR2_X1 U655 ( .A1(n585), .A2(n576), .ZN(n578) );
  INV_X1 U656 ( .A(n579), .ZN(n621) );
  NOR2_X1 U657 ( .A1(n580), .A2(n621), .ZN(n581) );
  NAND2_X1 U658 ( .A1(n596), .A2(n581), .ZN(n632) );
  INV_X1 U659 ( .A(n632), .ZN(n583) );
  INV_X1 U660 ( .A(KEYINPUT79), .ZN(n613) );
  NOR2_X1 U661 ( .A1(KEYINPUT47), .A2(n613), .ZN(n582) );
  NOR2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n595) );
  INV_X1 U663 ( .A(n691), .ZN(n584) );
  NOR2_X1 U664 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n601) );
  INV_X1 U666 ( .A(n601), .ZN(n590) );
  NOR2_X1 U667 ( .A1(n588), .A2(n633), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n617) );
  INV_X1 U669 ( .A(n591), .ZN(n592) );
  NOR2_X1 U670 ( .A1(n617), .A2(n592), .ZN(n593) );
  XNOR2_X1 U671 ( .A(n593), .B(KEYINPUT36), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n594), .A2(n533), .ZN(n684) );
  XNOR2_X1 U673 ( .A(n621), .B(KEYINPUT38), .ZN(n701) );
  AND2_X1 U674 ( .A1(n596), .A2(n701), .ZN(n597) );
  XNOR2_X1 U675 ( .A(KEYINPUT39), .B(n597), .ZN(n624) );
  NOR2_X1 U676 ( .A1(n624), .A2(n633), .ZN(n600) );
  XNOR2_X1 U677 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n598) );
  XNOR2_X1 U678 ( .A(n598), .B(KEYINPUT107), .ZN(n599) );
  XNOR2_X1 U679 ( .A(n600), .B(n599), .ZN(n762) );
  INV_X1 U680 ( .A(n574), .ZN(n602) );
  NOR2_X1 U681 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U682 ( .A(KEYINPUT28), .B(n603), .Z(n604) );
  NOR2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n609) );
  XNOR2_X1 U684 ( .A(n606), .B(KEYINPUT42), .ZN(n763) );
  NAND2_X1 U685 ( .A1(n762), .A2(n763), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n612), .A2(KEYINPUT47), .ZN(n610) );
  NOR2_X1 U688 ( .A1(KEYINPUT79), .A2(n610), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n705), .A2(n611), .ZN(n616) );
  INV_X1 U690 ( .A(n612), .ZN(n681) );
  NAND2_X1 U691 ( .A1(n705), .A2(n613), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n681), .A2(n614), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n533), .A2(n617), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n700), .A2(n618), .ZN(n619) );
  XOR2_X1 U695 ( .A(KEYINPUT43), .B(n619), .Z(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT105), .ZN(n622) );
  AND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n639) );
  NOR2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n686) );
  NOR2_X1 U699 ( .A1(n639), .A2(n686), .ZN(n625) );
  INV_X1 U700 ( .A(n751), .ZN(n627) );
  INV_X1 U701 ( .A(n628), .ZN(n738) );
  INV_X1 U702 ( .A(G952), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(G143), .ZN(G45) );
  INV_X1 U704 ( .A(n633), .ZN(n680) );
  NAND2_X1 U705 ( .A1(n672), .A2(n680), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n634), .B(G104), .ZN(G6) );
  XOR2_X1 U707 ( .A(G110), .B(n635), .Z(G12) );
  XOR2_X1 U708 ( .A(G101), .B(n636), .Z(G3) );
  XNOR2_X1 U709 ( .A(G119), .B(KEYINPUT127), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(G21) );
  XOR2_X1 U711 ( .A(n639), .B(G140), .Z(G42) );
  NAND2_X1 U712 ( .A1(n642), .A2(n680), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n640), .B(G113), .ZN(G15) );
  INV_X1 U714 ( .A(n641), .ZN(n677) );
  NAND2_X1 U715 ( .A1(n642), .A2(n677), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(G116), .ZN(G18) );
  XOR2_X1 U717 ( .A(n361), .B(G122), .Z(G24) );
  NAND2_X1 U718 ( .A1(n645), .A2(n687), .ZN(n655) );
  XOR2_X1 U719 ( .A(KEYINPUT116), .B(KEYINPUT59), .Z(n647) );
  XNOR2_X1 U720 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(n651) );
  INV_X1 U722 ( .A(n734), .ZN(n667) );
  NAND2_X1 U723 ( .A1(n651), .A2(n667), .ZN(n653) );
  XNOR2_X1 U724 ( .A(KEYINPUT117), .B(KEYINPUT60), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(G60) );
  INV_X1 U726 ( .A(G472), .ZN(n654) );
  XOR2_X1 U727 ( .A(KEYINPUT108), .B(KEYINPUT62), .Z(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n660), .A2(n667), .ZN(n661) );
  XNOR2_X1 U731 ( .A(n661), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U732 ( .A1(n725), .A2(G210), .ZN(n666) );
  XNOR2_X1 U733 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n662) );
  XOR2_X1 U734 ( .A(n662), .B(KEYINPUT85), .Z(n663) );
  XNOR2_X1 U735 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n666), .B(n665), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n671) );
  XNOR2_X1 U738 ( .A(KEYINPUT115), .B(KEYINPUT56), .ZN(n669) );
  XNOR2_X1 U739 ( .A(n669), .B(KEYINPUT82), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(G51) );
  NAND2_X1 U741 ( .A1(n672), .A2(n677), .ZN(n674) );
  XOR2_X1 U742 ( .A(KEYINPUT109), .B(KEYINPUT27), .Z(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(n676) );
  XOR2_X1 U744 ( .A(G107), .B(KEYINPUT26), .Z(n675) );
  XNOR2_X1 U745 ( .A(n676), .B(n675), .ZN(G9) );
  NAND2_X1 U746 ( .A1(n681), .A2(n677), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(G30) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(G146), .ZN(G48) );
  XOR2_X1 U750 ( .A(KEYINPUT37), .B(KEYINPUT110), .Z(n683) );
  XNOR2_X1 U751 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U752 ( .A(G125), .B(n685), .ZN(G27) );
  XOR2_X1 U753 ( .A(G134), .B(n686), .Z(G36) );
  XOR2_X1 U754 ( .A(KEYINPUT114), .B(KEYINPUT53), .Z(n724) );
  NAND2_X1 U755 ( .A1(n688), .A2(n366), .ZN(n689) );
  XOR2_X1 U756 ( .A(KEYINPUT50), .B(n689), .Z(n690) );
  XNOR2_X1 U757 ( .A(n690), .B(KEYINPUT111), .ZN(n695) );
  NOR2_X1 U758 ( .A1(n354), .A2(n691), .ZN(n692) );
  XOR2_X1 U759 ( .A(KEYINPUT49), .B(n692), .Z(n693) );
  NOR2_X1 U760 ( .A1(n574), .A2(n693), .ZN(n694) );
  NAND2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U763 ( .A(KEYINPUT51), .B(n698), .Z(n699) );
  NAND2_X1 U764 ( .A1(n699), .A2(n717), .ZN(n712) );
  NOR2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n709), .A2(n719), .ZN(n710) );
  XOR2_X1 U770 ( .A(KEYINPUT112), .B(n710), .Z(n711) );
  NAND2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n713), .B(KEYINPUT113), .ZN(n714) );
  XNOR2_X1 U773 ( .A(n714), .B(KEYINPUT52), .ZN(n715) );
  NOR2_X1 U774 ( .A1(n716), .A2(n715), .ZN(n721) );
  INV_X1 U775 ( .A(n717), .ZN(n718) );
  NOR2_X1 U776 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U777 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n724), .B(n723), .ZN(G75) );
  NAND2_X1 U779 ( .A1(n725), .A2(G469), .ZN(n729) );
  XOR2_X1 U780 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n727) );
  XOR2_X1 U781 ( .A(n727), .B(n726), .Z(n728) );
  XNOR2_X1 U782 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n734), .A2(n730), .ZN(G54) );
  NAND2_X1 U784 ( .A1(n725), .A2(G478), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n732), .B(n731), .ZN(n733) );
  NOR2_X1 U786 ( .A1(n734), .A2(n733), .ZN(G63) );
  XOR2_X1 U787 ( .A(KEYINPUT122), .B(n735), .Z(n737) );
  NAND2_X1 U788 ( .A1(n737), .A2(n736), .ZN(n748) );
  NOR2_X1 U789 ( .A1(n738), .A2(G953), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n739), .B(KEYINPUT121), .ZN(n745) );
  XOR2_X1 U791 ( .A(KEYINPUT61), .B(KEYINPUT120), .Z(n741) );
  NAND2_X1 U792 ( .A1(G224), .A2(G953), .ZN(n740) );
  XNOR2_X1 U793 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U794 ( .A(KEYINPUT119), .B(n742), .ZN(n743) );
  NAND2_X1 U795 ( .A1(n743), .A2(G898), .ZN(n744) );
  NAND2_X1 U796 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n746), .B(KEYINPUT123), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n748), .B(n747), .ZN(G69) );
  XOR2_X1 U799 ( .A(n750), .B(n749), .Z(n755) );
  XNOR2_X1 U800 ( .A(n755), .B(n751), .ZN(n753) );
  NAND2_X1 U801 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U802 ( .A(KEYINPUT124), .B(n754), .ZN(n761) );
  XNOR2_X1 U803 ( .A(G227), .B(n755), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(G900), .ZN(n757) );
  XOR2_X1 U805 ( .A(KEYINPUT125), .B(n757), .Z(n758) );
  NAND2_X1 U806 ( .A1(G953), .A2(n758), .ZN(n759) );
  XNOR2_X1 U807 ( .A(KEYINPUT126), .B(n759), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(G72) );
  XNOR2_X1 U809 ( .A(n762), .B(G131), .ZN(G33) );
  XNOR2_X1 U810 ( .A(G137), .B(n763), .ZN(G39) );
endmodule

