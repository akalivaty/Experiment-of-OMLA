//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G137), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n196), .A3(new_n200), .A4(new_n197), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  OR2_X1    g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n203), .B(new_n204), .C1(new_n206), .C2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT64), .B1(new_n205), .B2(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n207), .A3(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n205), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(new_n203), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n191), .B1(new_n202), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n218));
  OAI21_X1  g032(.A(G128), .B1(new_n206), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n206), .B2(new_n208), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n193), .A2(G137), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n195), .A2(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n201), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n216), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n199), .A2(new_n201), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT68), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n217), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT2), .B(G113), .Z(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT67), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n234), .A2(new_n235), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT70), .B(G237), .ZN(new_n240));
  INV_X1    g054(.A(G953), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(G210), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT27), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G101), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n216), .A2(KEYINPUT65), .B1(new_n199), .B2(new_n201), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n209), .A2(new_n215), .A3(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n249), .A2(new_n251), .B1(new_n224), .B2(new_n228), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n248), .B1(new_n252), .B2(KEYINPUT30), .ZN(new_n253));
  AND4_X1   g067(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n254));
  XNOR2_X1  g068(.A(G143), .B(G146), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT0), .B(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT65), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n231), .A3(new_n251), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n229), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(KEYINPUT66), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n217), .A2(KEYINPUT30), .A3(new_n229), .A4(new_n232), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n264), .A2(new_n238), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT69), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT69), .B1(new_n263), .B2(new_n265), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n247), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT66), .B1(new_n260), .B2(new_n261), .ZN(new_n272));
  AOI211_X1 g086(.A(new_n248), .B(KEYINPUT30), .C1(new_n259), .C2(new_n229), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n264), .A2(new_n238), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT31), .A3(new_n247), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n270), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n238), .B1(new_n224), .B2(new_n228), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n230), .A2(new_n231), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT28), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n260), .A2(new_n238), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n239), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g099(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(new_n245), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT72), .B1(new_n280), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n291), .B(new_n288), .C1(new_n270), .C2(new_n279), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n190), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n294));
  INV_X1    g108(.A(new_n239), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n276), .B2(new_n277), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n296), .B2(new_n245), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n239), .B1(new_n266), .B2(new_n267), .ZN(new_n298));
  INV_X1    g112(.A(new_n245), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(KEYINPUT73), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n287), .B2(new_n245), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n233), .B(new_n238), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n283), .B1(new_n303), .B2(KEYINPUT28), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n245), .A2(KEYINPUT29), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G472), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT31), .B1(new_n278), .B2(new_n247), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n269), .B(new_n246), .C1(new_n276), .C2(new_n277), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n289), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n291), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n280), .A2(KEYINPUT72), .A3(new_n289), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n188), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n293), .B(new_n308), .C1(new_n314), .C2(KEYINPUT32), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(G234), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT77), .ZN(new_n324));
  XNOR2_X1  g138(.A(G125), .B(G140), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n327), .A3(new_n207), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G146), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT24), .B(G110), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n221), .A2(G119), .ZN(new_n336));
  INV_X1    g150(.A(G119), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G128), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n335), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(G128), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n221), .A2(G119), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT74), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n334), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n346), .B(new_n340), .C1(new_n338), .C2(KEYINPUT23), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(G110), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n348), .B1(new_n343), .B2(new_n344), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n332), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G110), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n347), .B2(KEYINPUT75), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(KEYINPUT75), .B2(new_n347), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n339), .A2(new_n334), .A3(new_n342), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n329), .A2(new_n330), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n207), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n331), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(KEYINPUT78), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n361));
  INV_X1    g175(.A(new_n359), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(new_n350), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT22), .B(G137), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n241), .A2(G221), .A3(G234), .ZN(new_n365));
  XOR2_X1   g179(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n351), .A2(new_n359), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n361), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT25), .B1(new_n371), .B2(new_n317), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n373));
  AOI211_X1 g187(.A(new_n373), .B(G902), .C1(new_n368), .C2(new_n370), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n318), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n318), .A2(G902), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n219), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n223), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(new_n382), .B2(G107), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G104), .ZN(new_n386));
  INV_X1    g200(.A(G101), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(G107), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n383), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT80), .B1(new_n382), .B2(G107), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n388), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n382), .A2(KEYINPUT80), .A3(G107), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n381), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n395), .A2(KEYINPUT10), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n383), .A2(new_n386), .A3(new_n388), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(G101), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(G101), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n230), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n393), .A2(new_n405), .A3(new_n389), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n393), .B2(new_n389), .ZN(new_n408));
  OAI211_X1 g222(.A(KEYINPUT10), .B(new_n224), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n396), .A2(new_n202), .A3(new_n404), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n393), .A2(new_n389), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT81), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n412), .A2(new_n223), .A3(new_n220), .A4(new_n406), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n202), .B1(new_n413), .B2(new_n394), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT82), .A3(KEYINPUT12), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n407), .A2(new_n408), .A3(new_n224), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n231), .B1(new_n416), .B2(new_n395), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT12), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n418), .B(new_n202), .C1(new_n413), .C2(new_n394), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(KEYINPUT82), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n410), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n241), .A2(G227), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n410), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n396), .A2(new_n404), .A3(new_n409), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n231), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n423), .A2(new_n426), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G469), .ZN(new_n433));
  INV_X1    g247(.A(G469), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n415), .A2(new_n419), .ZN(new_n435));
  INV_X1    g249(.A(new_n422), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n428), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n427), .B1(new_n431), .B2(new_n410), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n434), .B(new_n317), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n434), .A2(new_n317), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n433), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G221), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT9), .B(G234), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n445), .B2(new_n317), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(KEYINPUT70), .A2(G237), .ZN(new_n449));
  NOR2_X1   g263(.A1(KEYINPUT70), .A2(G237), .ZN(new_n450));
  OAI211_X1 g264(.A(G214), .B(new_n241), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n205), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n240), .A2(G143), .A3(G214), .A4(new_n241), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT18), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(new_n200), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT84), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(KEYINPUT84), .A3(new_n456), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n328), .B1(new_n207), .B2(new_n325), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n452), .B(new_n453), .C1(new_n455), .C2(new_n200), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n382), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n452), .A2(new_n453), .A3(new_n200), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n200), .B1(new_n452), .B2(new_n453), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT86), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n358), .B1(KEYINPUT17), .B2(new_n470), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n454), .A2(G131), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n452), .A2(new_n453), .A3(new_n200), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(KEYINPUT86), .A3(new_n472), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n466), .B(new_n468), .C1(new_n473), .C2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n468), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n464), .B1(new_n459), .B2(new_n460), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT19), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n324), .A2(new_n327), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n323), .A2(KEYINPUT85), .A3(KEYINPUT19), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n325), .B2(new_n482), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n483), .A2(new_n207), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n487), .B(new_n331), .C1(new_n470), .C2(new_n469), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n480), .B1(new_n481), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n479), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G475), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n317), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT20), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n479), .A2(new_n490), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n492), .A4(new_n317), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n466), .B1(new_n478), .B2(new_n473), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n480), .ZN(new_n500));
  AOI21_X1  g314(.A(G902), .B1(new_n500), .B2(new_n479), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G475), .B1(new_n501), .B2(new_n502), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n498), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(G234), .A2(G237), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n508), .A2(G952), .A3(new_n241), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(G902), .A3(G953), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n510), .B(KEYINPUT92), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT21), .B(G898), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G116), .B(G122), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n385), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n205), .A2(G128), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n221), .A2(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G134), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n519), .A3(new_n193), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n526));
  INV_X1    g340(.A(G122), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(G116), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n385), .B1(new_n528), .B2(KEYINPUT14), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n525), .B2(new_n529), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n517), .B(new_n523), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G116), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G122), .ZN(new_n534));
  OAI21_X1  g348(.A(G107), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT89), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n517), .A2(new_n535), .B1(new_n536), .B2(new_n522), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n522), .A2(new_n536), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n221), .B2(G143), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n205), .A2(KEYINPUT13), .A3(G128), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n519), .A3(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n542), .A2(KEYINPUT88), .A3(G134), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT88), .B1(new_n542), .B2(G134), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n537), .B(new_n538), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n532), .A2(new_n545), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n444), .A2(new_n316), .A3(G953), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n532), .A2(new_n545), .A3(new_n547), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n546), .A2(KEYINPUT91), .A3(new_n548), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n317), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G478), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n554), .B(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n507), .A2(new_n515), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G214), .B1(G237), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G224), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G953), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT7), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n224), .A2(G125), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n230), .A2(new_n321), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n563), .A2(KEYINPUT83), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI221_X1 g385(.A(new_n565), .B1(KEYINPUT83), .B2(new_n563), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G122), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT8), .Z(new_n575));
  NAND2_X1  g389(.A1(new_n234), .A2(new_n235), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n337), .A2(G116), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n577), .B(G113), .C1(KEYINPUT5), .C2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n576), .B(new_n579), .C1(new_n407), .C2(new_n408), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n576), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n411), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n575), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n573), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n401), .A2(new_n238), .A3(new_n403), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n580), .A3(new_n574), .ZN(new_n586));
  AOI21_X1  g400(.A(G902), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n580), .ZN(new_n588));
  INV_X1    g402(.A(new_n574), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(KEYINPUT6), .A3(new_n586), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT6), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(new_n592), .A3(new_n589), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n569), .B(new_n564), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G210), .B1(G237), .B2(G902), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n587), .A2(new_n597), .A3(new_n595), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n561), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n448), .A2(new_n559), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n315), .A2(new_n378), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  OAI21_X1  g419(.A(new_n317), .B1(new_n290), .B2(new_n292), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G472), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n187), .B1(new_n290), .B2(new_n292), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n378), .A2(new_n442), .A3(new_n447), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n549), .A2(KEYINPUT33), .A3(new_n551), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n552), .A2(new_n612), .A3(new_n553), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT93), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n552), .A2(new_n615), .A3(new_n612), .A4(new_n553), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n611), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n555), .A2(G902), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n554), .A2(new_n555), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n506), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n601), .A2(new_n515), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n610), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT34), .B(G104), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  INV_X1    g440(.A(new_n505), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n503), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n498), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n494), .A2(KEYINPUT94), .A3(new_n497), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n628), .A2(new_n630), .A3(new_n557), .A4(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n610), .A2(new_n623), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT95), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  INV_X1    g450(.A(new_n376), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n367), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n369), .B(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n375), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n442), .A2(new_n641), .A3(new_n601), .A4(new_n447), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n559), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n607), .A3(new_n608), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  NAND2_X1  g460(.A1(new_n312), .A2(new_n313), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n647), .A2(new_n190), .B1(G472), .B2(new_n307), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n608), .A2(new_n189), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n642), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n509), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT96), .B(G900), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n651), .B1(new_n511), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n630), .A2(new_n631), .A3(new_n653), .ZN(new_n654));
  AOI211_X1 g468(.A(new_n558), .B(new_n654), .C1(new_n503), .C2(new_n627), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  INV_X1    g471(.A(G472), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n303), .A2(new_n299), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n268), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n660), .A2(KEYINPUT97), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n660), .B2(KEYINPUT97), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n647), .B2(new_n190), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n649), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n653), .B(KEYINPUT39), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n442), .A2(new_n447), .A3(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n599), .A2(new_n600), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT38), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n599), .A2(KEYINPUT38), .A3(new_n600), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n557), .A2(new_n560), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n674), .A2(new_n641), .A3(new_n507), .A4(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n665), .A2(new_n668), .A3(new_n669), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  NAND3_X1  g492(.A1(new_n506), .A2(new_n621), .A3(new_n653), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT98), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n506), .A2(new_n621), .A3(KEYINPUT98), .A4(new_n653), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n650), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NAND2_X1  g500(.A1(new_n435), .A2(new_n436), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n438), .B1(new_n687), .B2(new_n429), .ZN(new_n688));
  OAI21_X1  g502(.A(G469), .B1(new_n688), .B2(G902), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n447), .A3(new_n439), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n623), .A2(new_n690), .A3(new_n622), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n315), .A2(new_n378), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NOR3_X1   g508(.A1(new_n623), .A2(new_n632), .A3(new_n690), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n315), .A2(new_n378), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  INV_X1    g511(.A(new_n690), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n601), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n507), .A2(new_n641), .A3(new_n515), .A4(new_n558), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n315), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NOR4_X1   g517(.A1(new_n623), .A2(new_n690), .A3(new_n507), .A4(new_n558), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT99), .B(G472), .Z(new_n706));
  OAI21_X1  g520(.A(new_n280), .B1(new_n245), .B2(new_n304), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n606), .A2(new_n706), .B1(new_n187), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(KEYINPUT100), .A3(new_n378), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n187), .ZN(new_n710));
  AOI21_X1  g524(.A(G902), .B1(new_n312), .B2(new_n313), .ZN(new_n711));
  INV_X1    g525(.A(new_n706), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n378), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n705), .B1(new_n709), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n527), .ZN(G24));
  INV_X1    g531(.A(new_n699), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n708), .A2(new_n684), .A3(new_n718), .A4(new_n641), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NOR2_X1   g534(.A1(new_n446), .A2(new_n561), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n599), .A2(new_n600), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n423), .A2(new_n426), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n429), .A2(new_n431), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(KEYINPUT101), .A3(G469), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n439), .A3(new_n441), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT101), .B1(new_n432), .B2(G469), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n722), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n722), .B(KEYINPUT102), .C1(new_n726), .C2(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n315), .A3(new_n378), .A4(new_n684), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n314), .B2(KEYINPUT32), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n608), .A2(KEYINPUT104), .A3(new_n189), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n648), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n683), .B1(new_n730), .B2(new_n731), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n740), .A4(new_n378), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT105), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n732), .A2(KEYINPUT42), .A3(new_n684), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n378), .A4(new_n739), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n735), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n200), .ZN(G33));
  NAND4_X1  g561(.A1(new_n732), .A2(new_n315), .A3(new_n378), .A4(new_n655), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  OAI21_X1  g563(.A(G469), .B1(new_n432), .B2(KEYINPUT45), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n750), .A2(KEYINPUT106), .B1(KEYINPUT45), .B2(new_n432), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n752), .B(G469), .C1(new_n432), .C2(KEYINPUT45), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n440), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n439), .B1(new_n754), .B2(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n750), .A2(KEYINPUT106), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n432), .A2(KEYINPUT45), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n441), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n447), .B(new_n666), .C1(new_n755), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n607), .A2(new_n608), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n617), .A2(new_n618), .B1(new_n555), .B2(new_n554), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n506), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT43), .B1(new_n506), .B2(new_n764), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n767), .A2(new_n641), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT44), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n762), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n763), .A2(new_n769), .A3(KEYINPUT44), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n587), .A2(new_n597), .A3(new_n595), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n597), .B1(new_n587), .B2(new_n595), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n774), .A3(new_n561), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n772), .A2(KEYINPUT107), .A3(new_n775), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n771), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT108), .B(G137), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  NAND2_X1  g596(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n447), .B(new_n783), .C1(new_n755), .C2(new_n761), .ZN(new_n784));
  INV_X1    g598(.A(new_n775), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n315), .A2(new_n378), .A3(new_n683), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n439), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n759), .B2(new_n760), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n754), .A2(KEYINPUT46), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n446), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n791));
  OAI211_X1 g605(.A(new_n784), .B(new_n786), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NOR2_X1   g607(.A1(new_n507), .A2(new_n558), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n726), .A2(new_n727), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n653), .A2(new_n447), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n795), .A2(new_n641), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n665), .A2(new_n601), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n642), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n315), .B(new_n799), .C1(new_n684), .C2(new_n655), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n800), .A3(new_n719), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n798), .A2(new_n800), .A3(KEYINPUT52), .A4(new_n719), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n801), .A2(KEYINPUT113), .A3(new_n802), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n742), .A2(new_n745), .ZN(new_n810));
  INV_X1    g624(.A(new_n735), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n732), .A2(new_n708), .A3(new_n641), .A4(new_n684), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n641), .A2(new_n775), .A3(new_n628), .A4(new_n558), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n814), .A2(new_n448), .A3(new_n654), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n315), .A2(KEYINPUT112), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT112), .B1(new_n315), .B2(new_n815), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n748), .B(new_n813), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n692), .A2(new_n696), .A3(new_n702), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n507), .A2(new_n557), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n623), .B1(new_n820), .B2(new_n622), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n607), .A2(new_n821), .A3(new_n608), .A4(new_n609), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n604), .A2(new_n644), .A3(new_n822), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n818), .A2(new_n716), .A3(new_n819), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n808), .A2(new_n809), .A3(new_n812), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n803), .A2(new_n805), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n812), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n809), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n748), .A2(new_n813), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n604), .A2(new_n644), .A3(new_n822), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n315), .A2(new_n815), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n315), .A2(KEYINPUT112), .A3(new_n815), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n831), .A2(new_n832), .A3(new_n837), .A4(KEYINPUT53), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n746), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n709), .A2(new_n715), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n704), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n692), .A2(new_n696), .A3(new_n702), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT114), .B1(new_n716), .B2(new_n819), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n839), .A2(new_n807), .A3(new_n806), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n830), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n829), .B1(KEYINPUT54), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n690), .A2(new_n785), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n378), .A2(new_n509), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n665), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n507), .A3(new_n764), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n767), .A2(new_n768), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n509), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n851), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n641), .A3(new_n708), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n856), .B1(new_n709), .B2(new_n715), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(new_n561), .A3(new_n674), .A4(new_n698), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n859), .B1(new_n861), .B2(KEYINPUT50), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(KEYINPUT50), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n784), .B1(new_n790), .B2(new_n791), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n689), .A2(new_n439), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n447), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n775), .A3(new_n860), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT51), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n857), .A2(new_n378), .A3(new_n739), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT48), .ZN(new_n875));
  INV_X1    g689(.A(G952), .ZN(new_n876));
  INV_X1    g690(.A(new_n622), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n876), .B(G953), .C1(new_n853), .C2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n860), .A2(KEYINPUT117), .A3(new_n718), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT117), .B1(new_n860), .B2(new_n718), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n875), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n862), .A2(new_n872), .A3(new_n863), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT116), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n873), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n849), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n867), .A2(KEYINPUT49), .B1(new_n673), .B2(new_n672), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(KEYINPUT49), .B2(new_n867), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n378), .A2(KEYINPUT110), .A3(new_n721), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n765), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT110), .B1(new_n378), .B2(new_n721), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n889), .B1(new_n893), .B2(KEYINPUT111), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(KEYINPUT111), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n887), .B1(new_n665), .B2(new_n895), .ZN(G75));
  NAND2_X1  g710(.A1(new_n876), .A2(G953), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT118), .Z(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n848), .A2(G902), .ZN(new_n901));
  INV_X1    g715(.A(G210), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n591), .A2(new_n593), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(new_n594), .Z(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT55), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n906), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n900), .B(new_n908), .C1(new_n901), .C2(new_n902), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n907), .B2(new_n909), .ZN(G51));
  XNOR2_X1  g724(.A(new_n440), .B(KEYINPUT57), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n830), .A2(new_n912), .A3(new_n847), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n830), .B2(new_n847), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n688), .B(KEYINPUT119), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n901), .A2(new_n758), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n899), .B1(new_n917), .B2(new_n918), .ZN(G54));
  NAND2_X1  g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n901), .A2(new_n495), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n495), .B1(new_n901), .B2(new_n920), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n899), .B1(new_n921), .B2(new_n922), .ZN(G60));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n617), .B1(new_n849), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n617), .B(new_n926), .C1(new_n913), .C2(new_n914), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n898), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(G63));
  XNOR2_X1  g744(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n830), .B2(new_n847), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n898), .B1(new_n935), .B2(new_n371), .ZN(new_n936));
  AOI211_X1 g750(.A(new_n640), .B(new_n934), .C1(new_n830), .C2(new_n847), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n818), .A2(new_n809), .A3(new_n823), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n846), .A2(new_n812), .A3(new_n939), .ZN(new_n940));
  AOI22_X1  g754(.A1(new_n940), .A2(new_n808), .B1(new_n827), .B2(new_n809), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n370), .B(new_n368), .C1(new_n941), .C2(new_n934), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n935), .A2(new_n639), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n942), .A2(new_n898), .A3(new_n943), .A4(new_n931), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n938), .A2(new_n944), .ZN(G66));
  OAI21_X1  g759(.A(G953), .B1(new_n513), .B2(new_n562), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n716), .A2(new_n819), .A3(new_n823), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n904), .B1(G898), .B2(new_n241), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G69));
  AOI211_X1 g764(.A(new_n785), .B(new_n667), .C1(new_n622), .C2(new_n820), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n315), .A3(new_n378), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n677), .A2(new_n800), .A3(new_n719), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n780), .A2(new_n792), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n677), .A2(new_n800), .A3(new_n956), .A4(new_n719), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT121), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n241), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n263), .A2(new_n264), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(KEYINPUT122), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n739), .A2(new_n378), .A3(new_n601), .A4(new_n794), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n792), .B(new_n748), .C1(new_n762), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n746), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n800), .A2(new_n719), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n780), .A2(KEYINPUT123), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT123), .B1(new_n780), .B2(new_n968), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n967), .B(new_n241), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n972));
  AOI22_X1  g786(.A1(new_n963), .A2(KEYINPUT122), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n241), .B1(G227), .B2(G900), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT124), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n964), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n964), .B2(new_n973), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  NAND3_X1  g794(.A1(new_n297), .A2(new_n300), .A3(new_n268), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n825), .A2(new_n828), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  AND4_X1   g796(.A1(new_n780), .A2(new_n792), .A3(new_n952), .A4(new_n954), .ZN(new_n983));
  INV_X1    g797(.A(new_n958), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(new_n947), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n980), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n298), .B(KEYINPUT125), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n988), .A2(new_n299), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT126), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  INV_X1    g805(.A(new_n989), .ZN(new_n992));
  AOI211_X1 g806(.A(new_n991), .B(new_n992), .C1(new_n985), .C2(new_n980), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n982), .B(new_n898), .C1(new_n990), .C2(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n967), .B(new_n947), .C1(new_n969), .C2(new_n970), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n995), .A2(new_n996), .A3(new_n980), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n995), .B2(new_n980), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n988), .A2(new_n299), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n994), .A2(new_n1000), .ZN(G57));
endmodule


