//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n192), .A3(new_n195), .A4(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT79), .A2(G107), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT79), .A2(G107), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n198), .B(new_n199), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT79), .A2(G107), .ZN(new_n206));
  AOI21_X1  g020(.A(G104), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(G104), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT81), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n202), .B(G101), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT82), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n200), .A2(new_n201), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n199), .A2(KEYINPUT3), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n204), .B2(G104), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n213), .A2(new_n214), .B1(new_n208), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G143), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(G143), .B2(new_n219), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n220), .A2(new_n222), .A3(new_n224), .A4(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT81), .B(new_n208), .C1(new_n213), .C2(G104), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n230), .A2(KEYINPUT82), .A3(G101), .A4(new_n202), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n218), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n229), .B1(new_n218), .B2(new_n231), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT12), .B(new_n197), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT83), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n210), .A2(new_n211), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n214), .A2(new_n205), .A3(new_n206), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n216), .A2(new_n208), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n212), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n231), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n229), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n218), .A2(new_n229), .A3(new_n231), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT83), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT12), .A4(new_n197), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n197), .B1(new_n232), .B2(new_n233), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n235), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT10), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n197), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n254));
  XNOR2_X1  g068(.A(G143), .B(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(KEYINPUT0), .B2(G128), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n255), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT0), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT64), .B1(new_n261), .B2(new_n226), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n256), .B1(new_n223), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n254), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n257), .B1(new_n255), .B2(new_n259), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n221), .A2(G146), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n219), .A2(G143), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n262), .B(new_n256), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(KEYINPUT68), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n237), .A2(new_n238), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n212), .A2(KEYINPUT80), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n239), .A2(KEYINPUT4), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n271), .A2(KEYINPUT4), .A3(new_n272), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n218), .A2(KEYINPUT10), .A3(new_n229), .A4(new_n231), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n252), .A2(new_n253), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n250), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G227), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT78), .ZN(new_n281));
  XNOR2_X1  g095(.A(G110), .B(G140), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n277), .A2(new_n283), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n252), .A2(new_n276), .A3(new_n275), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n197), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n285), .A2(G469), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n250), .A2(new_n286), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n277), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n284), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n295), .A2(new_n296), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  OAI21_X1  g115(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT76), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n303), .B(KEYINPUT77), .Z(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G125), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT16), .ZN(new_n311));
  OR3_X1    g125(.A1(new_n309), .A2(KEYINPUT16), .A3(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n219), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n312), .A3(G146), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT69), .A2(G237), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT69), .A2(G237), .ZN(new_n318));
  OAI211_X1 g132(.A(G214), .B(new_n279), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT88), .B(G143), .Z(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(KEYINPUT69), .A2(G237), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT69), .A2(G237), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n221), .A2(KEYINPUT88), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n324), .A2(G214), .A3(new_n279), .A4(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n195), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n316), .B1(KEYINPUT17), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT88), .B(G143), .ZN(new_n329));
  AOI21_X1  g143(.A(G953), .B1(new_n322), .B2(new_n323), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(G214), .ZN(new_n331));
  INV_X1    g145(.A(new_n325), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n319), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G131), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n321), .A2(new_n326), .A3(new_n195), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n328), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT89), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT18), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n321), .A2(new_n326), .A3(new_n195), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(new_n327), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n321), .B(new_n326), .C1(new_n339), .C2(new_n340), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT75), .B1(new_n345), .B2(new_n219), .ZN(new_n346));
  AND4_X1   g160(.A1(KEYINPUT75), .A2(new_n308), .A3(new_n310), .A4(new_n219), .ZN(new_n347));
  OAI22_X1  g161(.A1(new_n346), .A2(new_n347), .B1(new_n219), .B2(new_n345), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G113), .B(G122), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT91), .B(G104), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n338), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n338), .B2(new_n350), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n296), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G475), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT20), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n338), .A2(new_n350), .A3(new_n353), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT19), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n345), .B(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n315), .B1(new_n361), .B2(G146), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n334), .A2(new_n336), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(KEYINPUT90), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT90), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n334), .A2(new_n365), .A3(new_n336), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n364), .A2(new_n366), .B1(new_n343), .B2(new_n349), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n359), .B1(new_n367), .B2(new_n353), .ZN(new_n368));
  NOR2_X1   g182(.A1(G475), .A2(G902), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n358), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT90), .B1(new_n342), .B2(new_n327), .ZN(new_n371));
  INV_X1    g185(.A(new_n315), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n345), .B(KEYINPUT19), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(new_n219), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n366), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n353), .B1(new_n375), .B2(new_n350), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n358), .B(new_n369), .C1(new_n354), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n357), .B1(new_n370), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n301), .A2(new_n380), .A3(G953), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT14), .ZN(new_n383));
  INV_X1    g197(.A(G116), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G122), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n384), .B2(G122), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n383), .B1(new_n384), .B2(G122), .ZN(new_n387));
  OAI21_X1  g201(.A(G107), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G116), .B(G122), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n213), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n221), .A2(G128), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n226), .A2(G143), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT92), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT92), .B1(new_n392), .B2(new_n393), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n188), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n396), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(G134), .A3(new_n394), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n391), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n213), .B(new_n389), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT13), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n393), .B1(new_n392), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT13), .B1(new_n221), .B2(G128), .ZN(new_n404));
  OAI21_X1  g218(.A(G134), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n397), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n382), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n399), .A2(new_n397), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n390), .A3(new_n388), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n406), .A3(new_n381), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n296), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n379), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT67), .ZN(new_n418));
  OR2_X1    g232(.A1(KEYINPUT2), .A2(G113), .ZN(new_n419));
  AND3_X1   g233(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G119), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G116), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n384), .A2(G119), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n418), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(KEYINPUT2), .A2(G113), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT65), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G116), .B(G119), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n432), .A2(KEYINPUT67), .A3(new_n433), .A4(new_n419), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G113), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n384), .A2(G119), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT5), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n240), .A2(new_n435), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n441), .ZN(new_n446));
  INV_X1    g260(.A(new_n439), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n435), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n231), .A3(new_n218), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT8), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n435), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT66), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n422), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n432), .A2(KEYINPUT66), .A3(new_n419), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n455), .A2(new_n456), .A3(new_n426), .ZN(new_n457));
  OAI22_X1  g271(.A1(new_n453), .A2(new_n457), .B1(new_n273), .B2(new_n274), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n218), .A2(new_n444), .A3(new_n435), .A4(new_n231), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n450), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n260), .A2(new_n263), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n229), .A2(new_n309), .ZN(new_n463));
  INV_X1    g277(.A(G224), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(new_n464), .B2(G953), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n463), .ZN(new_n467));
  INV_X1    g281(.A(new_n465), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n452), .A2(new_n460), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n470), .A2(new_n296), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n464), .A2(G953), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT86), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n467), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n458), .A2(new_n459), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n450), .A2(KEYINPUT85), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n460), .A2(KEYINPUT6), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n475), .A2(KEYINPUT6), .A3(new_n476), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n471), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n481), .ZN(new_n483));
  INV_X1    g297(.A(new_n474), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n460), .A2(KEYINPUT6), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n475), .A2(new_n476), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(KEYINPUT6), .A3(new_n476), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n470), .A2(new_n296), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n483), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n471), .A2(new_n479), .A3(new_n481), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(KEYINPUT87), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(G234), .A2(G237), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(G952), .A3(new_n279), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT21), .B(G898), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(G902), .A3(G953), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G214), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n417), .A2(new_n482), .A3(new_n493), .A4(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n306), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n188), .A2(G137), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n191), .A2(G134), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n196), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n228), .B2(new_n227), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n270), .B2(new_n197), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n433), .B1(new_n422), .B2(new_n454), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n427), .A2(new_n434), .B1(new_n512), .B2(new_n456), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT28), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n196), .A2(new_n508), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n461), .A2(new_n197), .B1(new_n516), .B2(new_n229), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n517), .B2(new_n513), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n265), .A2(KEYINPUT68), .A3(new_n268), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT68), .B1(new_n265), .B2(new_n268), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n197), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n510), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n513), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n512), .A2(new_n456), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n435), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n265), .A2(new_n268), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n194), .B2(new_n196), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n525), .B(KEYINPUT71), .C1(new_n527), .C2(new_n510), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n518), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n514), .B1(new_n529), .B2(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n330), .A2(G210), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT27), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(G101), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n521), .A2(KEYINPUT30), .A3(new_n522), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n527), .B2(new_n510), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n525), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n523), .ZN(new_n541));
  INV_X1    g355(.A(new_n534), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n535), .A2(KEYINPUT73), .A3(new_n536), .A4(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n521), .A2(new_n522), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n525), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n547), .B2(new_n523), .ZN(new_n548));
  OR4_X1    g362(.A1(new_n536), .A2(new_n548), .A3(new_n542), .A4(new_n514), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(new_n549), .A3(new_n296), .ZN(new_n550));
  INV_X1    g364(.A(new_n543), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(KEYINPUT29), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT73), .B1(new_n552), .B2(new_n535), .ZN(new_n553));
  OAI21_X1  g367(.A(G472), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n540), .A2(new_n534), .A3(new_n523), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT70), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n540), .A2(new_n557), .A3(new_n534), .A4(new_n523), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(KEYINPUT31), .A3(new_n558), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n555), .A2(KEYINPUT31), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n529), .A2(KEYINPUT28), .ZN(new_n561));
  INV_X1    g375(.A(new_n514), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT72), .B1(new_n563), .B2(new_n542), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT72), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n530), .A2(new_n565), .A3(new_n534), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n559), .B(new_n560), .C1(new_n564), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT32), .ZN(new_n568));
  NOR2_X1   g382(.A1(G472), .A2(G902), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n554), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n380), .B1(G234), .B2(new_n296), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n226), .A2(G119), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n423), .A2(G128), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT24), .B(G110), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(KEYINPUT74), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT23), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT23), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n575), .A2(KEYINPUT74), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n576), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n579), .B1(new_n584), .B2(G110), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(new_n315), .C1(new_n346), .C2(new_n347), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(G110), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n316), .B(new_n587), .C1(new_n577), .C2(new_n578), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT22), .B(G137), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n588), .A3(new_n592), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n296), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n594), .A2(KEYINPUT25), .A3(new_n296), .A4(new_n595), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n574), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n594), .A2(new_n595), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n573), .A2(G902), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n505), .A2(new_n572), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NAND2_X1  g423(.A1(new_n567), .A2(new_n296), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n567), .A2(new_n569), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n613), .A2(new_n306), .A3(new_n606), .ZN(new_n614));
  INV_X1    g428(.A(new_n492), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n481), .B1(new_n471), .B2(new_n479), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n412), .A2(KEYINPUT33), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n412), .A2(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(G478), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n412), .A2(new_n414), .A3(new_n296), .ZN(new_n621));
  NAND2_X1  g435(.A1(G478), .A2(G902), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n379), .ZN(new_n624));
  INV_X1    g438(.A(new_n503), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n617), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n614), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  XOR2_X1   g443(.A(new_n413), .B(new_n415), .Z(new_n630));
  NOR4_X1   g444(.A1(new_n617), .A2(new_n630), .A3(new_n379), .A4(new_n625), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n614), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n204), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NOR2_X1   g449(.A1(new_n613), .A2(new_n306), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n589), .B(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n638), .A2(new_n604), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n600), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT94), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n504), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  OAI21_X1  g459(.A(new_n369), .B1(new_n354), .B2(new_n376), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT20), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n377), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n498), .A2(G900), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n495), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n648), .A2(new_n416), .A3(new_n357), .A4(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(G902), .B1(new_n291), .B2(new_n293), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n298), .B1(new_n652), .B2(new_n295), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n304), .B(new_n651), .C1(new_n653), .C2(new_n290), .ZN(new_n654));
  INV_X1    g468(.A(new_n641), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n502), .B1(new_n491), .B2(new_n492), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n654), .A2(new_n572), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  AOI21_X1  g472(.A(new_n304), .B1(new_n653), .B2(new_n290), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n650), .B(KEYINPUT39), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT40), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n493), .A2(new_n482), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n556), .A2(new_n558), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n534), .B1(new_n523), .B2(new_n547), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n296), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(G472), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n570), .B2(new_n571), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n640), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n379), .A2(new_n416), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n672), .A2(new_n502), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n662), .A2(new_n666), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  AOI22_X1  g491(.A1(new_n647), .A2(new_n377), .B1(G475), .B2(new_n356), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n679));
  INV_X1    g493(.A(new_n650), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n300), .A2(new_n305), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n682), .A2(new_n572), .A3(new_n655), .A4(new_n656), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  AOI22_X1  g498(.A1(new_n250), .A2(new_n286), .B1(new_n292), .B2(new_n284), .ZN(new_n685));
  OAI21_X1  g499(.A(G469), .B1(new_n685), .B2(G902), .ZN(new_n686));
  INV_X1    g500(.A(new_n303), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n297), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n572), .A2(new_n607), .A3(new_n626), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT96), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n690), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n572), .A2(new_n607), .A3(new_n631), .A4(new_n689), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  NAND2_X1  g509(.A1(new_n612), .A2(KEYINPUT32), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n641), .B1(new_n698), .B2(new_n554), .ZN(new_n699));
  INV_X1    g513(.A(new_n656), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n688), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n379), .A2(new_n416), .A3(new_n500), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n699), .A2(new_n703), .A3(KEYINPUT97), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n572), .A2(new_n655), .A3(new_n701), .A4(new_n702), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT97), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT98), .B(G119), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G21));
  OAI21_X1  g524(.A(new_n542), .B1(new_n548), .B2(new_n514), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n559), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT99), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT99), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n559), .A2(new_n714), .A3(new_n711), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n560), .A3(new_n715), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n716), .A2(new_n569), .B1(new_n610), .B2(G472), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT100), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n678), .B2(new_n630), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n379), .A2(KEYINPUT100), .A3(new_n416), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n499), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n717), .A2(new_n701), .A3(new_n721), .A4(new_n607), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NAND4_X1  g537(.A1(new_n717), .A2(new_n701), .A3(new_n673), .A4(new_n681), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  AOI21_X1  g539(.A(new_n502), .B1(new_n493), .B2(new_n482), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n572), .A2(new_n607), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n300), .A2(KEYINPUT101), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT101), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n653), .A2(new_n729), .A3(new_n290), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(new_n687), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n681), .B1(KEYINPUT102), .B2(KEYINPUT42), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n727), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT102), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n572), .A2(new_n607), .A3(new_n726), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n731), .ZN(new_n741));
  INV_X1    g555(.A(new_n738), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n734), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n195), .ZN(G33));
  NOR3_X1   g559(.A1(new_n740), .A2(new_n651), .A3(new_n731), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT103), .B(G134), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G36));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n379), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n678), .A2(KEYINPUT106), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT43), .A4(new_n623), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n379), .B2(new_n679), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n752), .A2(KEYINPUT107), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n613), .A2(new_n673), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n726), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n278), .A2(new_n284), .B1(new_n288), .B2(new_n286), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT104), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n768), .A3(KEYINPUT45), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(G469), .B1(new_n765), .B2(KEYINPUT45), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT46), .B(new_n299), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n771), .B1(new_n767), .B2(new_n769), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(new_n298), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n297), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n687), .A3(new_n660), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n764), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n762), .A2(new_n779), .A3(new_n763), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n760), .B1(new_n758), .B2(new_n757), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT108), .B1(new_n781), .B2(KEYINPUT44), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  NAND2_X1  g599(.A1(new_n776), .A2(new_n687), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n786), .B1(new_n787), .B2(KEYINPUT47), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(KEYINPUT47), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(KEYINPUT47), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n776), .B(new_n687), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n663), .A2(new_n501), .A3(new_n681), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n554), .A2(new_n792), .A3(new_n698), .A4(new_n606), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  NOR3_X1   g609(.A1(new_n606), .A2(new_n304), .A3(new_n502), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n623), .A3(new_n751), .A4(new_n750), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n297), .A2(new_n686), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n797), .A2(KEYINPUT110), .B1(KEYINPUT49), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(KEYINPUT110), .B2(new_n797), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT111), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n798), .A2(KEYINPUT49), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n665), .A3(new_n672), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n606), .B1(new_n698), .B2(new_n554), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n495), .B1(new_n752), .B2(new_n754), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n689), .A2(new_n726), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n279), .A2(G952), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n805), .A2(new_n607), .A3(new_n717), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n812), .B1(new_n813), .B2(new_n701), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n606), .A2(new_n495), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n672), .A2(new_n806), .A3(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n811), .B(new_n814), .C1(new_n624), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n813), .A2(new_n726), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n788), .A2(new_n791), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n297), .A2(new_n686), .A3(new_n304), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n688), .A2(new_n501), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT113), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n813), .A3(new_n665), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n678), .A2(new_n679), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n816), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n806), .A2(new_n673), .A3(new_n717), .A4(new_n805), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n829), .A2(KEYINPUT51), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n817), .B1(new_n822), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n829), .A2(KEYINPUT114), .A3(new_n834), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT114), .B1(new_n829), .B2(new_n834), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n837), .A2(new_n821), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n836), .B1(new_n839), .B2(KEYINPUT51), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n792), .A2(new_n717), .A3(new_n673), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n630), .A2(new_n648), .A3(new_n357), .A4(new_n650), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n659), .A2(new_n726), .A3(new_n843), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n842), .A2(new_n732), .B1(new_n699), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n651), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n727), .A2(new_n846), .A3(new_n732), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n493), .A2(new_n482), .A3(new_n503), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n624), .A2(KEYINPUT112), .B1(new_n416), .B2(new_n678), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT112), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n613), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n607), .A4(new_n659), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n804), .A2(new_n505), .B1(new_n636), .B2(new_n642), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n845), .A2(new_n847), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n690), .A2(new_n694), .A3(new_n722), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n708), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n744), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n303), .B1(new_n300), .B2(KEYINPUT101), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n600), .A2(new_n639), .A3(new_n680), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n656), .A2(new_n719), .A3(new_n720), .A4(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n671), .A2(new_n859), .A3(new_n861), .A4(new_n730), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n683), .A2(new_n657), .A3(new_n862), .A4(new_n724), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT52), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n742), .B1(new_n741), .B2(new_n734), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n740), .A2(new_n731), .A3(new_n738), .A4(new_n733), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n853), .A2(new_n643), .A3(new_n608), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n663), .A2(new_n501), .A3(new_n843), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n572), .A2(new_n871), .A3(new_n659), .A4(new_n655), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n792), .A2(new_n717), .A3(new_n673), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n731), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n870), .A2(new_n746), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n690), .A2(new_n694), .A3(new_n722), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n707), .B2(new_n704), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n869), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n878), .A2(new_n879), .A3(new_n864), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n841), .B1(new_n866), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n858), .A2(new_n865), .A3(KEYINPUT53), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n878), .B2(new_n864), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n883), .A3(KEYINPUT54), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n840), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(G952), .A2(G953), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n803), .B1(new_n885), .B2(new_n886), .ZN(G75));
  AOI21_X1  g701(.A(new_n296), .B1(new_n882), .B2(new_n883), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(G210), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n477), .A2(new_n478), .A3(new_n474), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n489), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT55), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n279), .A2(G952), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  XOR2_X1   g710(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n897));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n889), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n894), .A2(new_n899), .ZN(G51));
  AND2_X1   g714(.A1(new_n888), .A2(new_n774), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n298), .B(KEYINPUT57), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n881), .A2(new_n884), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n294), .B(KEYINPUT117), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n901), .B1(new_n905), .B2(KEYINPUT118), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n907), .A3(new_n904), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n895), .B1(new_n906), .B2(new_n908), .ZN(G54));
  NAND2_X1  g723(.A1(KEYINPUT58), .A2(G475), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT119), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n888), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n368), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n896), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n913), .B2(new_n912), .ZN(G60));
  XNOR2_X1  g729(.A(new_n622), .B(KEYINPUT120), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT59), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n881), .A2(new_n884), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n618), .A2(new_n619), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n895), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n882), .B2(new_n883), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(new_n603), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n638), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n896), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n926), .A2(KEYINPUT61), .A3(new_n896), .A4(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(G66));
  NAND3_X1  g746(.A1(new_n497), .A2(G224), .A3(G953), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n857), .A2(new_n870), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n935), .B2(G953), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n487), .B(new_n488), .C1(G898), .C2(new_n279), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n936), .B(new_n937), .Z(G69));
  NAND4_X1  g752(.A1(new_n804), .A2(new_n656), .A3(new_n719), .A4(new_n720), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n777), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n744), .A2(new_n746), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n794), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n683), .A2(new_n657), .A3(new_n724), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT122), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n683), .A2(new_n657), .A3(new_n946), .A4(new_n724), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n784), .A2(new_n943), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n943), .B1(new_n784), .B2(new_n948), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n942), .B(new_n279), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n537), .A2(new_n539), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT121), .Z(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(new_n373), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(G900), .B2(G953), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT125), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n849), .A2(new_n850), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n661), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n959), .B2(new_n740), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n727), .A2(KEYINPUT123), .A3(new_n661), .A4(new_n958), .ZN(new_n961));
  AOI22_X1  g775(.A1(new_n778), .A2(new_n783), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n948), .A2(new_n676), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n948), .A2(new_n965), .A3(new_n676), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n962), .A2(new_n964), .A3(new_n794), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n279), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT124), .B1(new_n968), .B2(new_n954), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n970));
  INV_X1    g784(.A(new_n954), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n970), .B(new_n971), .C1(new_n967), .C2(new_n279), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n956), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n279), .B1(G227), .B2(G900), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n974), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n956), .B(new_n976), .C1(new_n969), .C2(new_n972), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(G72));
  OAI211_X1 g792(.A(new_n942), .B(new_n934), .C1(new_n949), .C2(new_n950), .ZN(new_n979));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT127), .Z(new_n982));
  AOI211_X1 g796(.A(new_n534), .B(new_n541), .C1(new_n979), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n541), .A2(new_n534), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n967), .A2(new_n935), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n982), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n981), .B1(new_n667), .B2(new_n551), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n882), .B2(new_n883), .ZN(new_n988));
  NOR4_X1   g802(.A1(new_n983), .A2(new_n986), .A3(new_n895), .A4(new_n988), .ZN(G57));
endmodule


