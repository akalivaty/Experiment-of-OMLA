

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761;

  AND2_X1 U354 ( .A1(n414), .A2(n410), .ZN(n409) );
  OR2_X1 U355 ( .A1(n653), .A2(n617), .ZN(n625) );
  NOR2_X1 U356 ( .A1(n654), .A2(n690), .ZN(n616) );
  XNOR2_X1 U357 ( .A(n429), .B(KEYINPUT104), .ZN(n661) );
  INV_X1 U358 ( .A(n668), .ZN(n398) );
  XNOR2_X1 U359 ( .A(n538), .B(n537), .ZN(n588) );
  XNOR2_X1 U360 ( .A(n568), .B(n567), .ZN(n575) );
  NOR2_X1 U361 ( .A1(G953), .A2(G237), .ZN(n530) );
  INV_X2 U362 ( .A(G953), .ZN(n750) );
  NAND2_X1 U363 ( .A1(n333), .A2(n339), .ZN(n648) );
  XNOR2_X1 U364 ( .A(n583), .B(n472), .ZN(n333) );
  NAND2_X1 U365 ( .A1(n378), .A2(n381), .ZN(n615) );
  NAND2_X2 U366 ( .A1(n382), .A2(n384), .ZN(n381) );
  NOR2_X2 U367 ( .A1(n371), .A2(n372), .ZN(n353) );
  NAND2_X1 U368 ( .A1(G234), .A2(G237), .ZN(n518) );
  NAND2_X1 U369 ( .A1(n575), .A2(n673), .ZN(n457) );
  BUF_X1 U370 ( .A(G113), .Z(n446) );
  AND2_X2 U371 ( .A1(n370), .A2(n369), .ZN(n368) );
  XNOR2_X2 U372 ( .A(n447), .B(n458), .ZN(n416) );
  AND2_X2 U373 ( .A1(n380), .A2(n379), .ZN(n378) );
  NOR2_X2 U374 ( .A1(n758), .A2(n760), .ZN(n480) );
  XNOR2_X2 U375 ( .A(n461), .B(n460), .ZN(n760) );
  XNOR2_X2 U376 ( .A(n614), .B(KEYINPUT1), .ZN(n668) );
  XNOR2_X2 U377 ( .A(G469), .B(n557), .ZN(n614) );
  INV_X1 U378 ( .A(G472), .ZN(n354) );
  NAND2_X1 U379 ( .A1(n408), .A2(n412), .ZN(n407) );
  XNOR2_X1 U380 ( .A(n581), .B(n580), .ZN(n598) );
  XOR2_X1 U381 ( .A(KEYINPUT31), .B(n593), .Z(n660) );
  AND2_X1 U382 ( .A1(n478), .A2(n398), .ZN(n663) );
  XNOR2_X1 U383 ( .A(n607), .B(KEYINPUT6), .ZN(n627) );
  XNOR2_X1 U384 ( .A(n732), .B(n731), .ZN(n733) );
  NOR2_X1 U385 ( .A1(n732), .A2(G902), .ZN(n568) );
  OR2_X1 U386 ( .A1(n635), .A2(G902), .ZN(n355) );
  XOR2_X1 U387 ( .A(n720), .B(KEYINPUT59), .Z(n722) );
  XNOR2_X1 U388 ( .A(n404), .B(n402), .ZN(n732) );
  XNOR2_X1 U389 ( .A(n716), .B(n715), .ZN(n717) );
  INV_X1 U390 ( .A(n437), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n562), .B(n405), .ZN(n404) );
  XNOR2_X1 U392 ( .A(n424), .B(n511), .ZN(n385) );
  XNOR2_X1 U393 ( .A(n494), .B(n503), .ZN(n505) );
  XNOR2_X1 U394 ( .A(n502), .B(n501), .ZN(n494) );
  XNOR2_X1 U395 ( .A(n508), .B(G134), .ZN(n542) );
  XNOR2_X1 U396 ( .A(n506), .B(G122), .ZN(n493) );
  OR2_X1 U397 ( .A1(G237), .A2(G902), .ZN(n515) );
  XOR2_X1 U398 ( .A(KEYINPUT72), .B(KEYINPUT16), .Z(n506) );
  XOR2_X1 U399 ( .A(KEYINPUT15), .B(G902), .Z(n547) );
  NAND2_X1 U400 ( .A1(n365), .A2(n367), .ZN(n335) );
  NAND2_X1 U401 ( .A1(n365), .A2(n367), .ZN(n730) );
  XNOR2_X2 U402 ( .A(n553), .B(n554), .ZN(n570) );
  OR2_X1 U403 ( .A1(n483), .A2(n547), .ZN(n438) );
  XNOR2_X1 U404 ( .A(n663), .B(KEYINPUT80), .ZN(n477) );
  XNOR2_X1 U405 ( .A(n514), .B(n484), .ZN(n483) );
  INV_X1 U406 ( .A(KEYINPUT87), .ZN(n484) );
  NOR2_X1 U407 ( .A1(n620), .A2(n336), .ZN(n437) );
  NAND2_X1 U408 ( .A1(n563), .A2(G221), .ZN(n405) );
  INV_X1 U409 ( .A(KEYINPUT97), .ZN(n441) );
  INV_X1 U410 ( .A(KEYINPUT17), .ZN(n426) );
  INV_X1 U411 ( .A(n666), .ZN(n413) );
  INV_X1 U412 ( .A(KEYINPUT79), .ZN(n412) );
  INV_X1 U413 ( .A(KEYINPUT48), .ZN(n458) );
  NOR2_X1 U414 ( .A1(n477), .A2(n625), .ZN(n459) );
  XNOR2_X1 U415 ( .A(n507), .B(n500), .ZN(n482) );
  XOR2_X1 U416 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n500) );
  XNOR2_X1 U417 ( .A(n512), .B(G125), .ZN(n526) );
  INV_X1 U418 ( .A(G146), .ZN(n512) );
  XOR2_X1 U419 ( .A(G101), .B(KEYINPUT67), .Z(n507) );
  XNOR2_X1 U420 ( .A(n499), .B(n542), .ZN(n748) );
  XNOR2_X1 U421 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U422 ( .A(G131), .B(KEYINPUT4), .Z(n498) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n683) );
  INV_X1 U424 ( .A(KEYINPUT41), .ZN(n363) );
  NOR2_X1 U425 ( .A1(n688), .A2(n620), .ZN(n362) );
  NOR2_X1 U426 ( .A1(n457), .A2(n614), .ZN(n605) );
  XNOR2_X1 U427 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n554) );
  XOR2_X1 U428 ( .A(G119), .B(G110), .Z(n496) );
  INV_X1 U429 ( .A(KEYINPUT91), .ZN(n462) );
  XNOR2_X1 U430 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U431 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n560) );
  AND2_X1 U432 ( .A1(n360), .A2(n341), .ZN(n352) );
  XNOR2_X1 U433 ( .A(n543), .B(n406), .ZN(n563) );
  INV_X1 U434 ( .A(KEYINPUT8), .ZN(n406) );
  XNOR2_X1 U435 ( .A(n540), .B(n433), .ZN(n432) );
  XNOR2_X1 U436 ( .A(KEYINPUT103), .B(KEYINPUT7), .ZN(n433) );
  XNOR2_X1 U437 ( .A(G116), .B(G122), .ZN(n540) );
  XNOR2_X1 U438 ( .A(n539), .B(KEYINPUT102), .ZN(n431) );
  XNOR2_X1 U439 ( .A(G107), .B(KEYINPUT9), .ZN(n539) );
  XOR2_X1 U440 ( .A(KEYINPUT99), .B(G104), .Z(n528) );
  XNOR2_X1 U441 ( .A(G143), .B(G131), .ZN(n527) );
  XOR2_X1 U442 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n532) );
  XNOR2_X1 U443 ( .A(n526), .B(n463), .ZN(n747) );
  XNOR2_X1 U444 ( .A(G140), .B(KEYINPUT10), .ZN(n463) );
  XNOR2_X1 U445 ( .A(n737), .B(n507), .ZN(n424) );
  XNOR2_X1 U446 ( .A(n748), .B(G146), .ZN(n556) );
  NAND2_X1 U447 ( .A1(n393), .A2(n392), .ZN(n704) );
  NAND2_X1 U448 ( .A1(n400), .A2(KEYINPUT33), .ZN(n392) );
  NAND2_X1 U449 ( .A1(n396), .A2(n394), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n422), .B(n624), .ZN(n633) );
  NAND2_X1 U451 ( .A1(n358), .A2(n357), .ZN(n629) );
  NOR2_X1 U452 ( .A1(n655), .A2(n620), .ZN(n357) );
  XNOR2_X1 U453 ( .A(n481), .B(n359), .ZN(n358) );
  INV_X1 U454 ( .A(KEYINPUT108), .ZN(n359) );
  NOR2_X1 U455 ( .A1(n334), .A2(n425), .ZN(n383) );
  NOR2_X1 U456 ( .A1(n430), .A2(n614), .ZN(n621) );
  XNOR2_X1 U457 ( .A(n443), .B(n340), .ZN(n430) );
  NAND2_X1 U458 ( .A1(n671), .A2(n626), .ZN(n443) );
  XNOR2_X1 U459 ( .A(n474), .B(n473), .ZN(n737) );
  INV_X1 U460 ( .A(G110), .ZN(n473) );
  XNOR2_X1 U461 ( .A(G107), .B(G104), .ZN(n474) );
  NOR2_X1 U462 ( .A1(G952), .A2(n750), .ZN(n736) );
  XNOR2_X1 U463 ( .A(n492), .B(n714), .ZN(n491) );
  INV_X1 U464 ( .A(KEYINPUT47), .ZN(n349) );
  INV_X1 U465 ( .A(KEYINPUT84), .ZN(n485) );
  INV_X1 U466 ( .A(KEYINPUT82), .ZN(n468) );
  NAND2_X1 U467 ( .A1(n685), .A2(n684), .ZN(n689) );
  XOR2_X1 U468 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n510) );
  XNOR2_X1 U469 ( .A(n513), .B(n387), .ZN(n386) );
  XNOR2_X1 U470 ( .A(n526), .B(n388), .ZN(n387) );
  XNOR2_X1 U471 ( .A(n426), .B(n389), .ZN(n388) );
  AND2_X1 U472 ( .A1(n411), .A2(n665), .ZN(n410) );
  NAND2_X1 U473 ( .A1(n413), .A2(n412), .ZN(n411) );
  NAND2_X1 U474 ( .A1(n398), .A2(n397), .ZN(n396) );
  NAND2_X1 U475 ( .A1(n627), .A2(n399), .ZN(n397) );
  INV_X1 U476 ( .A(KEYINPUT33), .ZN(n395) );
  XNOR2_X1 U477 ( .A(KEYINPUT86), .B(KEYINPUT0), .ZN(n524) );
  NOR2_X1 U478 ( .A1(n375), .A2(n517), .ZN(n374) );
  NOR2_X1 U479 ( .A1(n334), .A2(n376), .ZN(n375) );
  INV_X1 U480 ( .A(n438), .ZN(n376) );
  XNOR2_X1 U481 ( .A(n556), .B(n356), .ZN(n635) );
  XNOR2_X1 U482 ( .A(n504), .B(n442), .ZN(n356) );
  XNOR2_X1 U483 ( .A(n482), .B(n495), .ZN(n442) );
  INV_X1 U484 ( .A(KEYINPUT45), .ZN(n452) );
  XNOR2_X1 U485 ( .A(n577), .B(n578), .ZN(n456) );
  XNOR2_X1 U486 ( .A(n606), .B(n421), .ZN(n420) );
  INV_X1 U487 ( .A(KEYINPUT74), .ZN(n421) );
  NAND2_X1 U488 ( .A1(n595), .A2(n487), .ZN(n451) );
  XNOR2_X1 U489 ( .A(n448), .B(KEYINPUT95), .ZN(n595) );
  NAND2_X1 U490 ( .A1(n594), .A2(n605), .ZN(n448) );
  XNOR2_X1 U491 ( .A(n635), .B(KEYINPUT62), .ZN(n636) );
  XNOR2_X1 U492 ( .A(n747), .B(n403), .ZN(n402) );
  XNOR2_X1 U493 ( .A(n496), .B(n462), .ZN(n403) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n541) );
  XNOR2_X1 U495 ( .A(n535), .B(n534), .ZN(n720) );
  XNOR2_X1 U496 ( .A(n556), .B(n434), .ZN(n716) );
  XNOR2_X1 U497 ( .A(n555), .B(G140), .ZN(n435) );
  BUF_X1 U498 ( .A(G953), .Z(n427) );
  XNOR2_X1 U499 ( .A(n622), .B(n444), .ZN(n758) );
  XNOR2_X1 U500 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n444) );
  INV_X1 U501 ( .A(KEYINPUT40), .ZN(n460) );
  NOR2_X1 U502 ( .A1(n629), .A2(n631), .ZN(n628) );
  XNOR2_X1 U503 ( .A(n574), .B(KEYINPUT32), .ZN(n486) );
  INV_X1 U504 ( .A(KEYINPUT65), .ZN(n574) );
  NAND2_X1 U505 ( .A1(n621), .A2(n351), .ZN(n654) );
  INV_X1 U506 ( .A(KEYINPUT107), .ZN(n472) );
  INV_X1 U507 ( .A(n451), .ZN(n644) );
  INV_X1 U508 ( .A(KEYINPUT56), .ZN(n488) );
  INV_X1 U509 ( .A(n736), .ZN(n490) );
  INV_X1 U510 ( .A(G122), .ZN(n391) );
  AND2_X1 U511 ( .A1(n483), .A2(n547), .ZN(n336) );
  NAND2_X1 U512 ( .A1(n634), .A2(n476), .ZN(n337) );
  INV_X1 U513 ( .A(n671), .ZN(n487) );
  XOR2_X1 U514 ( .A(KEYINPUT88), .B(n516), .Z(n620) );
  XOR2_X1 U515 ( .A(n344), .B(KEYINPUT83), .Z(n338) );
  AND2_X1 U516 ( .A1(n487), .A2(n569), .ZN(n339) );
  INV_X1 U517 ( .A(n428), .ZN(n690) );
  OR2_X1 U518 ( .A1(n661), .A2(n657), .ZN(n428) );
  XOR2_X1 U519 ( .A(KEYINPUT109), .B(KEYINPUT28), .Z(n340) );
  AND2_X1 U520 ( .A1(n547), .A2(KEYINPUT64), .ZN(n341) );
  NAND2_X1 U521 ( .A1(n667), .A2(n476), .ZN(n367) );
  NAND2_X1 U522 ( .A1(n368), .A2(n360), .ZN(n667) );
  NAND2_X1 U523 ( .A1(n407), .A2(KEYINPUT2), .ZN(n372) );
  INV_X1 U524 ( .A(n409), .ZN(n371) );
  XNOR2_X1 U525 ( .A(n453), .B(KEYINPUT45), .ZN(n342) );
  XNOR2_X1 U526 ( .A(n599), .B(KEYINPUT68), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n759), .A2(n648), .ZN(n343) );
  XNOR2_X1 U528 ( .A(n343), .B(n485), .ZN(n344) );
  XNOR2_X1 U529 ( .A(n445), .B(n485), .ZN(n600) );
  INV_X1 U530 ( .A(n457), .ZN(n401) );
  NOR2_X1 U531 ( .A1(n457), .A2(KEYINPUT33), .ZN(n399) );
  BUF_X1 U532 ( .A(n423), .Z(n345) );
  BUF_X1 U533 ( .A(n711), .Z(n346) );
  NOR2_X1 U534 ( .A1(KEYINPUT44), .A2(n598), .ZN(n599) );
  NAND2_X1 U535 ( .A1(n668), .A2(n395), .ZN(n394) );
  XNOR2_X1 U536 ( .A(n347), .B(n348), .ZN(n534) );
  XNOR2_X1 U537 ( .A(n533), .B(KEYINPUT11), .ZN(n347) );
  XOR2_X1 U538 ( .A(n446), .B(G122), .Z(n348) );
  XNOR2_X1 U539 ( .A(n349), .B(n616), .ZN(n617) );
  XNOR2_X1 U540 ( .A(n453), .B(n452), .ZN(n350) );
  NAND2_X1 U541 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U542 ( .A1(n759), .A2(n648), .ZN(n445) );
  BUF_X1 U543 ( .A(n576), .Z(n592) );
  NAND2_X1 U544 ( .A1(n381), .A2(n378), .ZN(n351) );
  NAND2_X1 U545 ( .A1(n342), .A2(n353), .ZN(n360) );
  AND2_X2 U546 ( .A1(n373), .A2(n383), .ZN(n382) );
  INV_X1 U547 ( .A(n436), .ZN(n384) );
  NAND2_X1 U548 ( .A1(n335), .A2(G210), .ZN(n492) );
  INV_X1 U549 ( .A(n592), .ZN(n594) );
  AND2_X2 U550 ( .A1(n711), .A2(n483), .ZN(n436) );
  NAND2_X1 U551 ( .A1(n352), .A2(n368), .ZN(n366) );
  XNOR2_X2 U552 ( .A(n355), .B(n354), .ZN(n607) );
  NOR2_X1 U553 ( .A1(n436), .A2(n336), .ZN(n439) );
  XNOR2_X2 U554 ( .A(n361), .B(n385), .ZN(n711) );
  XNOR2_X2 U555 ( .A(n423), .B(n386), .ZN(n361) );
  NAND2_X1 U556 ( .A1(n685), .A2(n362), .ZN(n364) );
  XNOR2_X2 U557 ( .A(n631), .B(n619), .ZN(n685) );
  AND2_X2 U558 ( .A1(n366), .A2(n337), .ZN(n365) );
  OR2_X2 U559 ( .A1(n711), .A2(n438), .ZN(n373) );
  NAND2_X1 U560 ( .A1(n711), .A2(n437), .ZN(n377) );
  NAND2_X1 U561 ( .A1(n749), .A2(n475), .ZN(n369) );
  NAND2_X1 U562 ( .A1(n350), .A2(n475), .ZN(n370) );
  NAND2_X1 U563 ( .A1(n409), .A2(n407), .ZN(n749) );
  NAND2_X2 U564 ( .A1(n439), .A2(n373), .ZN(n631) );
  NAND2_X1 U565 ( .A1(n377), .A2(n374), .ZN(n379) );
  NAND2_X1 U566 ( .A1(n615), .A2(n523), .ZN(n525) );
  NAND2_X1 U567 ( .A1(n436), .A2(n425), .ZN(n380) );
  XNOR2_X2 U568 ( .A(n505), .B(n493), .ZN(n423) );
  INV_X1 U569 ( .A(KEYINPUT4), .ZN(n389) );
  NAND2_X1 U570 ( .A1(n600), .A2(n390), .ZN(n582) );
  INV_X1 U571 ( .A(n598), .ZN(n390) );
  XNOR2_X1 U572 ( .A(n598), .B(n391), .ZN(G24) );
  NOR2_X1 U573 ( .A1(n668), .A2(n457), .ZN(n591) );
  NAND2_X1 U574 ( .A1(n627), .A2(n401), .ZN(n400) );
  XNOR2_X2 U575 ( .A(G143), .B(G128), .ZN(n508) );
  INV_X1 U576 ( .A(n416), .ZN(n408) );
  NAND2_X1 U577 ( .A1(n416), .A2(n415), .ZN(n414) );
  AND2_X1 U578 ( .A1(n666), .A2(KEYINPUT79), .ZN(n415) );
  NAND2_X1 U579 ( .A1(n417), .A2(n420), .ZN(n422) );
  NOR2_X1 U580 ( .A1(n609), .A2(n418), .ZN(n417) );
  INV_X1 U581 ( .A(n685), .ZN(n418) );
  NOR2_X1 U582 ( .A1(n609), .A2(n419), .ZN(n623) );
  INV_X1 U583 ( .A(n420), .ZN(n419) );
  XNOR2_X1 U584 ( .A(n345), .B(G101), .ZN(n738) );
  XNOR2_X1 U585 ( .A(n424), .B(n435), .ZN(n434) );
  INV_X1 U586 ( .A(n517), .ZN(n425) );
  NAND2_X1 U587 ( .A1(n627), .A2(n626), .ZN(n481) );
  NOR2_X1 U588 ( .A1(n590), .A2(n589), .ZN(n429) );
  XNOR2_X1 U589 ( .A(n721), .B(n722), .ZN(n723) );
  AND2_X1 U590 ( .A1(n440), .A2(n428), .ZN(n596) );
  XNOR2_X1 U591 ( .A(n449), .B(n441), .ZN(n440) );
  NOR2_X2 U592 ( .A1(n592), .A2(n678), .ZN(n593) );
  XNOR2_X2 U593 ( .A(n525), .B(n524), .ZN(n576) );
  NOR2_X2 U594 ( .A1(n576), .A2(n552), .ZN(n553) );
  XNOR2_X1 U595 ( .A(n469), .B(n468), .ZN(n467) );
  NAND2_X1 U596 ( .A1(n467), .A2(n465), .ZN(n453) );
  NAND2_X1 U597 ( .A1(n470), .A2(n464), .ZN(n469) );
  NAND2_X1 U598 ( .A1(n459), .A2(n479), .ZN(n447) );
  NAND2_X1 U599 ( .A1(n491), .A2(n490), .ZN(n489) );
  XNOR2_X2 U600 ( .A(n573), .B(n486), .ZN(n759) );
  NOR2_X2 U601 ( .A1(n638), .A2(n736), .ZN(n640) );
  NAND2_X1 U602 ( .A1(n451), .A2(n450), .ZN(n449) );
  INV_X1 U603 ( .A(n660), .ZN(n450) );
  XNOR2_X1 U604 ( .A(n454), .B(KEYINPUT126), .ZN(G66) );
  NOR2_X2 U605 ( .A1(n735), .A2(n736), .ZN(n454) );
  NOR2_X2 U606 ( .A1(n570), .A2(n398), .ZN(n583) );
  NAND2_X1 U607 ( .A1(n338), .A2(n466), .ZN(n465) );
  XNOR2_X1 U608 ( .A(n455), .B(KEYINPUT122), .ZN(G54) );
  NOR2_X2 U609 ( .A1(n719), .A2(n736), .ZN(n455) );
  NAND2_X1 U610 ( .A1(n456), .A2(n579), .ZN(n581) );
  NAND2_X1 U611 ( .A1(n668), .A2(n457), .ZN(n669) );
  NAND2_X1 U612 ( .A1(n633), .A2(n657), .ZN(n461) );
  NAND2_X1 U613 ( .A1(n582), .A2(KEYINPUT44), .ZN(n470) );
  NOR2_X1 U614 ( .A1(n596), .A2(n597), .ZN(n464) );
  INV_X1 U615 ( .A(KEYINPUT2), .ZN(n475) );
  INV_X1 U616 ( .A(KEYINPUT64), .ZN(n476) );
  XNOR2_X1 U617 ( .A(n628), .B(KEYINPUT36), .ZN(n478) );
  XNOR2_X1 U618 ( .A(n480), .B(KEYINPUT46), .ZN(n479) );
  INV_X1 U619 ( .A(n607), .ZN(n671) );
  NAND2_X1 U620 ( .A1(n730), .A2(G475), .ZN(n721) );
  XNOR2_X1 U621 ( .A(n489), .B(n488), .ZN(G51) );
  XNOR2_X1 U622 ( .A(n718), .B(n717), .ZN(n719) );
  AND2_X1 U623 ( .A1(n530), .A2(G210), .ZN(n495) );
  XNOR2_X1 U624 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U625 ( .A(KEYINPUT73), .ZN(n618) );
  XNOR2_X1 U626 ( .A(n618), .B(KEYINPUT38), .ZN(n619) );
  INV_X1 U627 ( .A(KEYINPUT125), .ZN(n731) );
  XNOR2_X1 U628 ( .A(KEYINPUT76), .B(KEYINPUT35), .ZN(n580) );
  XNOR2_X1 U629 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U630 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U631 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U632 ( .A(KEYINPUT69), .B(G137), .ZN(n497) );
  XNOR2_X2 U633 ( .A(G116), .B(G113), .ZN(n502) );
  INV_X1 U634 ( .A(KEYINPUT3), .ZN(n501) );
  XOR2_X1 U635 ( .A(KEYINPUT70), .B(G119), .Z(n503) );
  BUF_X1 U636 ( .A(n505), .Z(n504) );
  INV_X1 U637 ( .A(n508), .ZN(n509) );
  NAND2_X1 U638 ( .A1(G224), .A2(n750), .ZN(n513) );
  NAND2_X1 U639 ( .A1(G210), .A2(n515), .ZN(n514) );
  NAND2_X1 U640 ( .A1(n515), .A2(G214), .ZN(n516) );
  XOR2_X1 U641 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n517) );
  XNOR2_X1 U642 ( .A(n518), .B(KEYINPUT14), .ZN(n520) );
  NAND2_X1 U643 ( .A1(G952), .A2(n520), .ZN(n701) );
  NOR2_X1 U644 ( .A1(n701), .A2(n427), .ZN(n519) );
  XNOR2_X1 U645 ( .A(n519), .B(KEYINPUT89), .ZN(n604) );
  NAND2_X1 U646 ( .A1(G902), .A2(n520), .ZN(n601) );
  INV_X1 U647 ( .A(n601), .ZN(n521) );
  NOR2_X1 U648 ( .A1(G898), .A2(n750), .ZN(n739) );
  NAND2_X1 U649 ( .A1(n521), .A2(n739), .ZN(n522) );
  NAND2_X1 U650 ( .A1(n604), .A2(n522), .ZN(n523) );
  XNOR2_X1 U651 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U652 ( .A(n747), .B(n529), .ZN(n535) );
  NAND2_X1 U653 ( .A1(G214), .A2(n530), .ZN(n531) );
  XNOR2_X1 U654 ( .A(n532), .B(n531), .ZN(n533) );
  NOR2_X1 U655 ( .A1(n720), .A2(G902), .ZN(n538) );
  XOR2_X1 U656 ( .A(G475), .B(KEYINPUT13), .Z(n536) );
  XNOR2_X1 U657 ( .A(KEYINPUT100), .B(n536), .ZN(n537) );
  XOR2_X1 U658 ( .A(n542), .B(n541), .Z(n545) );
  NAND2_X1 U659 ( .A1(G234), .A2(n750), .ZN(n543) );
  NAND2_X1 U660 ( .A1(G217), .A2(n563), .ZN(n544) );
  XNOR2_X1 U661 ( .A(n545), .B(n544), .ZN(n726) );
  NOR2_X1 U662 ( .A1(n726), .A2(G902), .ZN(n546) );
  XNOR2_X1 U663 ( .A(n546), .B(G478), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n588), .A2(n589), .ZN(n688) );
  INV_X1 U665 ( .A(n688), .ZN(n551) );
  XOR2_X1 U666 ( .A(KEYINPUT21), .B(KEYINPUT94), .Z(n550) );
  INV_X1 U667 ( .A(n547), .ZN(n634) );
  NAND2_X1 U668 ( .A1(G234), .A2(n634), .ZN(n548) );
  XNOR2_X1 U669 ( .A(KEYINPUT20), .B(n548), .ZN(n564) );
  NAND2_X1 U670 ( .A1(G221), .A2(n564), .ZN(n549) );
  XNOR2_X1 U671 ( .A(n550), .B(n549), .ZN(n673) );
  NAND2_X1 U672 ( .A1(n551), .A2(n673), .ZN(n552) );
  NAND2_X1 U673 ( .A1(G227), .A2(n750), .ZN(n555) );
  NOR2_X1 U674 ( .A1(G902), .A2(n716), .ZN(n557) );
  XOR2_X1 U675 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n559) );
  XNOR2_X1 U676 ( .A(G128), .B(G137), .ZN(n558) );
  XNOR2_X1 U677 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U678 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n566) );
  NAND2_X1 U679 ( .A1(G217), .A2(n564), .ZN(n565) );
  XNOR2_X1 U680 ( .A(n566), .B(n565), .ZN(n567) );
  INV_X1 U681 ( .A(n575), .ZN(n569) );
  XOR2_X1 U682 ( .A(n569), .B(KEYINPUT105), .Z(n584) );
  INV_X1 U683 ( .A(n584), .ZN(n672) );
  NOR2_X1 U684 ( .A1(n570), .A2(n672), .ZN(n572) );
  NOR2_X1 U685 ( .A1(n668), .A2(n627), .ZN(n571) );
  NOR2_X1 U686 ( .A1(n588), .A2(n589), .ZN(n610) );
  XOR2_X1 U687 ( .A(n610), .B(KEYINPUT77), .Z(n579) );
  XOR2_X1 U688 ( .A(KEYINPUT34), .B(KEYINPUT78), .Z(n578) );
  NAND2_X1 U689 ( .A1(n704), .A2(n594), .ZN(n577) );
  BUF_X1 U690 ( .A(n583), .Z(n586) );
  NOR2_X1 U691 ( .A1(n627), .A2(n584), .ZN(n585) );
  NAND2_X1 U692 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U693 ( .A(KEYINPUT106), .B(n587), .ZN(n761) );
  INV_X1 U694 ( .A(n761), .ZN(n597) );
  XNOR2_X1 U695 ( .A(KEYINPUT101), .B(n588), .ZN(n590) );
  NAND2_X1 U696 ( .A1(n589), .A2(n590), .ZN(n655) );
  INV_X1 U697 ( .A(n655), .ZN(n657) );
  NAND2_X1 U698 ( .A1(n671), .A2(n591), .ZN(n678) );
  NOR2_X1 U699 ( .A1(G900), .A2(n601), .ZN(n602) );
  NAND2_X1 U700 ( .A1(n427), .A2(n602), .ZN(n603) );
  NAND2_X1 U701 ( .A1(n604), .A2(n603), .ZN(n612) );
  NAND2_X1 U702 ( .A1(n605), .A2(n612), .ZN(n606) );
  NOR2_X1 U703 ( .A1(n620), .A2(n607), .ZN(n608) );
  XOR2_X1 U704 ( .A(KEYINPUT30), .B(n608), .Z(n609) );
  NAND2_X1 U705 ( .A1(n623), .A2(n610), .ZN(n611) );
  NOR2_X1 U706 ( .A1(n631), .A2(n611), .ZN(n653) );
  NAND2_X1 U707 ( .A1(n673), .A2(n612), .ZN(n613) );
  NOR2_X1 U708 ( .A1(n575), .A2(n613), .ZN(n626) );
  INV_X1 U709 ( .A(n620), .ZN(n684) );
  INV_X1 U710 ( .A(n683), .ZN(n703) );
  AND2_X1 U711 ( .A1(n703), .A2(n621), .ZN(n622) );
  XOR2_X1 U712 ( .A(KEYINPUT81), .B(KEYINPUT39), .Z(n624) );
  OR2_X1 U713 ( .A1(n398), .A2(n629), .ZN(n630) );
  XNOR2_X1 U714 ( .A(n630), .B(KEYINPUT43), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n666) );
  NAND2_X1 U716 ( .A1(n633), .A2(n661), .ZN(n665) );
  NAND2_X1 U717 ( .A1(n730), .A2(G472), .ZN(n637) );
  XNOR2_X1 U718 ( .A(KEYINPUT63), .B(KEYINPUT111), .ZN(n639) );
  XNOR2_X1 U719 ( .A(n640), .B(n639), .ZN(G57) );
  XOR2_X1 U720 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n642) );
  NAND2_X1 U721 ( .A1(n644), .A2(n657), .ZN(n641) );
  XNOR2_X1 U722 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U723 ( .A(G104), .B(n643), .ZN(G6) );
  XOR2_X1 U724 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n646) );
  NAND2_X1 U725 ( .A1(n644), .A2(n661), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U727 ( .A(G107), .B(n647), .ZN(G9) );
  XNOR2_X1 U728 ( .A(n648), .B(G110), .ZN(G12) );
  INV_X1 U729 ( .A(n661), .ZN(n649) );
  NOR2_X1 U730 ( .A1(n649), .A2(n654), .ZN(n651) );
  XNOR2_X1 U731 ( .A(KEYINPUT29), .B(KEYINPUT114), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U733 ( .A(G128), .B(n652), .ZN(G30) );
  XOR2_X1 U734 ( .A(G143), .B(n653), .Z(G45) );
  NOR2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U736 ( .A(G146), .B(n656), .Z(G48) );
  XOR2_X1 U737 ( .A(n446), .B(KEYINPUT115), .Z(n659) );
  NAND2_X1 U738 ( .A1(n660), .A2(n657), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n659), .B(n658), .ZN(G15) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n662), .B(G116), .ZN(G18) );
  XNOR2_X1 U742 ( .A(n663), .B(G125), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n664), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U744 ( .A(G134), .B(n665), .ZN(G36) );
  XNOR2_X1 U745 ( .A(G140), .B(n666), .ZN(G42) );
  BUF_X1 U746 ( .A(n667), .Z(n709) );
  XOR2_X1 U747 ( .A(KEYINPUT50), .B(n669), .Z(n670) );
  NOR2_X1 U748 ( .A1(n671), .A2(n670), .ZN(n677) );
  NOR2_X1 U749 ( .A1(n673), .A2(n672), .ZN(n675) );
  XNOR2_X1 U750 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n674) );
  XNOR2_X1 U751 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U753 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U754 ( .A(n680), .B(KEYINPUT117), .ZN(n681) );
  XOR2_X1 U755 ( .A(KEYINPUT51), .B(n681), .Z(n682) );
  NOR2_X1 U756 ( .A1(n683), .A2(n682), .ZN(n697) );
  NOR2_X1 U757 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n686), .B(KEYINPUT118), .ZN(n687) );
  NOR2_X1 U759 ( .A1(n688), .A2(n687), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U761 ( .A(KEYINPUT119), .B(n691), .Z(n692) );
  NOR2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n695) );
  INV_X1 U763 ( .A(n704), .ZN(n694) );
  NOR2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U766 ( .A(n698), .B(KEYINPUT120), .ZN(n699) );
  XNOR2_X1 U767 ( .A(KEYINPUT52), .B(n699), .ZN(n700) );
  NOR2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U769 ( .A(n702), .B(KEYINPUT121), .ZN(n706) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n427), .A2(n707), .ZN(n708) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U774 ( .A(KEYINPUT53), .B(n710), .Z(G75) );
  XOR2_X1 U775 ( .A(KEYINPUT85), .B(KEYINPUT55), .Z(n713) );
  XNOR2_X1 U776 ( .A(n346), .B(KEYINPUT54), .ZN(n712) );
  XNOR2_X1 U777 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U778 ( .A1(n730), .A2(G469), .ZN(n718) );
  XOR2_X1 U779 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n715) );
  NOR2_X2 U780 ( .A1(n723), .A2(n736), .ZN(n724) );
  XNOR2_X1 U781 ( .A(n724), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U782 ( .A1(G478), .A2(n335), .ZN(n728) );
  XOR2_X1 U783 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n725) );
  NOR2_X1 U784 ( .A1(n736), .A2(n729), .ZN(G63) );
  NAND2_X1 U785 ( .A1(n335), .A2(G217), .ZN(n734) );
  XNOR2_X1 U786 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n737), .B(n738), .ZN(n740) );
  NOR2_X1 U788 ( .A1(n740), .A2(n739), .ZN(n746) );
  NAND2_X1 U789 ( .A1(n427), .A2(G224), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n741), .B(KEYINPUT61), .ZN(n742) );
  NAND2_X1 U791 ( .A1(n742), .A2(G898), .ZN(n744) );
  OR2_X1 U792 ( .A1(n427), .A2(n350), .ZN(n743) );
  NAND2_X1 U793 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(G69) );
  XNOR2_X1 U795 ( .A(n748), .B(n747), .ZN(n752) );
  XNOR2_X1 U796 ( .A(n749), .B(n752), .ZN(n751) );
  NAND2_X1 U797 ( .A1(n751), .A2(n750), .ZN(n757) );
  XNOR2_X1 U798 ( .A(G227), .B(n752), .ZN(n753) );
  NAND2_X1 U799 ( .A1(n753), .A2(G900), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n754), .A2(n427), .ZN(n755) );
  XOR2_X1 U801 ( .A(KEYINPUT127), .B(n755), .Z(n756) );
  NAND2_X1 U802 ( .A1(n757), .A2(n756), .ZN(G72) );
  XOR2_X1 U803 ( .A(n758), .B(G137), .Z(G39) );
  XNOR2_X1 U804 ( .A(G119), .B(n759), .ZN(G21) );
  XOR2_X1 U805 ( .A(G131), .B(n760), .Z(G33) );
  XNOR2_X1 U806 ( .A(G101), .B(n761), .ZN(G3) );
endmodule

