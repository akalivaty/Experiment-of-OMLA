

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725;

  XNOR2_X1 U363 ( .A(n430), .B(n366), .ZN(n613) );
  NAND2_X2 U364 ( .A1(n389), .A2(n387), .ZN(n557) );
  XNOR2_X2 U365 ( .A(n557), .B(KEYINPUT19), .ZN(n560) );
  INV_X1 U366 ( .A(G953), .ZN(n713) );
  BUF_X1 U367 ( .A(G143), .Z(n367) );
  AND2_X2 U368 ( .A1(n353), .A2(n352), .ZN(n351) );
  OR2_X2 U369 ( .A1(n591), .A2(G902), .ZN(n383) );
  XNOR2_X2 U370 ( .A(n535), .B(KEYINPUT39), .ZN(n583) );
  OR2_X2 U371 ( .A1(n565), .A2(n537), .ZN(n535) );
  NAND2_X2 U372 ( .A1(n347), .A2(n393), .ZN(n346) );
  XNOR2_X2 U373 ( .A(n346), .B(n344), .ZN(n508) );
  XNOR2_X2 U374 ( .A(n459), .B(n458), .ZN(n534) );
  OR2_X2 U375 ( .A1(n680), .A2(n590), .ZN(n459) );
  NAND2_X2 U376 ( .A1(n370), .A2(n368), .ZN(n379) );
  NAND2_X1 U377 ( .A1(n375), .A2(n374), .ZN(n677) );
  NOR2_X1 U378 ( .A1(n638), .A2(n469), .ZN(n360) );
  XNOR2_X1 U379 ( .A(n556), .B(KEYINPUT106), .ZN(n577) );
  NAND2_X1 U380 ( .A1(n567), .A2(n388), .ZN(n387) );
  AND2_X1 U381 ( .A1(n391), .A2(n390), .ZN(n389) );
  XNOR2_X1 U382 ( .A(n544), .B(n409), .ZN(n410) );
  XNOR2_X1 U383 ( .A(n383), .B(n382), .ZN(n544) );
  XNOR2_X1 U384 ( .A(n434), .B(n701), .ZN(n454) );
  OR2_X2 U385 ( .A1(n611), .A2(G902), .ZN(n442) );
  XNOR2_X1 U386 ( .A(n408), .B(G469), .ZN(n382) );
  XNOR2_X1 U387 ( .A(n355), .B(n522), .ZN(n693) );
  NOR2_X1 U388 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U389 ( .A(n515), .B(KEYINPUT99), .ZN(n626) );
  NAND2_X1 U390 ( .A1(n379), .A2(G472), .ZN(n386) );
  INV_X1 U391 ( .A(KEYINPUT44), .ZN(n354) );
  NOR2_X1 U392 ( .A1(n722), .A2(n354), .ZN(n349) );
  XNOR2_X1 U393 ( .A(n677), .B(KEYINPUT85), .ZN(n559) );
  XOR2_X1 U394 ( .A(G137), .B(KEYINPUT67), .Z(n418) );
  XNOR2_X1 U395 ( .A(n417), .B(n447), .ZN(n475) );
  XNOR2_X1 U396 ( .A(G113), .B(n367), .ZN(n470) );
  XNOR2_X1 U397 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n446) );
  INV_X1 U398 ( .A(n656), .ZN(n362) );
  XNOR2_X1 U399 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U400 ( .A(KEYINPUT3), .B(G119), .Z(n432) );
  XNOR2_X1 U401 ( .A(G116), .B(G113), .ZN(n431) );
  XOR2_X1 U402 ( .A(G104), .B(KEYINPUT88), .Z(n404) );
  XNOR2_X1 U403 ( .A(n422), .B(n421), .ZN(n423) );
  INV_X1 U404 ( .A(KEYINPUT23), .ZN(n421) );
  XNOR2_X1 U405 ( .A(G119), .B(G128), .ZN(n422) );
  XNOR2_X1 U406 ( .A(n475), .B(n418), .ZN(n712) );
  XNOR2_X1 U407 ( .A(G122), .B(G107), .ZN(n488) );
  AND2_X1 U408 ( .A1(n378), .A2(n410), .ZN(n377) );
  OR2_X1 U409 ( .A1(n555), .A2(n554), .ZN(n556) );
  OR2_X1 U410 ( .A1(n544), .A2(n617), .ZN(n523) );
  XNOR2_X1 U411 ( .A(n429), .B(KEYINPUT25), .ZN(n366) );
  OR2_X1 U412 ( .A1(n689), .A2(G902), .ZN(n430) );
  NAND2_X1 U413 ( .A1(n373), .A2(n369), .ZN(n368) );
  NAND2_X1 U414 ( .A1(n612), .A2(n587), .ZN(n370) );
  NOR2_X1 U415 ( .A1(n392), .A2(n461), .ZN(n388) );
  XNOR2_X1 U416 ( .A(G137), .B(KEYINPUT5), .ZN(n436) );
  XNOR2_X1 U417 ( .A(n411), .B(G902), .ZN(n590) );
  XNOR2_X1 U418 ( .A(G107), .B(G140), .ZN(n398) );
  XNOR2_X1 U419 ( .A(n397), .B(n435), .ZN(n401) );
  NAND2_X1 U420 ( .A1(n350), .A2(n349), .ZN(n348) );
  AND2_X1 U421 ( .A1(n571), .A2(n396), .ZN(n572) );
  INV_X1 U422 ( .A(KEYINPUT46), .ZN(n548) );
  BUF_X1 U423 ( .A(n638), .Z(n645) );
  XNOR2_X1 U424 ( .A(n581), .B(n343), .ZN(n537) );
  XNOR2_X1 U425 ( .A(n444), .B(KEYINPUT33), .ZN(n638) );
  AND2_X1 U426 ( .A1(n514), .A2(n551), .ZN(n444) );
  XNOR2_X1 U427 ( .A(n380), .B(KEYINPUT75), .ZN(n514) );
  NAND2_X1 U428 ( .A1(n410), .A2(n381), .ZN(n380) );
  INV_X1 U429 ( .A(n617), .ZN(n381) );
  INV_X1 U430 ( .A(G128), .ZN(n402) );
  AND2_X1 U431 ( .A1(n589), .A2(n372), .ZN(n369) );
  AND2_X1 U432 ( .A1(n590), .A2(n588), .ZN(n372) );
  XOR2_X1 U433 ( .A(G122), .B(G104), .Z(n471) );
  XNOR2_X1 U434 ( .A(n454), .B(n453), .ZN(n680) );
  NAND2_X1 U435 ( .A1(n373), .A2(n589), .ZN(n612) );
  XNOR2_X1 U436 ( .A(n342), .B(n712), .ZN(n427) );
  XOR2_X1 U437 ( .A(n600), .B(KEYINPUT59), .Z(n601) );
  XNOR2_X1 U438 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U439 ( .A(n536), .B(KEYINPUT40), .ZN(n724) );
  AND2_X1 U440 ( .A1(n583), .A2(n670), .ZN(n536) );
  AND2_X1 U441 ( .A1(n376), .A2(n377), .ZN(n375) );
  AND2_X1 U442 ( .A1(n503), .A2(n504), .ZN(n393) );
  XNOR2_X1 U443 ( .A(n516), .B(KEYINPUT31), .ZN(n674) );
  XNOR2_X1 U444 ( .A(n365), .B(n364), .ZN(n659) );
  INV_X1 U445 ( .A(KEYINPUT98), .ZN(n364) );
  INV_X1 U446 ( .A(n692), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n345), .ZN(n358) );
  OR2_X1 U448 ( .A1(n674), .A2(n659), .ZN(n340) );
  OR2_X1 U449 ( .A1(n558), .A2(KEYINPUT36), .ZN(n341) );
  XOR2_X1 U450 ( .A(n424), .B(n423), .Z(n342) );
  OR2_X1 U451 ( .A1(n507), .A2(n506), .ZN(n663) );
  XOR2_X1 U452 ( .A(KEYINPUT74), .B(KEYINPUT38), .Z(n343) );
  XOR2_X1 U453 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n344) );
  XOR2_X1 U454 ( .A(n611), .B(n610), .Z(n345) );
  INV_X1 U455 ( .A(n629), .ZN(n392) );
  INV_X1 U456 ( .A(n508), .ZN(n609) );
  INV_X1 U457 ( .A(n507), .ZN(n347) );
  NAND2_X1 U458 ( .A1(n351), .A2(n348), .ZN(n356) );
  INV_X1 U459 ( .A(n357), .ZN(n350) );
  NAND2_X1 U460 ( .A1(n722), .A2(n354), .ZN(n352) );
  NAND2_X1 U461 ( .A1(n357), .A2(n354), .ZN(n353) );
  NAND2_X1 U462 ( .A1(n356), .A2(n521), .ZN(n355) );
  NAND2_X1 U463 ( .A1(n508), .A2(n663), .ZN(n357) );
  XNOR2_X1 U464 ( .A(n384), .B(KEYINPUT63), .ZN(G57) );
  AND2_X1 U465 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X2 U466 ( .A(n499), .B(n498), .ZN(n722) );
  NAND2_X1 U467 ( .A1(n358), .A2(n385), .ZN(n384) );
  BUF_X1 U468 ( .A(n693), .Z(n359) );
  XNOR2_X1 U469 ( .A(n360), .B(KEYINPUT34), .ZN(n496) );
  XNOR2_X1 U470 ( .A(n406), .B(n407), .ZN(n591) );
  NOR2_X2 U471 ( .A1(n560), .A2(n468), .ZN(n361) );
  XNOR2_X2 U472 ( .A(n361), .B(KEYINPUT0), .ZN(n502) );
  XNOR2_X2 U473 ( .A(n394), .B(KEYINPUT22), .ZN(n507) );
  NAND2_X1 U474 ( .A1(n363), .A2(n362), .ZN(n520) );
  NAND2_X1 U475 ( .A1(n340), .A2(n562), .ZN(n363) );
  NAND2_X1 U476 ( .A1(n502), .A2(n517), .ZN(n365) );
  XNOR2_X2 U477 ( .A(n710), .B(G101), .ZN(n434) );
  XNOR2_X2 U478 ( .A(n490), .B(KEYINPUT4), .ZN(n710) );
  XNOR2_X2 U479 ( .A(n403), .B(n402), .ZN(n490) );
  NOR2_X1 U480 ( .A1(n359), .A2(n371), .ZN(n652) );
  NAND2_X1 U481 ( .A1(n589), .A2(n588), .ZN(n371) );
  INV_X1 U482 ( .A(n693), .ZN(n373) );
  OR2_X1 U483 ( .A1(n577), .A2(n341), .ZN(n374) );
  NAND2_X1 U484 ( .A1(n577), .A2(KEYINPUT36), .ZN(n376) );
  NAND2_X1 U485 ( .A1(n558), .A2(KEYINPUT36), .ZN(n378) );
  NAND2_X1 U486 ( .A1(n379), .A2(G469), .ZN(n595) );
  NAND2_X1 U487 ( .A1(n379), .A2(G475), .ZN(n602) );
  NAND2_X1 U488 ( .A1(n379), .A2(G210), .ZN(n682) );
  NAND2_X1 U489 ( .A1(n379), .A2(G478), .ZN(n686) );
  NAND2_X1 U490 ( .A1(n379), .A2(G217), .ZN(n690) );
  INV_X1 U491 ( .A(n410), .ZN(n618) );
  NOR2_X2 U492 ( .A1(n683), .A2(n692), .ZN(n685) );
  NOR2_X2 U493 ( .A1(n603), .A2(n692), .ZN(n605) );
  NAND2_X1 U494 ( .A1(n392), .A2(n461), .ZN(n390) );
  NAND2_X1 U495 ( .A1(n534), .A2(n461), .ZN(n391) );
  NOR2_X1 U496 ( .A1(n507), .A2(n551), .ZN(n519) );
  NAND2_X1 U497 ( .A1(n502), .A2(n501), .ZN(n394) );
  AND2_X1 U498 ( .A1(G227), .A2(n713), .ZN(n395) );
  OR2_X1 U499 ( .A1(n570), .A2(KEYINPUT47), .ZN(n396) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n549), .B(n548), .ZN(n575) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n434), .B(n452), .ZN(n406) );
  XNOR2_X1 U504 ( .A(KEYINPUT60), .B(KEYINPUT66), .ZN(n604) );
  XNOR2_X1 U505 ( .A(n418), .B(n395), .ZN(n397) );
  XNOR2_X1 U506 ( .A(G131), .B(G134), .ZN(n709) );
  XNOR2_X1 U507 ( .A(n709), .B(G146), .ZN(n435) );
  XOR2_X1 U508 ( .A(KEYINPUT78), .B(KEYINPUT93), .Z(n399) );
  XNOR2_X1 U509 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U510 ( .A(n401), .B(n400), .Z(n407) );
  XNOR2_X2 U511 ( .A(KEYINPUT64), .B(G143), .ZN(n403) );
  XNOR2_X1 U512 ( .A(n404), .B(G110), .ZN(n703) );
  XNOR2_X1 U513 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n405) );
  XNOR2_X1 U514 ( .A(n703), .B(n405), .ZN(n452) );
  XNOR2_X1 U515 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n408) );
  INV_X1 U516 ( .A(KEYINPUT1), .ZN(n409) );
  INV_X1 U517 ( .A(KEYINPUT15), .ZN(n411) );
  INV_X1 U518 ( .A(n590), .ZN(n412) );
  NAND2_X1 U519 ( .A1(n412), .A2(G234), .ZN(n413) );
  XNOR2_X1 U520 ( .A(n413), .B(KEYINPUT20), .ZN(n428) );
  NAND2_X1 U521 ( .A1(n428), .A2(G221), .ZN(n415) );
  XNOR2_X1 U522 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n414) );
  XNOR2_X1 U523 ( .A(n415), .B(n414), .ZN(n614) );
  INV_X1 U524 ( .A(KEYINPUT97), .ZN(n416) );
  XNOR2_X1 U525 ( .A(n614), .B(n416), .ZN(n500) );
  XNOR2_X1 U526 ( .A(G140), .B(KEYINPUT10), .ZN(n417) );
  XNOR2_X2 U527 ( .A(G146), .B(G125), .ZN(n447) );
  XOR2_X1 U528 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n420) );
  XNOR2_X1 U529 ( .A(G110), .B(KEYINPUT95), .ZN(n419) );
  XNOR2_X1 U530 ( .A(n420), .B(n419), .ZN(n424) );
  NAND2_X1 U531 ( .A1(G234), .A2(n713), .ZN(n425) );
  XOR2_X1 U532 ( .A(KEYINPUT8), .B(n425), .Z(n485) );
  NAND2_X1 U533 ( .A1(G221), .A2(n485), .ZN(n426) );
  XNOR2_X1 U534 ( .A(n427), .B(n426), .ZN(n689) );
  NAND2_X1 U535 ( .A1(G217), .A2(n428), .ZN(n429) );
  OR2_X2 U536 ( .A1(n500), .A2(n613), .ZN(n617) );
  XNOR2_X1 U537 ( .A(n431), .B(KEYINPUT71), .ZN(n433) );
  XNOR2_X1 U538 ( .A(n433), .B(n432), .ZN(n701) );
  XNOR2_X1 U539 ( .A(n436), .B(KEYINPUT76), .ZN(n437) );
  XOR2_X1 U540 ( .A(n435), .B(n437), .Z(n440) );
  NOR2_X1 U541 ( .A1(G953), .A2(G237), .ZN(n438) );
  XOR2_X1 U542 ( .A(KEYINPUT77), .B(n438), .Z(n476) );
  NAND2_X1 U543 ( .A1(n476), .A2(G210), .ZN(n439) );
  XNOR2_X1 U544 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U545 ( .A(n454), .B(n441), .ZN(n611) );
  XNOR2_X2 U546 ( .A(n442), .B(G472), .ZN(n624) );
  INV_X1 U547 ( .A(KEYINPUT6), .ZN(n443) );
  XNOR2_X1 U548 ( .A(n624), .B(n443), .ZN(n551) );
  NAND2_X1 U549 ( .A1(n713), .A2(G224), .ZN(n445) );
  XNOR2_X1 U550 ( .A(n445), .B(KEYINPUT79), .ZN(n449) );
  XNOR2_X1 U551 ( .A(n488), .B(KEYINPUT16), .ZN(n699) );
  XNOR2_X1 U552 ( .A(n450), .B(n699), .ZN(n451) );
  XNOR2_X1 U553 ( .A(n452), .B(n451), .ZN(n453) );
  INV_X1 U554 ( .A(G902), .ZN(n493) );
  INV_X1 U555 ( .A(G237), .ZN(n455) );
  NAND2_X1 U556 ( .A1(n493), .A2(n455), .ZN(n460) );
  NAND2_X1 U557 ( .A1(n460), .A2(G210), .ZN(n457) );
  INV_X1 U558 ( .A(KEYINPUT89), .ZN(n456) );
  NAND2_X1 U559 ( .A1(n460), .A2(G214), .ZN(n629) );
  INV_X1 U560 ( .A(KEYINPUT86), .ZN(n461) );
  NAND2_X1 U561 ( .A1(G234), .A2(G237), .ZN(n462) );
  XNOR2_X1 U562 ( .A(n462), .B(KEYINPUT14), .ZN(n464) );
  NAND2_X1 U563 ( .A1(G952), .A2(n464), .ZN(n644) );
  NOR2_X1 U564 ( .A1(G953), .A2(n644), .ZN(n528) );
  NOR2_X1 U565 ( .A1(G898), .A2(n713), .ZN(n463) );
  XOR2_X1 U566 ( .A(KEYINPUT90), .B(n463), .Z(n704) );
  NAND2_X1 U567 ( .A1(G902), .A2(n464), .ZN(n524) );
  NOR2_X1 U568 ( .A1(n704), .A2(n524), .ZN(n465) );
  XOR2_X1 U569 ( .A(KEYINPUT91), .B(n465), .Z(n466) );
  NOR2_X1 U570 ( .A1(n528), .A2(n466), .ZN(n467) );
  XNOR2_X1 U571 ( .A(n467), .B(KEYINPUT92), .ZN(n468) );
  INV_X1 U572 ( .A(n502), .ZN(n469) );
  XNOR2_X1 U573 ( .A(n471), .B(n470), .ZN(n480) );
  XOR2_X1 U574 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n473) );
  XNOR2_X1 U575 ( .A(G131), .B(KEYINPUT100), .ZN(n472) );
  XNOR2_X1 U576 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U577 ( .A(n475), .B(n474), .ZN(n478) );
  NAND2_X1 U578 ( .A1(G214), .A2(n476), .ZN(n477) );
  XNOR2_X1 U579 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U580 ( .A(n480), .B(n479), .Z(n600) );
  NOR2_X1 U581 ( .A1(G902), .A2(n600), .ZN(n482) );
  XOR2_X1 U582 ( .A(KEYINPUT13), .B(G475), .Z(n481) );
  XNOR2_X1 U583 ( .A(n482), .B(n481), .ZN(n512) );
  XOR2_X1 U584 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n484) );
  XNOR2_X1 U585 ( .A(G116), .B(KEYINPUT9), .ZN(n483) );
  XNOR2_X1 U586 ( .A(n484), .B(n483), .ZN(n487) );
  NAND2_X1 U587 ( .A1(G217), .A2(n485), .ZN(n486) );
  XNOR2_X1 U588 ( .A(n487), .B(n486), .ZN(n492) );
  XNOR2_X1 U589 ( .A(n488), .B(G134), .ZN(n489) );
  XNOR2_X1 U590 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U591 ( .A(n492), .B(n491), .ZN(n687) );
  NAND2_X1 U592 ( .A1(n687), .A2(n493), .ZN(n495) );
  INV_X1 U593 ( .A(G478), .ZN(n494) );
  XNOR2_X1 U594 ( .A(n495), .B(n494), .ZN(n510) );
  NOR2_X1 U595 ( .A1(n512), .A2(n510), .ZN(n563) );
  NAND2_X1 U596 ( .A1(n496), .A2(n563), .ZN(n499) );
  XNOR2_X1 U597 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U598 ( .A(n497), .B(KEYINPUT80), .ZN(n498) );
  NAND2_X1 U599 ( .A1(n512), .A2(n510), .ZN(n633) );
  NOR2_X1 U600 ( .A1(n633), .A2(n500), .ZN(n501) );
  INV_X1 U601 ( .A(n551), .ZN(n503) );
  AND2_X1 U602 ( .A1(n410), .A2(n613), .ZN(n504) );
  INV_X1 U603 ( .A(n624), .ZN(n542) );
  AND2_X1 U604 ( .A1(n542), .A2(n613), .ZN(n505) );
  NAND2_X1 U605 ( .A1(n618), .A2(n505), .ZN(n506) );
  INV_X1 U606 ( .A(n512), .ZN(n509) );
  NOR2_X1 U607 ( .A1(n509), .A2(n510), .ZN(n673) );
  INV_X1 U608 ( .A(n510), .ZN(n511) );
  OR2_X1 U609 ( .A1(n512), .A2(n511), .ZN(n554) );
  INV_X1 U610 ( .A(n554), .ZN(n670) );
  NOR2_X1 U611 ( .A1(n673), .A2(n670), .ZN(n513) );
  XOR2_X1 U612 ( .A(KEYINPUT102), .B(n513), .Z(n562) );
  INV_X1 U613 ( .A(n562), .ZN(n634) );
  NAND2_X1 U614 ( .A1(n624), .A2(n514), .ZN(n515) );
  NAND2_X1 U615 ( .A1(n626), .A2(n502), .ZN(n516) );
  NOR2_X1 U616 ( .A1(n523), .A2(n624), .ZN(n517) );
  NOR2_X1 U617 ( .A1(n410), .A2(n613), .ZN(n518) );
  AND2_X1 U618 ( .A1(n519), .A2(n518), .ZN(n656) );
  XNOR2_X1 U619 ( .A(n520), .B(KEYINPUT103), .ZN(n521) );
  XNOR2_X1 U620 ( .A(KEYINPUT83), .B(KEYINPUT45), .ZN(n522) );
  XOR2_X1 U621 ( .A(KEYINPUT108), .B(n523), .Z(n533) );
  OR2_X1 U622 ( .A1(n713), .A2(n524), .ZN(n525) );
  XNOR2_X1 U623 ( .A(KEYINPUT104), .B(n525), .ZN(n526) );
  NOR2_X1 U624 ( .A1(G900), .A2(n526), .ZN(n527) );
  NOR2_X1 U625 ( .A1(n528), .A2(n527), .ZN(n539) );
  XOR2_X1 U626 ( .A(KEYINPUT30), .B(KEYINPUT109), .Z(n530) );
  NAND2_X1 U627 ( .A1(n624), .A2(n629), .ZN(n529) );
  XNOR2_X1 U628 ( .A(n530), .B(n529), .ZN(n531) );
  NOR2_X1 U629 ( .A1(n539), .A2(n531), .ZN(n532) );
  NAND2_X1 U630 ( .A1(n533), .A2(n532), .ZN(n565) );
  INV_X1 U631 ( .A(n534), .ZN(n567) );
  INV_X1 U632 ( .A(n567), .ZN(n581) );
  INV_X1 U633 ( .A(n537), .ZN(n630) );
  NAND2_X1 U634 ( .A1(n630), .A2(n629), .ZN(n635) );
  NOR2_X1 U635 ( .A1(n633), .A2(n635), .ZN(n538) );
  XNOR2_X1 U636 ( .A(KEYINPUT41), .B(n538), .ZN(n646) );
  NOR2_X1 U637 ( .A1(n539), .A2(n614), .ZN(n540) );
  XNOR2_X1 U638 ( .A(KEYINPUT68), .B(n540), .ZN(n541) );
  NAND2_X1 U639 ( .A1(n541), .A2(n613), .ZN(n550) );
  NOR2_X1 U640 ( .A1(n542), .A2(n550), .ZN(n543) );
  XNOR2_X1 U641 ( .A(n543), .B(KEYINPUT28), .ZN(n546) );
  XOR2_X1 U642 ( .A(n544), .B(KEYINPUT110), .Z(n545) );
  NAND2_X1 U643 ( .A1(n546), .A2(n545), .ZN(n561) );
  NOR2_X1 U644 ( .A1(n646), .A2(n561), .ZN(n547) );
  XNOR2_X1 U645 ( .A(n547), .B(KEYINPUT42), .ZN(n725) );
  NOR2_X1 U646 ( .A1(n724), .A2(n725), .ZN(n549) );
  INV_X1 U647 ( .A(n550), .ZN(n552) );
  XNOR2_X1 U648 ( .A(n553), .B(KEYINPUT105), .ZN(n555) );
  INV_X1 U649 ( .A(n557), .ZN(n558) );
  INV_X1 U650 ( .A(n559), .ZN(n573) );
  NOR2_X1 U651 ( .A1(n561), .A2(n560), .ZN(n667) );
  NAND2_X1 U652 ( .A1(n667), .A2(n562), .ZN(n570) );
  NAND2_X1 U653 ( .A1(n570), .A2(KEYINPUT47), .ZN(n568) );
  INV_X1 U654 ( .A(n563), .ZN(n564) );
  NOR2_X1 U655 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U656 ( .A1(n567), .A2(n566), .ZN(n606) );
  NAND2_X1 U657 ( .A1(n568), .A2(n606), .ZN(n569) );
  XNOR2_X1 U658 ( .A(n569), .B(KEYINPUT81), .ZN(n571) );
  NAND2_X1 U659 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U660 ( .A(n576), .B(KEYINPUT48), .ZN(n585) );
  XOR2_X1 U661 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n580) );
  NOR2_X1 U662 ( .A1(n410), .A2(n577), .ZN(n578) );
  NAND2_X1 U663 ( .A1(n578), .A2(n629), .ZN(n579) );
  XNOR2_X1 U664 ( .A(n580), .B(n579), .ZN(n582) );
  NAND2_X1 U665 ( .A1(n582), .A2(n581), .ZN(n607) );
  NAND2_X1 U666 ( .A1(n583), .A2(n673), .ZN(n678) );
  AND2_X1 U667 ( .A1(n607), .A2(n678), .ZN(n584) );
  AND2_X2 U668 ( .A1(n585), .A2(n584), .ZN(n589) );
  XNOR2_X1 U669 ( .A(n590), .B(KEYINPUT82), .ZN(n586) );
  AND2_X1 U670 ( .A1(KEYINPUT2), .A2(n586), .ZN(n587) );
  INV_X1 U671 ( .A(KEYINPUT2), .ZN(n588) );
  XOR2_X1 U672 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n593) );
  XNOR2_X1 U673 ( .A(n591), .B(KEYINPUT120), .ZN(n592) );
  XNOR2_X1 U674 ( .A(n595), .B(n594), .ZN(n597) );
  INV_X1 U675 ( .A(G952), .ZN(n596) );
  AND2_X1 U676 ( .A1(n596), .A2(G953), .ZN(n692) );
  NOR2_X2 U677 ( .A1(n597), .A2(n692), .ZN(n599) );
  INV_X1 U678 ( .A(KEYINPUT121), .ZN(n598) );
  XNOR2_X1 U679 ( .A(n599), .B(n598), .ZN(G54) );
  XNOR2_X1 U680 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n605), .B(n604), .ZN(G60) );
  XNOR2_X1 U682 ( .A(n606), .B(n367), .ZN(G45) );
  XNOR2_X1 U683 ( .A(n607), .B(G140), .ZN(G42) );
  XOR2_X1 U684 ( .A(G119), .B(KEYINPUT126), .Z(n608) );
  XNOR2_X1 U685 ( .A(n609), .B(n608), .ZN(G21) );
  XOR2_X1 U686 ( .A(KEYINPUT87), .B(KEYINPUT62), .Z(n610) );
  AND2_X1 U687 ( .A1(n612), .A2(KEYINPUT2), .ZN(n651) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n615), .B(KEYINPUT115), .ZN(n616) );
  XNOR2_X1 U690 ( .A(KEYINPUT49), .B(n616), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n619), .B(KEYINPUT50), .ZN(n620) );
  XNOR2_X1 U693 ( .A(KEYINPUT116), .B(n620), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U696 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U697 ( .A(KEYINPUT51), .B(n627), .Z(n628) );
  NOR2_X1 U698 ( .A1(n646), .A2(n628), .ZN(n641) );
  NOR2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U700 ( .A(KEYINPUT117), .B(n631), .Z(n632) );
  NOR2_X1 U701 ( .A1(n633), .A2(n632), .ZN(n637) );
  NOR2_X1 U702 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U703 ( .A1(n637), .A2(n636), .ZN(n639) );
  NOR2_X1 U704 ( .A1(n639), .A2(n645), .ZN(n640) );
  NOR2_X1 U705 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U706 ( .A(n642), .B(KEYINPUT52), .ZN(n643) );
  NOR2_X1 U707 ( .A1(n644), .A2(n643), .ZN(n649) );
  NOR2_X1 U708 ( .A1(n646), .A2(n645), .ZN(n647) );
  OR2_X1 U709 ( .A1(G953), .A2(n647), .ZN(n648) );
  OR2_X1 U710 ( .A1(n649), .A2(n648), .ZN(n650) );
  OR2_X1 U711 ( .A1(n651), .A2(n650), .ZN(n653) );
  NOR2_X1 U712 ( .A1(n653), .A2(n652), .ZN(n655) );
  XNOR2_X1 U713 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n654) );
  XNOR2_X1 U714 ( .A(n655), .B(n654), .ZN(G75) );
  XOR2_X1 U715 ( .A(G101), .B(n656), .Z(G3) );
  XOR2_X1 U716 ( .A(G104), .B(KEYINPUT111), .Z(n658) );
  NAND2_X1 U717 ( .A1(n670), .A2(n659), .ZN(n657) );
  XNOR2_X1 U718 ( .A(n658), .B(n657), .ZN(G6) );
  XOR2_X1 U719 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n661) );
  NAND2_X1 U720 ( .A1(n673), .A2(n659), .ZN(n660) );
  XNOR2_X1 U721 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U722 ( .A(G107), .B(n662), .ZN(G9) );
  XNOR2_X1 U723 ( .A(G110), .B(n663), .ZN(G12) );
  XOR2_X1 U724 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n665) );
  NAND2_X1 U725 ( .A1(n667), .A2(n673), .ZN(n664) );
  XNOR2_X1 U726 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U727 ( .A(G128), .B(n666), .ZN(G30) );
  XOR2_X1 U728 ( .A(G146), .B(KEYINPUT113), .Z(n669) );
  NAND2_X1 U729 ( .A1(n667), .A2(n670), .ZN(n668) );
  XNOR2_X1 U730 ( .A(n669), .B(n668), .ZN(G48) );
  NAND2_X1 U731 ( .A1(n674), .A2(n670), .ZN(n671) );
  XNOR2_X1 U732 ( .A(n671), .B(KEYINPUT114), .ZN(n672) );
  XNOR2_X1 U733 ( .A(G113), .B(n672), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U735 ( .A(n675), .B(G116), .ZN(G18) );
  XOR2_X1 U736 ( .A(G125), .B(KEYINPUT37), .Z(n676) );
  XNOR2_X1 U737 ( .A(n677), .B(n676), .ZN(G27) );
  XNOR2_X1 U738 ( .A(G134), .B(n678), .ZN(G36) );
  XOR2_X1 U739 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n679) );
  XNOR2_X1 U740 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U741 ( .A(n682), .B(n681), .ZN(n683) );
  XOR2_X1 U742 ( .A(KEYINPUT56), .B(KEYINPUT119), .Z(n684) );
  XNOR2_X1 U743 ( .A(n685), .B(n684), .ZN(G51) );
  XOR2_X1 U744 ( .A(n687), .B(n686), .Z(n688) );
  NOR2_X1 U745 ( .A1(n692), .A2(n688), .ZN(G63) );
  XNOR2_X1 U746 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U747 ( .A1(n692), .A2(n691), .ZN(G66) );
  OR2_X1 U748 ( .A1(n359), .A2(G953), .ZN(n697) );
  NAND2_X1 U749 ( .A1(G953), .A2(G224), .ZN(n694) );
  XNOR2_X1 U750 ( .A(KEYINPUT61), .B(n694), .ZN(n695) );
  NAND2_X1 U751 ( .A1(n695), .A2(G898), .ZN(n696) );
  NAND2_X1 U752 ( .A1(n697), .A2(n696), .ZN(n708) );
  XNOR2_X1 U753 ( .A(G101), .B(KEYINPUT122), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n706), .B(KEYINPUT123), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n708), .B(n707), .ZN(G69) );
  XNOR2_X1 U760 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U761 ( .A(n712), .B(n711), .ZN(n716) );
  XOR2_X1 U762 ( .A(n716), .B(n589), .Z(n714) );
  NAND2_X1 U763 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n715), .B(KEYINPUT124), .ZN(n721) );
  XNOR2_X1 U765 ( .A(G227), .B(n716), .ZN(n717) );
  NAND2_X1 U766 ( .A1(n717), .A2(G900), .ZN(n718) );
  XOR2_X1 U767 ( .A(KEYINPUT125), .B(n718), .Z(n719) );
  NAND2_X1 U768 ( .A1(G953), .A2(n719), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n721), .A2(n720), .ZN(G72) );
  BUF_X1 U770 ( .A(n722), .Z(n723) );
  XOR2_X1 U771 ( .A(G122), .B(n723), .Z(G24) );
  XOR2_X1 U772 ( .A(G131), .B(n724), .Z(G33) );
  XOR2_X1 U773 ( .A(G137), .B(n725), .Z(G39) );
endmodule

