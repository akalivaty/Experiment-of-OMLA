

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735;

  XNOR2_X1 U361 ( .A(n718), .B(n394), .ZN(n621) );
  NOR2_X1 U362 ( .A1(G953), .A2(G237), .ZN(n504) );
  INV_X1 U363 ( .A(n669), .ZN(n465) );
  XOR2_X1 U364 ( .A(G104), .B(G107), .Z(n338) );
  NAND2_X2 U365 ( .A1(n387), .A2(n413), .ZN(n428) );
  XNOR2_X2 U366 ( .A(n526), .B(n525), .ZN(n573) );
  XNOR2_X2 U367 ( .A(n352), .B(n435), .ZN(n424) );
  XNOR2_X2 U368 ( .A(n723), .B(n433), .ZN(n352) );
  NAND2_X1 U369 ( .A1(n522), .A2(n554), .ZN(n397) );
  AND2_X1 U370 ( .A1(n404), .A2(n347), .ZN(n383) );
  XNOR2_X1 U371 ( .A(n545), .B(n422), .ZN(n664) );
  NOR2_X1 U372 ( .A1(n547), .A2(n680), .ZN(n545) );
  AND2_X1 U373 ( .A1(n579), .A2(n578), .ZN(n604) );
  XNOR2_X1 U374 ( .A(n412), .B(KEYINPUT41), .ZN(n703) );
  XNOR2_X1 U375 ( .A(n576), .B(n575), .ZN(n661) );
  XOR2_X1 U376 ( .A(KEYINPUT59), .B(n621), .Z(n622) );
  BUF_X1 U377 ( .A(n452), .Z(n727) );
  BUF_X1 U378 ( .A(n634), .Z(n641) );
  NAND2_X1 U379 ( .A1(n398), .A2(n341), .ZN(n366) );
  XNOR2_X1 U380 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n432) );
  NOR2_X1 U381 ( .A1(n735), .A2(n548), .ZN(n371) );
  NAND2_X1 U382 ( .A1(n420), .A2(n419), .ZN(n548) );
  NAND2_X1 U383 ( .A1(n421), .A2(n343), .ZN(n419) );
  NAND2_X1 U384 ( .A1(n664), .A2(n588), .ZN(n420) );
  NAND2_X1 U385 ( .A1(n389), .A2(n373), .ZN(n358) );
  NOR2_X1 U386 ( .A1(n633), .A2(n732), .ZN(n389) );
  XNOR2_X1 U387 ( .A(n533), .B(KEYINPUT0), .ZN(n551) );
  NOR2_X1 U388 ( .A1(n585), .A2(n532), .ZN(n533) );
  XNOR2_X1 U389 ( .A(n363), .B(n497), .ZN(n527) );
  NAND2_X1 U390 ( .A1(n350), .A2(n611), .ZN(n363) );
  OR2_X1 U391 ( .A1(n614), .A2(G902), .ZN(n483) );
  INV_X1 U392 ( .A(G953), .ZN(n452) );
  XNOR2_X1 U393 ( .A(n489), .B(n490), .ZN(n707) );
  XNOR2_X1 U394 ( .A(n606), .B(n498), .ZN(n687) );
  XNOR2_X1 U395 ( .A(G902), .B(KEYINPUT15), .ZN(n611) );
  INV_X1 U396 ( .A(KEYINPUT3), .ZN(n476) );
  XNOR2_X1 U397 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n491) );
  XNOR2_X1 U398 ( .A(n393), .B(n602), .ZN(n351) );
  XNOR2_X1 U399 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n602) );
  NAND2_X1 U400 ( .A1(n687), .A2(n686), .ZN(n692) );
  XNOR2_X1 U401 ( .A(n486), .B(n417), .ZN(n416) );
  AND2_X1 U402 ( .A1(n677), .A2(n686), .ZN(n486) );
  BUF_X1 U403 ( .A(n543), .Z(n670) );
  AND2_X1 U404 ( .A1(n351), .A2(n610), .ZN(n388) );
  XNOR2_X1 U405 ( .A(n369), .B(KEYINPUT45), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n371), .B(n379), .ZN(n370) );
  XNOR2_X1 U407 ( .A(n403), .B(n402), .ZN(n515) );
  INV_X1 U408 ( .A(KEYINPUT8), .ZN(n402) );
  NAND2_X1 U409 ( .A1(n452), .A2(G234), .ZN(n403) );
  XNOR2_X1 U410 ( .A(n492), .B(KEYINPUT10), .ZN(n503) );
  XNOR2_X1 U411 ( .A(G134), .B(G116), .ZN(n511) );
  XOR2_X1 U412 ( .A(G122), .B(G107), .Z(n512) );
  XNOR2_X1 U413 ( .A(n503), .B(n502), .ZN(n718) );
  XNOR2_X1 U414 ( .A(G143), .B(G113), .ZN(n507) );
  XOR2_X1 U415 ( .A(G131), .B(G140), .Z(n502) );
  AND2_X1 U416 ( .A1(n661), .A2(n577), .ZN(n579) );
  XNOR2_X1 U417 ( .A(n537), .B(n536), .ZN(n562) );
  XNOR2_X1 U418 ( .A(KEYINPUT22), .B(KEYINPUT65), .ZN(n536) );
  XNOR2_X1 U419 ( .A(n349), .B(n528), .ZN(n585) );
  NOR2_X1 U420 ( .A1(G902), .A2(n638), .ZN(n521) );
  NAND2_X1 U421 ( .A1(n562), .A2(n670), .ZN(n557) );
  NAND2_X1 U422 ( .A1(n704), .A2(n727), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n600), .B(KEYINPUT82), .ZN(n601) );
  INV_X1 U424 ( .A(G237), .ZN(n484) );
  INV_X1 U425 ( .A(KEYINPUT107), .ZN(n379) );
  INV_X1 U426 ( .A(KEYINPUT44), .ZN(n357) );
  INV_X1 U427 ( .A(G137), .ZN(n434) );
  NAND2_X1 U428 ( .A1(G234), .A2(G237), .ZN(n468) );
  AND2_X1 U429 ( .A1(n465), .A2(KEYINPUT108), .ZN(n406) );
  INV_X1 U430 ( .A(n687), .ZN(n355) );
  INV_X1 U431 ( .A(G902), .ZN(n485) );
  XNOR2_X1 U432 ( .A(KEYINPUT5), .B(G131), .ZN(n479) );
  XNOR2_X1 U433 ( .A(G128), .B(KEYINPUT70), .ZN(n445) );
  XNOR2_X1 U434 ( .A(KEYINPUT77), .B(G140), .ZN(n451) );
  NAND2_X1 U435 ( .A1(n385), .A2(n613), .ZN(n384) );
  NAND2_X1 U436 ( .A1(n428), .A2(n612), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n364), .B(n707), .ZN(n350) );
  XNOR2_X1 U438 ( .A(n493), .B(n494), .ZN(n418) );
  OR2_X1 U439 ( .A1(n692), .A2(n689), .ZN(n412) );
  NOR2_X1 U440 ( .A1(n416), .A2(n344), .ZN(n415) );
  BUF_X1 U441 ( .A(n527), .Z(n606) );
  INV_X1 U442 ( .A(KEYINPUT102), .ZN(n510) );
  XNOR2_X1 U443 ( .A(n392), .B(n391), .ZN(n421) );
  INV_X1 U444 ( .A(KEYINPUT99), .ZN(n391) );
  NOR2_X1 U445 ( .A1(n547), .A2(n546), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n614), .B(KEYINPUT62), .ZN(n615) );
  INV_X1 U447 ( .A(n726), .ZN(n378) );
  AND2_X1 U448 ( .A1(n348), .A2(n727), .ZN(n714) );
  XNOR2_X1 U449 ( .A(n401), .B(n516), .ZN(n517) );
  XOR2_X1 U450 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n516) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n505), .B(n507), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n508), .B(n506), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n424), .B(n430), .ZN(n642) );
  AND2_X1 U455 ( .A1(n617), .A2(G953), .ZN(n646) );
  NAND2_X1 U456 ( .A1(n399), .A2(n377), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n400), .B(n582), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n410), .B(n409), .ZN(n373) );
  INV_X1 U459 ( .A(KEYINPUT35), .ZN(n409) );
  XNOR2_X1 U460 ( .A(n544), .B(KEYINPUT100), .ZN(n422) );
  NOR2_X1 U461 ( .A1(n585), .A2(n584), .ZN(n658) );
  NOR2_X1 U462 ( .A1(n557), .A2(n541), .ZN(n542) );
  XNOR2_X1 U463 ( .A(n361), .B(n360), .ZN(G75) );
  INV_X1 U464 ( .A(KEYINPUT53), .ZN(n360) );
  NAND2_X1 U465 ( .A1(n705), .A2(n342), .ZN(n361) );
  NAND2_X1 U466 ( .A1(n674), .A2(n340), .ZN(n669) );
  AND2_X1 U467 ( .A1(n610), .A2(KEYINPUT2), .ZN(n339) );
  NOR2_X1 U468 ( .A1(n557), .A2(n556), .ZN(n633) );
  XOR2_X1 U469 ( .A(n673), .B(KEYINPUT97), .Z(n340) );
  AND2_X1 U470 ( .A1(n595), .A2(n594), .ZN(n341) );
  NOR2_X1 U471 ( .A1(n706), .A2(n362), .ZN(n342) );
  AND2_X1 U472 ( .A1(n588), .A2(n555), .ZN(n343) );
  NOR2_X1 U473 ( .A1(n565), .A2(n475), .ZN(n344) );
  AND2_X1 U474 ( .A1(n421), .A2(n555), .ZN(n345) );
  XOR2_X1 U475 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n346) );
  AND2_X1 U476 ( .A1(n612), .A2(KEYINPUT64), .ZN(n347) );
  INV_X1 U477 ( .A(KEYINPUT2), .ZN(n413) );
  NAND2_X1 U478 ( .A1(n388), .A2(n348), .ZN(n387) );
  NAND2_X1 U479 ( .A1(n429), .A2(n348), .ZN(n404) );
  OR2_X1 U480 ( .A1(n580), .A2(n349), .ZN(n400) );
  NAND2_X1 U481 ( .A1(n527), .A2(n686), .ZN(n349) );
  XNOR2_X1 U482 ( .A(n350), .B(n627), .ZN(n628) );
  AND2_X1 U483 ( .A1(n351), .A2(n339), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n352), .B(n418), .ZN(n364) );
  NAND2_X1 U485 ( .A1(n354), .A2(n353), .ZN(n501) );
  INV_X1 U486 ( .A(n390), .ZN(n353) );
  NOR2_X1 U487 ( .A1(n426), .A2(n355), .ZN(n354) );
  NOR2_X1 U488 ( .A1(n426), .A2(n390), .ZN(n356) );
  NAND2_X1 U489 ( .A1(n356), .A2(n606), .ZN(n596) );
  XNOR2_X1 U490 ( .A(n546), .B(n467), .ZN(n427) );
  NOR2_X1 U491 ( .A1(n601), .A2(n366), .ZN(n365) );
  XNOR2_X1 U492 ( .A(n358), .B(n357), .ZN(n372) );
  NOR2_X1 U493 ( .A1(n427), .A2(n475), .ZN(n426) );
  NAND2_X1 U494 ( .A1(n573), .A2(n733), .ZN(n368) );
  NAND2_X1 U495 ( .A1(n367), .A2(n365), .ZN(n393) );
  XNOR2_X1 U496 ( .A(n368), .B(n574), .ZN(n367) );
  XNOR2_X1 U497 ( .A(n448), .B(n503), .ZN(n456) );
  XNOR2_X1 U498 ( .A(n359), .B(n449), .ZN(n454) );
  XNOR2_X1 U499 ( .A(n450), .B(n451), .ZN(n359) );
  XNOR2_X2 U500 ( .A(n405), .B(n461), .ZN(n674) );
  NAND2_X1 U501 ( .A1(n372), .A2(n370), .ZN(n369) );
  XNOR2_X1 U502 ( .A(n373), .B(n731), .ZN(G24) );
  NAND2_X1 U503 ( .A1(n375), .A2(n374), .ZN(n549) );
  NAND2_X1 U504 ( .A1(n377), .A2(n406), .ZN(n374) );
  NAND2_X1 U505 ( .A1(n376), .A2(n407), .ZN(n375) );
  NAND2_X1 U506 ( .A1(n377), .A2(n465), .ZN(n376) );
  INV_X1 U507 ( .A(n543), .ZN(n377) );
  XNOR2_X1 U508 ( .A(n388), .B(n378), .ZN(n728) );
  AND2_X2 U509 ( .A1(n382), .A2(n380), .ZN(n386) );
  NAND2_X1 U510 ( .A1(n381), .A2(n613), .ZN(n380) );
  INV_X1 U511 ( .A(n404), .ZN(n381) );
  NAND2_X1 U512 ( .A1(n383), .A2(n428), .ZN(n382) );
  NAND2_X2 U513 ( .A1(n386), .A2(n384), .ZN(n634) );
  NAND2_X1 U514 ( .A1(n414), .A2(n415), .ZN(n390) );
  NOR2_X2 U515 ( .A1(n621), .A2(G902), .ZN(n509) );
  XNOR2_X2 U516 ( .A(n397), .B(KEYINPUT105), .ZN(n576) );
  INV_X1 U517 ( .A(n398), .ZN(n666) );
  NAND2_X1 U518 ( .A1(n515), .A2(G217), .ZN(n401) );
  NAND2_X1 U519 ( .A1(n702), .A2(n404), .ZN(n705) );
  INV_X1 U520 ( .A(n674), .ZN(n558) );
  NAND2_X1 U521 ( .A1(n635), .A2(n485), .ZN(n405) );
  NAND2_X1 U522 ( .A1(n377), .A2(n465), .ZN(n408) );
  OR2_X1 U523 ( .A1(n408), .A2(n555), .ZN(n680) );
  INV_X1 U524 ( .A(KEYINPUT108), .ZN(n407) );
  NAND2_X1 U525 ( .A1(n411), .A2(n597), .ZN(n410) );
  XNOR2_X1 U526 ( .A(n552), .B(n346), .ZN(n411) );
  NAND2_X1 U527 ( .A1(n427), .A2(n425), .ZN(n414) );
  INV_X1 U528 ( .A(KEYINPUT30), .ZN(n417) );
  XNOR2_X2 U529 ( .A(n423), .B(G143), .ZN(n513) );
  XNOR2_X2 U530 ( .A(G128), .B(KEYINPUT80), .ZN(n423) );
  XNOR2_X1 U531 ( .A(n424), .B(n482), .ZN(n614) );
  AND2_X1 U532 ( .A1(n565), .A2(n475), .ZN(n425) );
  INV_X1 U533 ( .A(n428), .ZN(n701) );
  XNOR2_X1 U534 ( .A(n570), .B(n538), .ZN(n543) );
  XOR2_X1 U535 ( .A(n440), .B(n439), .Z(n430) );
  XOR2_X1 U536 ( .A(KEYINPUT13), .B(G475), .Z(n431) );
  INV_X1 U537 ( .A(KEYINPUT110), .ZN(n467) );
  INV_X1 U538 ( .A(KEYINPUT84), .ZN(n581) );
  XNOR2_X1 U539 ( .A(n581), .B(KEYINPUT36), .ZN(n582) );
  XNOR2_X1 U540 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U541 ( .A(n553), .B(n510), .ZN(n522) );
  XNOR2_X2 U542 ( .A(n513), .B(n432), .ZN(n723) );
  XNOR2_X1 U543 ( .A(KEYINPUT67), .B(G101), .ZN(n433) );
  XNOR2_X1 U544 ( .A(n434), .B(G134), .ZN(n719) );
  XNOR2_X1 U545 ( .A(n719), .B(G146), .ZN(n435) );
  XNOR2_X1 U546 ( .A(G110), .B(KEYINPUT86), .ZN(n436) );
  XNOR2_X1 U547 ( .A(n338), .B(n436), .ZN(n487) );
  XOR2_X1 U548 ( .A(n487), .B(n502), .Z(n440) );
  NAND2_X1 U549 ( .A1(G227), .A2(n727), .ZN(n437) );
  XNOR2_X1 U550 ( .A(KEYINPUT90), .B(n437), .ZN(n438) );
  XNOR2_X1 U551 ( .A(n438), .B(KEYINPUT70), .ZN(n439) );
  OR2_X2 U552 ( .A1(n642), .A2(G902), .ZN(n442) );
  XNOR2_X1 U553 ( .A(KEYINPUT72), .B(G469), .ZN(n441) );
  XNOR2_X2 U554 ( .A(n442), .B(n441), .ZN(n570) );
  XNOR2_X2 U555 ( .A(G146), .B(G125), .ZN(n492) );
  XNOR2_X1 U556 ( .A(G137), .B(G119), .ZN(n444) );
  XNOR2_X1 U557 ( .A(KEYINPUT24), .B(KEYINPUT94), .ZN(n443) );
  XNOR2_X1 U558 ( .A(n444), .B(n443), .ZN(n447) );
  XNOR2_X1 U559 ( .A(n445), .B(G110), .ZN(n446) );
  XNOR2_X1 U560 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U561 ( .A(KEYINPUT23), .B(KEYINPUT93), .ZN(n450) );
  XNOR2_X1 U562 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n449) );
  NAND2_X1 U563 ( .A1(n515), .A2(G221), .ZN(n453) );
  XNOR2_X1 U564 ( .A(n456), .B(n455), .ZN(n635) );
  NAND2_X1 U565 ( .A1(n611), .A2(G234), .ZN(n458) );
  XNOR2_X1 U566 ( .A(KEYINPUT20), .B(KEYINPUT96), .ZN(n457) );
  XNOR2_X1 U567 ( .A(n458), .B(n457), .ZN(n462) );
  NAND2_X1 U568 ( .A1(n462), .A2(G217), .ZN(n460) );
  XNOR2_X1 U569 ( .A(KEYINPUT95), .B(KEYINPUT25), .ZN(n459) );
  XNOR2_X1 U570 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U571 ( .A1(n462), .A2(G221), .ZN(n464) );
  INV_X1 U572 ( .A(KEYINPUT21), .ZN(n463) );
  XNOR2_X1 U573 ( .A(n464), .B(n463), .ZN(n673) );
  NAND2_X1 U574 ( .A1(n570), .A2(n465), .ZN(n466) );
  XNOR2_X2 U575 ( .A(n466), .B(KEYINPUT98), .ZN(n546) );
  XNOR2_X1 U576 ( .A(n468), .B(KEYINPUT88), .ZN(n469) );
  XNOR2_X1 U577 ( .A(KEYINPUT14), .B(n469), .ZN(n471) );
  NAND2_X1 U578 ( .A1(n471), .A2(G952), .ZN(n470) );
  XOR2_X1 U579 ( .A(KEYINPUT89), .B(n470), .Z(n700) );
  NOR2_X1 U580 ( .A1(n700), .A2(G953), .ZN(n531) );
  INV_X1 U581 ( .A(n531), .ZN(n474) );
  AND2_X1 U582 ( .A1(n471), .A2(G953), .ZN(n472) );
  NAND2_X1 U583 ( .A1(G902), .A2(n472), .ZN(n529) );
  OR2_X1 U584 ( .A1(n529), .A2(G900), .ZN(n473) );
  NAND2_X1 U585 ( .A1(n474), .A2(n473), .ZN(n565) );
  INV_X1 U586 ( .A(KEYINPUT76), .ZN(n475) );
  XNOR2_X1 U587 ( .A(n476), .B(G119), .ZN(n478) );
  XNOR2_X1 U588 ( .A(G116), .B(G113), .ZN(n477) );
  XNOR2_X1 U589 ( .A(n478), .B(n477), .ZN(n488) );
  NAND2_X1 U590 ( .A1(n504), .A2(G210), .ZN(n480) );
  XNOR2_X1 U591 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U592 ( .A(n488), .B(n481), .ZN(n482) );
  XNOR2_X2 U593 ( .A(n483), .B(G472), .ZN(n677) );
  NAND2_X1 U594 ( .A1(n485), .A2(n484), .ZN(n495) );
  NAND2_X1 U595 ( .A1(n495), .A2(G214), .ZN(n686) );
  XOR2_X1 U596 ( .A(G122), .B(KEYINPUT16), .Z(n490) );
  XNOR2_X1 U597 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U598 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U599 ( .A1(G224), .A2(n727), .ZN(n494) );
  NAND2_X1 U600 ( .A1(G210), .A2(n495), .ZN(n496) );
  XNOR2_X1 U601 ( .A(KEYINPUT87), .B(n496), .ZN(n497) );
  INV_X1 U602 ( .A(KEYINPUT38), .ZN(n498) );
  INV_X1 U603 ( .A(KEYINPUT73), .ZN(n499) );
  XNOR2_X1 U604 ( .A(n499), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U605 ( .A(n501), .B(n500), .ZN(n523) );
  XOR2_X1 U606 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n506) );
  NAND2_X1 U607 ( .A1(G214), .A2(n504), .ZN(n505) );
  XOR2_X1 U608 ( .A(G122), .B(G104), .Z(n508) );
  XNOR2_X2 U609 ( .A(n509), .B(n431), .ZN(n553) );
  XNOR2_X1 U610 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X1 U611 ( .A(n513), .B(n514), .ZN(n518) );
  XNOR2_X1 U612 ( .A(n518), .B(n517), .ZN(n638) );
  XNOR2_X1 U613 ( .A(G478), .B(KEYINPUT103), .ZN(n519) );
  XNOR2_X1 U614 ( .A(n519), .B(KEYINPUT104), .ZN(n520) );
  XOR2_X1 U615 ( .A(n521), .B(n520), .Z(n554) );
  NOR2_X1 U616 ( .A1(n522), .A2(n554), .ZN(n663) );
  AND2_X1 U617 ( .A1(n523), .A2(n663), .ZN(n609) );
  XOR2_X1 U618 ( .A(G134), .B(n609), .Z(G36) );
  NAND2_X1 U619 ( .A1(n523), .A2(n576), .ZN(n526) );
  INV_X1 U620 ( .A(KEYINPUT113), .ZN(n524) );
  XNOR2_X1 U621 ( .A(n524), .B(KEYINPUT40), .ZN(n525) );
  XNOR2_X1 U622 ( .A(n573), .B(G131), .ZN(G33) );
  INV_X1 U623 ( .A(KEYINPUT19), .ZN(n528) );
  NOR2_X1 U624 ( .A1(G898), .A2(n529), .ZN(n530) );
  NOR2_X1 U625 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U626 ( .A1(n554), .A2(n553), .ZN(n689) );
  INV_X1 U627 ( .A(n689), .ZN(n534) );
  AND2_X1 U628 ( .A1(n340), .A2(n534), .ZN(n535) );
  NAND2_X1 U629 ( .A1(n551), .A2(n535), .ZN(n537) );
  XOR2_X1 U630 ( .A(KEYINPUT66), .B(KEYINPUT1), .Z(n538) );
  INV_X1 U631 ( .A(KEYINPUT6), .ZN(n539) );
  XNOR2_X1 U632 ( .A(n677), .B(n539), .ZN(n578) );
  INV_X1 U633 ( .A(n578), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n540), .A2(n674), .ZN(n541) );
  XNOR2_X1 U635 ( .A(n542), .B(KEYINPUT106), .ZN(n735) );
  NOR2_X1 U636 ( .A1(n576), .A2(n663), .ZN(n691) );
  INV_X1 U637 ( .A(n551), .ZN(n547) );
  XNOR2_X1 U638 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n544) );
  INV_X1 U639 ( .A(n677), .ZN(n555) );
  NAND2_X1 U640 ( .A1(n549), .A2(n578), .ZN(n550) );
  XNOR2_X2 U641 ( .A(n550), .B(KEYINPUT33), .ZN(n685) );
  NAND2_X1 U642 ( .A1(n685), .A2(n551), .ZN(n552) );
  NOR2_X1 U643 ( .A1(n554), .A2(n553), .ZN(n597) );
  NAND2_X1 U644 ( .A1(n555), .A2(n558), .ZN(n556) );
  XOR2_X1 U645 ( .A(KEYINPUT78), .B(KEYINPUT32), .Z(n564) );
  XOR2_X1 U646 ( .A(KEYINPUT79), .B(n578), .Z(n560) );
  NAND2_X1 U647 ( .A1(n377), .A2(n558), .ZN(n559) );
  NOR2_X1 U648 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U649 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U650 ( .A(n564), .B(n563), .ZN(n732) );
  NAND2_X1 U651 ( .A1(n565), .A2(n673), .ZN(n566) );
  OR2_X1 U652 ( .A1(n566), .A2(n674), .ZN(n567) );
  XNOR2_X1 U653 ( .A(n567), .B(KEYINPUT71), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n577), .A2(n677), .ZN(n569) );
  XOR2_X1 U655 ( .A(KEYINPUT28), .B(KEYINPUT112), .Z(n568) );
  XNOR2_X1 U656 ( .A(n569), .B(n568), .ZN(n571) );
  AND2_X1 U657 ( .A1(n570), .A2(n571), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n703), .A2(n583), .ZN(n572) );
  XNOR2_X1 U659 ( .A(n572), .B(KEYINPUT42), .ZN(n733) );
  INV_X1 U660 ( .A(KEYINPUT46), .ZN(n574) );
  INV_X1 U661 ( .A(KEYINPUT109), .ZN(n575) );
  XOR2_X1 U662 ( .A(KEYINPUT114), .B(n604), .Z(n580) );
  INV_X1 U663 ( .A(n583), .ZN(n584) );
  INV_X1 U664 ( .A(n658), .ZN(n587) );
  NOR2_X1 U665 ( .A1(KEYINPUT75), .A2(KEYINPUT47), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(n592) );
  XOR2_X1 U667 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n589) );
  INV_X1 U668 ( .A(n691), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n589), .A2(n588), .ZN(n593) );
  OR2_X1 U670 ( .A1(n593), .A2(KEYINPUT75), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n658), .A2(n590), .ZN(n591) );
  NAND2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n593), .A2(KEYINPUT75), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n691), .A2(KEYINPUT47), .ZN(n599) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT111), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n657) );
  NAND2_X1 U677 ( .A1(n599), .A2(n657), .ZN(n600) );
  AND2_X1 U678 ( .A1(n670), .A2(n686), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n605), .B(KEYINPUT43), .ZN(n608) );
  INV_X1 U681 ( .A(n606), .ZN(n607) );
  AND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n668) );
  NOR2_X1 U683 ( .A1(n609), .A2(n668), .ZN(n610) );
  INV_X1 U684 ( .A(n611), .ZN(n612) );
  INV_X1 U685 ( .A(KEYINPUT64), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n634), .A2(G472), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n616), .B(n615), .ZN(n618) );
  INV_X1 U688 ( .A(G952), .ZN(n617) );
  NOR2_X2 U689 ( .A1(n618), .A2(n646), .ZN(n620) );
  INV_X1 U690 ( .A(KEYINPUT63), .ZN(n619) );
  XNOR2_X1 U691 ( .A(n620), .B(n619), .ZN(G57) );
  NAND2_X1 U692 ( .A1(n634), .A2(G475), .ZN(n623) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X2 U694 ( .A1(n624), .A2(n646), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U696 ( .A1(n634), .A2(G210), .ZN(n629) );
  XNOR2_X1 U697 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n626) );
  XOR2_X1 U698 ( .A(n626), .B(KEYINPUT55), .Z(n627) );
  XNOR2_X1 U699 ( .A(n629), .B(n628), .ZN(n630) );
  NOR2_X2 U700 ( .A1(n630), .A2(n646), .ZN(n632) );
  XNOR2_X1 U701 ( .A(KEYINPUT122), .B(KEYINPUT56), .ZN(n631) );
  XNOR2_X1 U702 ( .A(n632), .B(n631), .ZN(G51) );
  XOR2_X1 U703 ( .A(G110), .B(n633), .Z(G12) );
  AND2_X1 U704 ( .A1(n641), .A2(G217), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(n637) );
  NOR2_X1 U706 ( .A1(n637), .A2(n646), .ZN(G66) );
  NAND2_X1 U707 ( .A1(n641), .A2(G478), .ZN(n639) );
  XNOR2_X1 U708 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X1 U709 ( .A1(n640), .A2(n646), .ZN(G63) );
  NAND2_X1 U710 ( .A1(n641), .A2(G469), .ZN(n645) );
  XOR2_X1 U711 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n643) );
  XNOR2_X1 U712 ( .A(n642), .B(n643), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n645), .B(n644), .ZN(n647) );
  NOR2_X1 U714 ( .A1(n647), .A2(n646), .ZN(G54) );
  NAND2_X1 U715 ( .A1(n345), .A2(n661), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n648), .B(G104), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT115), .B(KEYINPUT26), .Z(n650) );
  NAND2_X1 U718 ( .A1(n345), .A2(n663), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(n652) );
  XOR2_X1 U720 ( .A(G107), .B(KEYINPUT27), .Z(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(G9) );
  AND2_X1 U722 ( .A1(n658), .A2(n663), .ZN(n656) );
  XOR2_X1 U723 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n654) );
  XNOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n656), .B(n655), .ZN(G30) );
  XNOR2_X1 U727 ( .A(G143), .B(n657), .ZN(G45) );
  NAND2_X1 U728 ( .A1(n658), .A2(n661), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n659), .B(KEYINPUT118), .ZN(n660) );
  XNOR2_X1 U730 ( .A(G146), .B(n660), .ZN(G48) );
  NAND2_X1 U731 ( .A1(n664), .A2(n661), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n662), .B(G113), .ZN(G15) );
  NAND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n665), .B(G116), .ZN(G18) );
  XNOR2_X1 U735 ( .A(G125), .B(n666), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n667), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U737 ( .A(G140), .B(n668), .Z(G42) );
  NAND2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n672) );
  XOR2_X1 U739 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n671) );
  XNOR2_X1 U740 ( .A(n672), .B(n671), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U742 ( .A(KEYINPUT49), .B(n675), .Z(n676) );
  NOR2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n683) );
  XOR2_X1 U746 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n682) );
  XNOR2_X1 U747 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n703), .A2(n684), .ZN(n697) );
  NOR2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U751 ( .A(n690), .B(KEYINPUT121), .ZN(n694) );
  OR2_X1 U752 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U753 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U754 ( .A1(n685), .A2(n695), .ZN(n696) );
  NAND2_X1 U755 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U756 ( .A(KEYINPUT52), .B(n698), .Z(n699) );
  NOR2_X1 U757 ( .A1(n700), .A2(n699), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n701), .B(KEYINPUT81), .ZN(n702) );
  NAND2_X1 U759 ( .A1(n703), .A2(n685), .ZN(n704) );
  XOR2_X1 U760 ( .A(G101), .B(n707), .Z(n709) );
  NOR2_X1 U761 ( .A1(G898), .A2(n727), .ZN(n708) );
  NOR2_X1 U762 ( .A1(n709), .A2(n708), .ZN(n717) );
  INV_X1 U763 ( .A(G898), .ZN(n713) );
  NAND2_X1 U764 ( .A1(G224), .A2(G953), .ZN(n710) );
  XNOR2_X1 U765 ( .A(n710), .B(KEYINPUT123), .ZN(n711) );
  XNOR2_X1 U766 ( .A(n711), .B(KEYINPUT61), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n713), .A2(n712), .ZN(n715) );
  NOR2_X1 U768 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U769 ( .A(n717), .B(n716), .Z(G69) );
  XNOR2_X1 U770 ( .A(n718), .B(KEYINPUT124), .ZN(n721) );
  XNOR2_X1 U771 ( .A(n719), .B(KEYINPUT70), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U773 ( .A(n723), .B(n722), .ZN(n726) );
  XNOR2_X1 U774 ( .A(n726), .B(G227), .ZN(n724) );
  NAND2_X1 U775 ( .A1(G900), .A2(n724), .ZN(n725) );
  NAND2_X1 U776 ( .A1(n725), .A2(G953), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U778 ( .A1(n730), .A2(n729), .ZN(G72) );
  XOR2_X1 U779 ( .A(G122), .B(KEYINPUT125), .Z(n731) );
  XOR2_X1 U780 ( .A(G119), .B(n732), .Z(G21) );
  XNOR2_X1 U781 ( .A(G137), .B(n733), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(KEYINPUT126), .ZN(G39) );
  XOR2_X1 U783 ( .A(n735), .B(G101), .Z(G3) );
endmodule

