//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(G2104), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR3_X1   g037(.A1(new_n462), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n463));
  OAI21_X1  g038(.A(G101), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(KEYINPUT65), .A3(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n460), .A4(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n470), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n472), .B1(G2105), .B2(new_n476), .ZN(G160));
  INV_X1    g052(.A(new_n471), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n469), .A2(new_n470), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(G2105), .A3(new_n468), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n460), .B2(G112), .ZN(new_n484));
  OAI221_X1 g059(.A(new_n479), .B1(new_n481), .B2(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  AND2_X1   g061(.A1(KEYINPUT4), .A2(G138), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(G102), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n468), .A2(new_n469), .A3(G126), .A4(new_n470), .ZN(new_n491));
  NAND2_X1  g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n460), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n460), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT4), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n490), .A2(new_n493), .A3(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G62), .ZN(new_n500));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(KEYINPUT67), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n499), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n502), .A2(KEYINPUT67), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  INV_X1    g090(.A(G89), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n505), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n499), .A2(G63), .A3(G651), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n507), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n517), .A2(new_n520), .ZN(G168));
  INV_X1    g096(.A(G90), .ZN(new_n522));
  INV_X1    g097(.A(G52), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n505), .A2(new_n522), .B1(new_n507), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT68), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(new_n498), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(G171));
  INV_X1    g103(.A(G81), .ZN(new_n529));
  INV_X1    g104(.A(G43), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n505), .A2(new_n529), .B1(new_n507), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n498), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(KEYINPUT69), .B1(new_n531), .B2(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  NAND4_X1  g115(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT70), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  AND2_X1   g120(.A1(KEYINPUT71), .A2(G53), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n504), .A2(G543), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT9), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n499), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n548), .A2(new_n549), .B1(G651), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n505), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n499), .A2(new_n504), .A3(KEYINPUT72), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(G91), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G299));
  NAND2_X1  g134(.A1(new_n525), .A2(new_n527), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  OR2_X1    g136(.A1(new_n499), .A2(G74), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n504), .A2(G543), .ZN(new_n563));
  AOI22_X1  g138(.A1(G651), .A2(new_n562), .B1(new_n563), .B2(G49), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n556), .A2(G87), .A3(new_n557), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT73), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n568), .A2(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n551), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(new_n563), .B2(G48), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n556), .A2(new_n557), .ZN(new_n576));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(G305));
  XOR2_X1   g153(.A(KEYINPUT74), .B(G85), .Z(new_n579));
  INV_X1    g154(.A(G47), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n505), .A2(new_n579), .B1(new_n507), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G72), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G60), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n551), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n581), .B1(G651), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n556), .A2(G92), .A3(new_n557), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n563), .A2(KEYINPUT76), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n593), .B1(new_n507), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n551), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n592), .A2(new_n595), .B1(new_n598), .B2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n591), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n589), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n589), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  XNOR2_X1  g181(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND3_X1  g184(.A1(new_n601), .A2(new_n608), .A3(G868), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n539), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT11), .Z(G282));
  INV_X1    g189(.A(new_n613), .ZN(G323));
  OR2_X1    g190(.A1(new_n461), .A2(new_n463), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n494), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n478), .A2(G135), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n625));
  OAI221_X1 g200(.A(new_n622), .B1(new_n481), .B2(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n621), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT79), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT81), .ZN(new_n645));
  INV_X1    g220(.A(G14), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n643), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(KEYINPUT80), .A3(new_n643), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n645), .A2(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT82), .ZN(new_n654));
  NOR2_X1   g229(.A1(G2072), .A2(G2078), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n442), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2084), .B(G2090), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n656), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(KEYINPUT17), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n660), .B(new_n657), .C1(new_n654), .C2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n657), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n654), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n627), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(G2096), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(new_n620), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT83), .ZN(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n676), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n677), .A2(KEYINPUT20), .A3(new_n676), .ZN(new_n682));
  OAI221_X1 g257(.A(new_n678), .B1(new_n676), .B2(new_n674), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  INV_X1    g262(.A(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n689), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(G229));
  OR2_X1    g267(.A1(G16), .A2(G22), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(G303), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1971), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n694), .A2(G6), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G305), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n569), .A2(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n694), .A2(G23), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(KEYINPUT33), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n701), .A2(new_n705), .A3(new_n702), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n704), .A2(G1976), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G1976), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n696), .A2(new_n700), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n713), .A2(new_n714), .A3(KEYINPUT34), .ZN(new_n715));
  MUX2_X1   g290(.A(G24), .B(G290), .S(G16), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1986), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  OR2_X1    g294(.A1(G95), .A2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n720), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n721));
  INV_X1    g296(.A(G131), .ZN(new_n722));
  INV_X1    g297(.A(G119), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n721), .B1(new_n722), .B2(new_n471), .C1(new_n481), .C2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n719), .B1(new_n728), .B2(G29), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT35), .B(G1991), .Z(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n731), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n732), .A2(KEYINPUT85), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(KEYINPUT85), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n717), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n715), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(KEYINPUT34), .B1(new_n713), .B2(new_n714), .ZN(new_n738));
  OAI21_X1  g313(.A(KEYINPUT36), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n713), .A2(new_n714), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT34), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n742), .A2(new_n743), .A3(new_n715), .A4(new_n736), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n694), .A2(G4), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n601), .B2(new_n694), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT87), .B(G1348), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n718), .B1(KEYINPUT24), .B2(G34), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(KEYINPUT24), .B2(G34), .ZN(new_n751));
  INV_X1    g326(.A(G160), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(G29), .ZN(new_n753));
  INV_X1    g328(.A(G2084), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT91), .ZN(new_n756));
  INV_X1    g331(.A(G2090), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n718), .A2(G35), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n718), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT29), .Z(new_n760));
  AOI21_X1  g335(.A(new_n756), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n749), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n694), .A2(G20), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT23), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1956), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n760), .B2(new_n757), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n694), .A2(G19), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n539), .B2(new_n694), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT88), .B(G1341), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n718), .A2(G33), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT90), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT25), .Z(new_n777));
  AOI22_X1  g352(.A1(new_n494), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n778));
  INV_X1    g353(.A(G139), .ZN(new_n779));
  OAI22_X1  g354(.A1(new_n778), .A2(new_n460), .B1(new_n779), .B2(new_n471), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n774), .B1(new_n781), .B2(new_n718), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G2072), .Z(new_n783));
  NOR2_X1   g358(.A1(G164), .A2(new_n718), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G27), .B2(new_n718), .ZN(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n718), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  OAI21_X1  g364(.A(KEYINPUT89), .B1(G104), .B2(G2105), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(KEYINPUT89), .A2(G104), .A3(G2105), .ZN(new_n792));
  OAI221_X1 g367(.A(G2104), .B1(G116), .B2(new_n460), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G128), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n481), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G140), .B2(new_n478), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n789), .B1(new_n796), .B2(new_n718), .ZN(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n773), .A2(new_n783), .A3(new_n787), .A4(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G28), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT30), .ZN(new_n802));
  AOI21_X1  g377(.A(G29), .B1(new_n801), .B2(KEYINPUT30), .ZN(new_n803));
  OR2_X1    g378(.A1(KEYINPUT31), .A2(G11), .ZN(new_n804));
  NAND2_X1  g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G168), .A2(new_n694), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n694), .B2(G21), .ZN(new_n808));
  INV_X1    g383(.A(G1966), .ZN(new_n809));
  OAI221_X1 g384(.A(new_n806), .B1(new_n718), .B2(new_n626), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n694), .A2(G5), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G171), .B2(new_n694), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n810), .B1(G1961), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n786), .B2(new_n785), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n808), .A2(new_n809), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n753), .A2(new_n754), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n816), .B(new_n817), .C1(G1961), .C2(new_n812), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n800), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT26), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n616), .A2(G105), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n478), .A2(G141), .ZN(new_n825));
  INV_X1    g400(.A(G129), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n481), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(new_n718), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT92), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(KEYINPUT92), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n829), .A2(new_n830), .B1(G29), .B2(G32), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT27), .B(G1996), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n769), .A2(new_n819), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT95), .B1(new_n745), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n838));
  AOI211_X1 g413(.A(new_n838), .B(new_n835), .C1(new_n739), .C2(new_n744), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(G311));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n745), .B2(new_n836), .ZN(new_n842));
  AOI211_X1 g417(.A(KEYINPUT96), .B(new_n835), .C1(new_n739), .C2(new_n744), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(G150));
  XOR2_X1   g419(.A(KEYINPUT97), .B(G93), .Z(new_n845));
  INV_X1    g420(.A(G55), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n505), .A2(new_n845), .B1(new_n507), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT98), .Z(new_n848));
  AOI22_X1  g423(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(new_n498), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n538), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n848), .A2(new_n534), .A3(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n601), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n851), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(G145));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n728), .A2(KEYINPUT100), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n728), .A2(KEYINPUT100), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n618), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(new_n618), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n866), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(G106), .A2(G2105), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(new_n460), .B2(G118), .ZN(new_n876));
  OAI22_X1  g451(.A1(new_n481), .A2(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(G142), .B2(new_n478), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n869), .A2(new_n872), .A3(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n796), .B(G164), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n883), .A2(new_n827), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n827), .ZN(new_n885));
  INV_X1    g460(.A(new_n781), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n886), .B1(new_n884), .B2(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n865), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n881), .A3(new_n880), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n626), .B(G160), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(G162), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n892), .A2(new_n865), .A3(new_n881), .A4(new_n880), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n882), .B2(new_n890), .ZN(new_n899));
  AOI21_X1  g474(.A(G37), .B1(new_n899), .B2(new_n893), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g477(.A1(new_n601), .A2(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n600), .A2(new_n605), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT41), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n601), .A2(new_n608), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n854), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n904), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n910), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G303), .B(G305), .ZN(new_n916));
  NAND2_X1  g491(.A1(G290), .A2(new_n569), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n586), .A2(new_n566), .A3(new_n587), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n919), .B2(KEYINPUT102), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(KEYINPUT102), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n913), .B2(KEYINPUT42), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n914), .B1(new_n910), .B2(new_n912), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n915), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n915), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n851), .A2(new_n611), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(G295));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n928), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  NAND2_X1  g506(.A1(G286), .A2(KEYINPUT104), .ZN(new_n932));
  OR2_X1    g507(.A1(G286), .A2(KEYINPUT104), .ZN(new_n933));
  NAND3_X1  g508(.A1(G171), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(G301), .A2(KEYINPUT104), .A3(G286), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n936), .A2(new_n854), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n854), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n906), .B2(new_n905), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n911), .A3(new_n938), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n922), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n922), .A2(new_n940), .A3(new_n941), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n931), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n944), .A2(new_n946), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n947), .A3(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(G397));
  NAND2_X1  g529(.A1(new_n491), .A2(new_n492), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n496), .B1(new_n955), .B2(G2105), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n488), .A2(new_n489), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n460), .ZN(new_n958));
  AOI21_X1  g533(.A(G1384), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT105), .B(G40), .Z(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n475), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n494), .B2(G125), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n964), .B2(new_n460), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT106), .B1(new_n965), .B2(new_n472), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n961), .B1(new_n476), .B2(G2105), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n480), .A2(G137), .A3(new_n460), .A4(new_n468), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n464), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n960), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(G290), .A2(G1986), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n974), .A2(KEYINPUT107), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(KEYINPUT107), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT108), .Z(new_n979));
  OAI21_X1  g554(.A(new_n973), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n796), .B(new_n798), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n973), .A2(new_n981), .A3(KEYINPUT109), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n827), .B(G1996), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n984), .A2(new_n985), .B1(new_n973), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n728), .A2(new_n731), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n730), .B1(new_n726), .B2(new_n727), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n973), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n980), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n955), .A2(G2105), .ZN(new_n994));
  INV_X1    g569(.A(new_n496), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n958), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n971), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n809), .B1(new_n1000), .B2(new_n960), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n996), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT114), .B(G2084), .Z(new_n1006));
  NAND4_X1  g581(.A1(new_n1002), .A2(new_n971), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1001), .A2(KEYINPUT120), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT120), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g584(.A(G168), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n993), .B1(new_n1010), .B2(G8), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1007), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n970), .A2(new_n966), .B1(new_n996), .B2(new_n998), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n997), .B1(G164), .B2(G1384), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1966), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1012), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1001), .A2(KEYINPUT120), .A3(new_n1007), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  NOR2_X1   g594(.A1(G168), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1001), .A2(new_n1007), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n993), .B(G8), .C1(new_n1022), .C2(G286), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT62), .B1(new_n1011), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT110), .B1(new_n959), .B2(KEYINPUT45), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1027), .B(new_n997), .C1(G164), .C2(G1384), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1014), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1971), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1002), .A2(new_n757), .A3(new_n1005), .A4(new_n971), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT111), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1019), .B1(new_n510), .B2(new_n511), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1035), .A2(KEYINPUT55), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT112), .B1(new_n1035), .B2(KEYINPUT55), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1031), .A2(new_n1043), .A3(new_n1032), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1034), .A2(G8), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1042), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1033), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n1019), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT113), .B(G1976), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n568), .A2(new_n570), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1019), .B1(new_n971), .B2(new_n959), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n709), .B2(new_n569), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n575), .B1(new_n577), .B2(new_n505), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G1981), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT49), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n575), .B(new_n688), .C1(new_n577), .C2(new_n576), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1053), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1054), .A2(KEYINPUT52), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1055), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1045), .A2(new_n1048), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G286), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT51), .B1(new_n1066), .B2(new_n1019), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1029), .B2(G2078), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1014), .A2(KEYINPUT53), .A3(new_n786), .A4(new_n1015), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT121), .B(new_n1071), .C1(new_n1029), .C2(G2078), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1002), .A2(new_n971), .A3(new_n1005), .ZN(new_n1077));
  INV_X1    g652(.A(G1961), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G171), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1025), .A2(new_n1065), .A3(new_n1070), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1081), .B1(new_n1086), .B2(KEYINPUT62), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1087), .A2(KEYINPUT123), .A3(new_n1065), .A4(new_n1070), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  NOR4_X1   g664(.A1(new_n1060), .A2(G288), .A3(new_n1061), .A4(G1976), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1059), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1053), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1064), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(new_n1045), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT63), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1045), .A2(new_n1048), .A3(new_n1064), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1022), .A2(G8), .A3(G168), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1034), .A2(G8), .A3(new_n1044), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n1046), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1097), .A2(new_n1095), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1100), .A2(new_n1045), .A3(new_n1064), .A4(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1094), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n554), .A2(new_n558), .A3(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1077), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1026), .A2(new_n1014), .A3(new_n1028), .A4(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1110), .A2(new_n1112), .A3(KEYINPUT117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1108), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1348), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1077), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n971), .A2(new_n959), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n798), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1127));
  OR3_X1    g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n600), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1114), .B1(new_n1120), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1108), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1114), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT58), .B(G1341), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n1029), .A2(G1996), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n538), .B1(KEYINPUT118), .B2(KEYINPUT59), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1134), .B(new_n1135), .C1(KEYINPUT118), .C2(KEYINPUT59), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1132), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT60), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n601), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT60), .B(new_n600), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OR3_X1    g719(.A1(new_n1126), .A2(new_n1127), .A3(KEYINPUT60), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1113), .A2(KEYINPUT61), .ZN(new_n1148));
  OR3_X1    g723(.A1(new_n1119), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1119), .B2(new_n1148), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1129), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1072), .A2(new_n1073), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n1154));
  INV_X1    g729(.A(G40), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n752), .B2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1071), .B(G2078), .C1(new_n996), .C2(new_n998), .ZN(new_n1157));
  NAND3_X1  g732(.A1(G160), .A2(KEYINPUT122), .A3(G40), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1015), .A4(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1153), .A2(G301), .A3(new_n1076), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1081), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1153), .A2(G301), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1153), .A2(new_n1076), .A3(new_n1159), .ZN(new_n1165));
  OAI211_X1 g740(.A(KEYINPUT54), .B(new_n1164), .C1(new_n1165), .C2(G301), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1163), .A2(new_n1166), .A3(new_n1065), .A4(new_n1086), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1103), .B1(new_n1152), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n992), .B1(new_n1089), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n973), .B1(new_n981), .B2(new_n827), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT46), .ZN(new_n1171));
  OR3_X1    g746(.A1(new_n972), .A2(new_n1171), .A3(G1996), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1171), .B1(new_n972), .B2(G1996), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1175));
  XNOR2_X1  g750(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n975), .A2(new_n973), .A3(new_n976), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT48), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1176), .B1(new_n1178), .B2(new_n991), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n987), .A2(new_n988), .B1(new_n798), .B2(new_n796), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT124), .B1(new_n1180), .B2(new_n972), .ZN(new_n1181));
  OR3_X1    g756(.A1(new_n1180), .A2(KEYINPUT124), .A3(new_n972), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1169), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g761(.A1(new_n952), .A2(new_n947), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n667), .A2(new_n669), .A3(G319), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1190));
  OR2_X1    g764(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n1191), .B(new_n1192), .C1(new_n690), .C2(new_n691), .ZN(new_n1193));
  AOI21_X1  g767(.A(new_n1193), .B1(new_n645), .B2(new_n651), .ZN(new_n1194));
  AND3_X1   g768(.A1(new_n1188), .A2(new_n1194), .A3(new_n901), .ZN(G308));
  NAND3_X1  g769(.A1(new_n1188), .A2(new_n1194), .A3(new_n901), .ZN(G225));
endmodule


