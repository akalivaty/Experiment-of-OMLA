//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n209), .B(new_n215), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n228), .B(new_n231), .Z(G358));
  XOR2_X1   g0032(.A(G58), .B(G77), .Z(new_n233));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  INV_X1    g0039(.A(G1), .ZN(new_n240));
  NAND3_X1  g0040(.A1(new_n240), .A2(G13), .A3(G20), .ZN(new_n241));
  NAND3_X1  g0041(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(new_n212), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n244), .B1(G1), .B2(new_n213), .ZN(new_n245));
  MUX2_X1   g0045(.A(new_n241), .B(new_n245), .S(G50), .Z(new_n246));
  INV_X1    g0046(.A(G150), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  OAI22_X1  g0049(.A1(new_n247), .A2(new_n249), .B1(new_n201), .B2(new_n213), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT8), .ZN(new_n251));
  INV_X1    g0051(.A(G58), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT67), .ZN(new_n253));
  OAI21_X1  g0053(.A(KEYINPUT67), .B1(new_n252), .B2(KEYINPUT68), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n253), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(new_n251), .B2(new_n254), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n250), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n246), .B1(new_n259), .B2(new_n244), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT9), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G222), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n265), .B1(new_n202), .B2(new_n263), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n212), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(KEYINPUT66), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT66), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G33), .A3(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(new_n269), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(G274), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n280), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G226), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n273), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G190), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT71), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT10), .B1(new_n285), .B2(G200), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n262), .A2(new_n288), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(G200), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(new_n261), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n277), .A2(G238), .A3(new_n282), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n281), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n263), .A2(G232), .A3(G1698), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G97), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT3), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G33), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n300), .A2(new_n302), .A3(G226), .A4(new_n264), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n298), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n272), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n297), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n297), .B2(new_n305), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G190), .ZN(new_n310));
  INV_X1    g0110(.A(G68), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n248), .A2(G50), .B1(G20), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n258), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n202), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n314), .A2(new_n243), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n315), .A2(KEYINPUT11), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(KEYINPUT11), .ZN(new_n317));
  OR3_X1    g0117(.A1(new_n241), .A2(KEYINPUT12), .A3(G68), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT12), .B1(new_n241), .B2(G68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n311), .B2(new_n245), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(G200), .B1(new_n307), .B2(new_n308), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n310), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n297), .A2(new_n305), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT13), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n297), .A2(new_n305), .A3(new_n306), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT14), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT72), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n333), .B(KEYINPUT14), .C1(new_n309), .C2(new_n326), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n309), .A2(G179), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n331), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n332), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n322), .B(KEYINPUT73), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n325), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n285), .A2(G179), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n285), .A2(new_n326), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n260), .A3(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT8), .B(G58), .Z(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT15), .B(G87), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n313), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n243), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT69), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n263), .A2(G232), .A3(new_n264), .ZN(new_n350));
  INV_X1    g0150(.A(G107), .ZN(new_n351));
  INV_X1    g0151(.A(G238), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n350), .B1(new_n351), .B2(new_n263), .C1(new_n266), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n272), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n283), .A2(G244), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n354), .A2(G190), .A3(new_n281), .A4(new_n355), .ZN(new_n356));
  MUX2_X1   g0156(.A(new_n241), .B(new_n245), .S(G77), .Z(new_n357));
  AND3_X1   g0157(.A1(new_n349), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(new_n281), .A3(new_n355), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G200), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n349), .A2(new_n357), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n359), .A2(G179), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n326), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n295), .A2(new_n339), .A3(new_n342), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n256), .A2(new_n245), .ZN(new_n368));
  INV_X1    g0168(.A(new_n241), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n256), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n300), .A2(new_n302), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT7), .B1(new_n371), .B2(new_n213), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  AOI211_X1 g0173(.A(new_n373), .B(G20), .C1(new_n300), .C2(new_n302), .ZN(new_n374));
  OAI21_X1  g0174(.A(G68), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n252), .A2(new_n311), .ZN(new_n376));
  NOR2_X1   g0176(.A1(G58), .A2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n248), .A2(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT16), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n373), .B1(new_n263), .B2(G20), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n371), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n311), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(KEYINPUT16), .A3(new_n379), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n243), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT74), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n382), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n386), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n244), .B1(new_n375), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n385), .B2(new_n380), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT74), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n370), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n277), .A2(G232), .A3(new_n282), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n281), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n300), .A2(new_n302), .A3(G226), .A4(G1698), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n300), .A2(new_n302), .A3(G223), .A4(new_n264), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT75), .A4(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n401), .A2(new_n272), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n397), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G179), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n272), .A3(new_n401), .ZN(new_n408));
  INV_X1    g0208(.A(new_n397), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G169), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n395), .A2(new_n412), .A3(KEYINPUT18), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT76), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n388), .B1(new_n382), .B2(new_n387), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n391), .A2(KEYINPUT74), .A3(new_n393), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n370), .B1(new_n411), .B2(new_n407), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(KEYINPUT76), .A3(KEYINPUT18), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n395), .A2(new_n412), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n415), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n256), .A2(new_n369), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n256), .B2(new_n245), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n416), .B2(new_n417), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n408), .A2(new_n286), .A3(new_n409), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n406), .B2(G200), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n427), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT17), .B1(new_n427), .B2(new_n429), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n424), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n240), .A2(G45), .ZN(new_n434));
  OR2_X1    g0234(.A1(KEYINPUT5), .A2(G41), .ZN(new_n435));
  NAND2_X1  g0235(.A1(KEYINPUT5), .A2(G41), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n277), .A3(G274), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n279), .A2(G1), .ZN(new_n439));
  AND2_X1   g0239(.A1(KEYINPUT5), .A2(G41), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n277), .A2(new_n442), .A3(G264), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n300), .A2(new_n302), .A3(G257), .A4(G1698), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n300), .A2(new_n302), .A3(G250), .A4(new_n264), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G294), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT84), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n272), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n448), .B2(new_n272), .ZN(new_n452));
  OAI21_X1  g0252(.A(G169), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n277), .A2(new_n442), .ZN(new_n454));
  AOI22_X1  g0254(.A1(G264), .A2(new_n454), .B1(new_n448), .B2(new_n272), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(G179), .A3(new_n438), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n300), .A2(new_n302), .A3(new_n213), .A4(G87), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT22), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n263), .A2(new_n460), .A3(new_n213), .A4(G87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G116), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT23), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n213), .B2(G107), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n351), .A2(KEYINPUT23), .A3(G20), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n462), .A2(new_n463), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n463), .B1(new_n462), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n243), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XOR2_X1   g0272(.A(KEYINPUT83), .B(KEYINPUT25), .Z(new_n473));
  NOR2_X1   g0273(.A1(new_n241), .A2(G107), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n240), .A2(G33), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n244), .A2(new_n241), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(G107), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n457), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n448), .A2(new_n272), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT84), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(new_n286), .A3(new_n450), .A4(new_n444), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n438), .A3(new_n443), .ZN(new_n485));
  INV_X1    g0285(.A(G200), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n472), .A3(new_n479), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n263), .A2(new_n213), .A3(G68), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n263), .A2(KEYINPUT81), .A3(new_n213), .A4(G68), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT19), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n258), .A2(new_n494), .A3(G97), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  INV_X1    g0296(.A(G87), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n496), .A2(new_n497), .B1(new_n299), .B2(new_n213), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(new_n494), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n492), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n243), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n345), .A2(new_n369), .ZN(new_n502));
  OR2_X1    g0302(.A1(new_n477), .A2(new_n497), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n434), .A2(G274), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n505), .B(new_n277), .C1(G250), .C2(new_n439), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n300), .A2(new_n302), .A3(G244), .A4(G1698), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n464), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT80), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n263), .A2(new_n509), .A3(G238), .A4(new_n264), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n300), .A2(new_n302), .A3(G238), .A4(new_n264), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT80), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G190), .B(new_n506), .C1(new_n513), .C2(new_n271), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n506), .B1(new_n513), .B2(new_n271), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G200), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n504), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n501), .B(new_n502), .C1(new_n345), .C2(new_n477), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n326), .ZN(new_n519));
  INV_X1    g0319(.A(G179), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n506), .C1(new_n513), .C2(new_n271), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n481), .A2(new_n489), .A3(new_n517), .A4(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT82), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n277), .A2(new_n442), .A3(G270), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n438), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n300), .A2(new_n302), .A3(G264), .A4(G1698), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n300), .A2(new_n302), .A3(G257), .A4(new_n264), .ZN(new_n528));
  INV_X1    g0328(.A(G303), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n263), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n272), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(G190), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G116), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n369), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n244), .A2(G116), .A3(new_n241), .A4(new_n476), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n242), .A2(new_n212), .B1(G20), .B2(new_n533), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  INV_X1    g0337(.A(G97), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n213), .C1(G33), .C2(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT20), .B1(new_n536), .B2(new_n539), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n534), .B(new_n535), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n532), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n486), .B1(new_n526), .B2(new_n531), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n524), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n526), .A2(new_n531), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(KEYINPUT82), .A3(new_n543), .A4(new_n532), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n547), .A2(KEYINPUT21), .A3(G169), .A4(new_n542), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n542), .A2(new_n526), .A3(G179), .A4(new_n531), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n326), .B1(new_n526), .B2(new_n531), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT21), .B1(new_n554), .B2(new_n542), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n523), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n300), .A2(new_n302), .A3(G244), .A4(new_n264), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT4), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n264), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n537), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n272), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n277), .A2(new_n442), .A3(G257), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n438), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n326), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n564), .A2(KEYINPUT78), .A3(new_n272), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT78), .B1(new_n564), .B2(new_n272), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n520), .B(new_n568), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  XNOR2_X1  g0373(.A(G97), .B(G107), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT6), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n575), .A2(new_n538), .A3(G107), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n213), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n249), .A2(new_n202), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT77), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT77), .ZN(new_n582));
  INV_X1    g0382(.A(new_n580), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n577), .B1(new_n575), .B2(new_n574), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n213), .ZN(new_n585));
  OAI21_X1  g0385(.A(G107), .B1(new_n372), .B2(new_n374), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n587), .A2(new_n243), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n369), .A2(new_n538), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n477), .B2(new_n538), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n570), .B(new_n573), .C1(new_n588), .C2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n587), .B2(new_n243), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n567), .B1(new_n272), .B2(new_n564), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G190), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT78), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n565), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n564), .A2(KEYINPUT78), .A3(new_n272), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n567), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n592), .B(new_n594), .C1(new_n598), .C2(new_n486), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT79), .B1(new_n591), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n591), .A2(new_n599), .A3(KEYINPUT79), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n558), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n367), .A2(new_n433), .A3(new_n602), .ZN(G372));
  NOR2_X1   g0403(.A1(new_n367), .A2(new_n433), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n504), .A2(new_n516), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT85), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT85), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n504), .A2(new_n607), .A3(new_n516), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n514), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(new_n522), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n573), .A2(new_n570), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n611), .A2(KEYINPUT86), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(KEYINPUT86), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n612), .A2(new_n613), .A3(new_n592), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n517), .A2(new_n522), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(new_n591), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n556), .A2(new_n481), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n609), .A2(new_n489), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n591), .A2(new_n599), .ZN(new_n621));
  OAI221_X1 g0421(.A(new_n522), .B1(new_n615), .B2(new_n618), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n604), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n342), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n423), .A2(new_n413), .ZN(new_n625));
  INV_X1    g0425(.A(new_n365), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n337), .A2(new_n338), .B1(new_n626), .B2(new_n324), .ZN(new_n627));
  INV_X1    g0427(.A(new_n432), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n624), .B1(new_n629), .B2(new_n295), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n623), .A2(new_n630), .ZN(G369));
  NAND3_X1  g0431(.A1(new_n240), .A2(new_n213), .A3(G13), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n556), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(new_n481), .A3(new_n489), .ZN(new_n639));
  INV_X1    g0439(.A(new_n637), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n457), .A2(new_n480), .A3(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT87), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT87), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n543), .A2(new_n640), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n553), .B2(new_n555), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n557), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n480), .A2(new_n637), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n481), .A2(new_n650), .A3(new_n489), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n457), .A2(new_n480), .A3(new_n637), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n645), .A2(new_n656), .ZN(G399));
  INV_X1    g0457(.A(KEYINPUT88), .ZN(new_n658));
  INV_X1    g0458(.A(new_n207), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(G41), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n207), .A2(KEYINPUT88), .A3(new_n278), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n496), .A2(new_n497), .A3(new_n533), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n663), .A2(new_n240), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n211), .B2(new_n663), .ZN(new_n666));
  XOR2_X1   g0466(.A(new_n666), .B(KEYINPUT28), .Z(new_n667));
  OAI21_X1  g0467(.A(new_n640), .B1(new_n622), .B2(new_n616), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT29), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT90), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n618), .A2(new_n615), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n673), .B(new_n522), .C1(new_n620), .C2(new_n621), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n615), .B1(new_n610), .B2(new_n614), .ZN(new_n675));
  OAI211_X1 g0475(.A(KEYINPUT29), .B(new_n640), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n668), .A2(KEYINPUT90), .A3(new_n669), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n672), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n438), .A2(new_n525), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n272), .B2(new_n530), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G179), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n680), .A2(new_n515), .A3(new_n485), .A4(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT89), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n526), .A2(G179), .A3(new_n531), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n569), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n482), .A2(new_n443), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n515), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n685), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n684), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n593), .A2(new_n682), .A3(G179), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n455), .B(new_n506), .C1(new_n271), .C2(new_n513), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT89), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(KEYINPUT30), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n637), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n520), .A2(new_n515), .A3(new_n547), .A4(new_n485), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n695), .A2(KEYINPUT30), .B1(new_n680), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n690), .A2(new_n691), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT31), .B1(new_n703), .B2(new_n637), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n558), .B(new_n640), .C1(new_n600), .C2(new_n601), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n679), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n678), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n667), .B1(new_n710), .B2(G1), .ZN(G364));
  INV_X1    g0511(.A(G13), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n240), .B1(new_n713), .B2(G45), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n663), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n648), .B2(G330), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(G330), .B2(new_n648), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G13), .A2(G33), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n212), .B1(G20), .B2(new_n326), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n659), .A2(new_n263), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n279), .B2(new_n211), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n726), .A2(new_n727), .B1(new_n235), .B2(new_n279), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n727), .B2(new_n726), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n659), .A2(new_n371), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT91), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G355), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G116), .B2(new_n207), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n723), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n716), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n213), .A2(G179), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(G190), .A3(G200), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n286), .A3(G200), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n497), .A2(new_n737), .B1(new_n738), .B2(new_n351), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G190), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G159), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(KEYINPUT95), .B(KEYINPUT32), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n213), .A2(new_n520), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G200), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT94), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G190), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n739), .B(new_n745), .C1(G68), .C2(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n286), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n213), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n746), .A2(G190), .A3(new_n486), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(new_n740), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n252), .B1(new_n755), .B2(new_n202), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n263), .B1(new_n538), .B2(new_n753), .C1(new_n756), .C2(KEYINPUT93), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(KEYINPUT93), .B2(new_n756), .ZN(new_n758));
  INV_X1    g0558(.A(G50), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n749), .A2(new_n286), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n751), .B(new_n758), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G326), .A2(new_n760), .B1(new_n750), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G294), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n753), .A2(new_n765), .B1(new_n738), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n737), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G303), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n741), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT96), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT96), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n371), .B1(new_n755), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n754), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n777), .B1(G322), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n764), .A2(new_n769), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n762), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n735), .B1(new_n722), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n721), .B(KEYINPUT97), .Z(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n648), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n718), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NOR2_X1   g0586(.A1(new_n722), .A2(new_n719), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT98), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n716), .B1(new_n788), .B2(G77), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT99), .Z(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n755), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n778), .A2(G143), .B1(new_n792), .B2(G159), .ZN(new_n793));
  INV_X1    g0593(.A(new_n750), .ZN(new_n794));
  INV_X1    g0594(.A(G137), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n793), .B1(new_n794), .B2(new_n247), .C1(new_n795), .C2(new_n761), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT34), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n738), .A2(new_n311), .ZN(new_n798));
  INV_X1    g0598(.A(new_n753), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(G58), .B2(new_n799), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n800), .B(new_n263), .C1(new_n759), .C2(new_n737), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G132), .B2(new_n774), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G283), .A2(new_n750), .B1(new_n760), .B2(G303), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n753), .A2(new_n538), .B1(new_n737), .B2(new_n351), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n738), .A2(new_n497), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n774), .A2(G311), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n371), .B1(new_n755), .B2(new_n533), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G294), .B2(new_n778), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n804), .A2(new_n807), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n803), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n791), .B1(new_n812), .B2(new_n722), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n640), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n358), .A2(new_n360), .B1(new_n362), .B2(new_n637), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n626), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n719), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n668), .A2(new_n816), .ZN(new_n819));
  INV_X1    g0619(.A(new_n816), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n640), .B(new_n820), .C1(new_n622), .C2(new_n616), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n708), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT100), .Z(new_n824));
  AOI21_X1  g0624(.A(new_n716), .B1(new_n822), .B2(new_n708), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n818), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G384));
  NOR2_X1   g0627(.A1(new_n713), .A2(new_n240), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n418), .A2(new_n429), .A3(new_n370), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n419), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  INV_X1    g0631(.A(new_n635), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n395), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n830), .A2(KEYINPUT101), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n427), .A2(new_n429), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n421), .A2(new_n833), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT101), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n391), .A2(new_n393), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n635), .B1(new_n840), .B2(new_n370), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n427), .B2(new_n429), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n370), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n412), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n831), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n433), .A2(new_n841), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n421), .A2(new_n833), .A3(new_n835), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n834), .A2(new_n838), .B1(KEYINPUT37), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n833), .B1(new_n625), .B2(new_n432), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT39), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n849), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n845), .B1(new_n834), .B2(new_n838), .ZN(new_n858));
  INV_X1    g0658(.A(new_n841), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n424), .B2(new_n432), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n857), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n855), .B1(new_n849), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT103), .B1(new_n856), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n337), .A2(new_n338), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n637), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT38), .B1(new_n847), .B2(new_n848), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n858), .A2(new_n860), .A3(new_n857), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT39), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT103), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n849), .A2(new_n854), .A3(new_n855), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n863), .A2(new_n865), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n625), .A2(new_n832), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n821), .A2(new_n814), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n338), .A2(new_n637), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n864), .A2(new_n324), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n338), .B(new_n637), .C1(new_n337), .C2(new_n325), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n849), .A2(new_n861), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n873), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n672), .A2(new_n676), .A3(new_n604), .A4(new_n677), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n630), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n883), .B(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT104), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n640), .B1(new_n701), .B2(new_n702), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n888), .B2(KEYINPUT31), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(KEYINPUT31), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n697), .A2(KEYINPUT104), .A3(new_n698), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n706), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n816), .B1(new_n876), .B2(new_n877), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n866), .B2(new_n867), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n849), .A2(new_n854), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n892), .A2(new_n893), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT105), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n898), .A2(new_n901), .A3(KEYINPUT40), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n604), .A2(new_n892), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n906), .A2(new_n907), .A3(new_n679), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n828), .B1(new_n886), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n886), .B2(new_n909), .ZN(new_n911));
  INV_X1    g0711(.A(new_n584), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n912), .A2(KEYINPUT35), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(KEYINPUT35), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n913), .A2(G116), .A3(new_n214), .A4(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT36), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n376), .A2(new_n210), .A3(new_n202), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n311), .A2(G50), .ZN(new_n918));
  OAI211_X1 g0718(.A(G1), .B(new_n712), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n916), .A3(new_n919), .ZN(G367));
  NAND2_X1  g0720(.A1(new_n231), .A2(new_n724), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(new_n723), .C1(new_n207), .C2(new_n345), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(KEYINPUT108), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(KEYINPUT108), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n716), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n738), .A2(new_n538), .ZN(new_n926));
  AOI22_X1  g0726(.A1(G283), .A2(new_n792), .B1(new_n770), .B2(G317), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n927), .B(new_n371), .C1(new_n529), .C2(new_n754), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n926), .B(new_n928), .C1(G107), .C2(new_n799), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n768), .A2(G116), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT46), .ZN(new_n931));
  AOI22_X1  g0731(.A1(G294), .A2(new_n750), .B1(new_n760), .B2(G311), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT109), .Z(new_n934));
  AOI22_X1  g0734(.A1(G143), .A2(new_n760), .B1(new_n750), .B2(G159), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n755), .A2(new_n759), .B1(new_n741), .B2(new_n795), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n371), .B(new_n936), .C1(G150), .C2(new_n778), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n738), .A2(new_n202), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n753), .A2(new_n311), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n938), .B(new_n939), .C1(G58), .C2(new_n768), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n935), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT47), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n923), .B(new_n925), .C1(new_n943), .C2(new_n722), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n504), .A2(new_n640), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n522), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n610), .B2(new_n945), .ZN(new_n947));
  INV_X1    g0747(.A(new_n783), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n614), .A2(new_n637), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n591), .B(new_n599), .C1(new_n592), .C2(new_n640), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n643), .B2(new_n644), .ZN(new_n955));
  XOR2_X1   g0755(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n643), .A2(new_n644), .A3(new_n954), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT44), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n655), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT44), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n958), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n955), .A2(new_n956), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n955), .A2(new_n956), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n962), .A2(new_n656), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n653), .A2(new_n638), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT107), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n639), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(new_n649), .Z(new_n973));
  AOI21_X1  g0773(.A(new_n709), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n662), .B(KEYINPUT41), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n714), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n953), .A2(new_n481), .A3(new_n489), .A4(new_n638), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT42), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n953), .A2(new_n457), .A3(new_n480), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n637), .B1(new_n979), .B2(new_n591), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT43), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n978), .A2(new_n980), .B1(new_n981), .B2(new_n947), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n947), .A2(new_n981), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n655), .A2(new_n953), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n950), .B1(new_n976), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(G387));
  OR2_X1    g0788(.A1(new_n710), .A2(new_n973), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n710), .A2(new_n973), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n663), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n654), .A2(new_n948), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n724), .B1(new_n228), .B2(new_n279), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n731), .A2(new_n664), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n343), .A2(new_n759), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n998));
  AOI211_X1 g0798(.A(G45), .B(new_n664), .C1(G68), .C2(G77), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n995), .A2(new_n1000), .B1(new_n351), .B2(new_n659), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n723), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n716), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n778), .A2(G50), .B1(new_n792), .B2(G68), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n345), .B2(new_n753), .C1(new_n761), .C2(new_n742), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n256), .B2(new_n750), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n737), .A2(new_n202), .B1(new_n741), .B2(new_n247), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n371), .B(new_n926), .C1(new_n1007), .C2(KEYINPUT110), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(KEYINPUT110), .B2(new_n1007), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT111), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n263), .B1(new_n770), .B2(G326), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n753), .A2(new_n766), .B1(new_n737), .B2(new_n765), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n778), .A2(G317), .B1(new_n792), .B2(G303), .ZN(new_n1014));
  INV_X1    g0814(.A(G322), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1014), .B1(new_n794), .B2(new_n776), .C1(new_n1015), .C2(new_n761), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1012), .B1(new_n533), .B2(new_n738), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1011), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1003), .B1(new_n1023), .B2(new_n722), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n973), .A2(new_n715), .B1(new_n992), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n991), .A2(new_n1025), .ZN(G393));
  NAND2_X1  g0826(.A1(new_n967), .A2(new_n715), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n954), .A2(new_n721), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n371), .B1(new_n741), .B2(new_n1015), .C1(new_n765), .C2(new_n755), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n737), .A2(new_n766), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n753), .A2(new_n533), .B1(new_n738), .B2(new_n351), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n794), .B2(new_n529), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n760), .A2(G317), .B1(G311), .B2(new_n778), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT52), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n760), .A2(G150), .B1(G159), .B2(new_n778), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT51), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n770), .A2(G143), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n371), .B(new_n1038), .C1(new_n343), .C2(new_n792), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n737), .A2(new_n311), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n806), .B(new_n1040), .C1(G77), .C2(new_n799), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1039), .B(new_n1041), .C1(new_n759), .C2(new_n794), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1033), .A2(new_n1035), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n722), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n723), .B1(new_n538), .B2(new_n207), .C1(new_n238), .C2(new_n725), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1028), .A2(new_n716), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n990), .A2(new_n966), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n663), .B1(new_n990), .B2(new_n966), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1027), .B(new_n1046), .C1(new_n1048), .C2(new_n1049), .ZN(G390));
  AND3_X1   g0850(.A1(new_n892), .A2(new_n893), .A3(G330), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n865), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n863), .A2(new_n871), .B1(new_n1052), .B2(new_n879), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n815), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n365), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n640), .B(new_n1055), .C1(new_n674), .C2(new_n675), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1056), .A2(new_n814), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n878), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n1059), .A2(new_n1052), .A3(new_n898), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1051), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n879), .A2(new_n1052), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n856), .A2(new_n862), .A3(KEYINPUT103), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1059), .A2(new_n1052), .A3(new_n898), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n704), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n706), .A3(new_n890), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1068), .A2(G330), .A3(new_n820), .A4(new_n878), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1065), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1061), .A2(new_n1070), .A3(new_n715), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n719), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n716), .B1(new_n788), .B2(new_n256), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G107), .A2(new_n750), .B1(new_n760), .B2(G283), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n753), .A2(new_n202), .B1(new_n754), .B2(new_n533), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT116), .Z(new_n1076));
  NAND2_X1  g0876(.A1(new_n774), .A2(G294), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n371), .B1(new_n755), .B2(new_n538), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n798), .B(new_n1078), .C1(G87), .C2(new_n768), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(KEYINPUT54), .B(G143), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n753), .A2(new_n742), .B1(new_n755), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n750), .B2(G137), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT115), .Z(new_n1084));
  INV_X1    g0884(.A(G132), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n263), .B1(new_n754), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n768), .A2(G150), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(KEYINPUT53), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n738), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1086), .B(new_n1088), .C1(G50), .C2(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n774), .A2(G125), .B1(KEYINPUT53), .B2(new_n1087), .ZN(new_n1091));
  INV_X1    g0891(.A(G128), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1090), .B(new_n1091), .C1(new_n1092), .C2(new_n761), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1080), .B1(new_n1084), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1073), .B1(new_n1094), .B2(new_n722), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1072), .A2(new_n1095), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1071), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1061), .A2(new_n1070), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n878), .B1(new_n707), .B2(new_n820), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n874), .B1(new_n1099), .B2(new_n1051), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT112), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(KEYINPUT112), .B(new_n874), .C1(new_n1099), .C2(new_n1051), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n892), .A2(G330), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n878), .B1(new_n1104), .B2(new_n820), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1069), .A2(new_n814), .A3(new_n1056), .ZN(new_n1106));
  OAI21_X1  g0906(.A(KEYINPUT113), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n892), .A2(G330), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1058), .B1(new_n1108), .B2(new_n816), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT113), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n1057), .A4(new_n1069), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1102), .A2(new_n1103), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n604), .A2(new_n1104), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n884), .A2(new_n630), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT114), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1098), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1061), .A2(new_n1070), .A3(new_n1118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n663), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1097), .B1(new_n1121), .B2(new_n1123), .ZN(G378));
  INV_X1    g0924(.A(new_n1114), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT57), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n897), .A2(G330), .A3(new_n903), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n260), .A2(new_n832), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n295), .A2(new_n342), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n295), .B2(new_n342), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  OR3_X1    g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1128), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n897), .A2(new_n1136), .A3(G330), .A4(new_n903), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n883), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n872), .A3(new_n882), .A4(new_n1139), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1127), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1126), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n663), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT57), .B1(new_n1126), .B2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n715), .B(new_n663), .C1(new_n759), .C2(new_n787), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT119), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1136), .A2(new_n720), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n538), .A2(new_n794), .B1(new_n761), .B2(new_n533), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n939), .B1(G77), .B2(new_n768), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n252), .B2(new_n738), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n773), .A2(new_n766), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n263), .A2(G41), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n755), .B2(new_n345), .C1(new_n351), .C2(new_n754), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .A4(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n759), .B1(G33), .B2(G41), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1158), .A2(KEYINPUT58), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT117), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(KEYINPUT58), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n753), .A2(new_n247), .B1(new_n755), .B2(new_n795), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n760), .B2(G125), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n754), .A2(new_n1092), .B1(new_n737), .B2(new_n1081), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT118), .Z(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(new_n1085), .C2(new_n794), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1089), .A2(G159), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n770), .C2(G124), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1163), .B1(KEYINPUT117), .B2(new_n1160), .C1(new_n1169), .C2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1150), .B(new_n1151), .C1(new_n722), .C2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1146), .B2(new_n715), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1148), .A2(new_n1176), .ZN(G375));
  NAND2_X1  g0977(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(new_n1125), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n975), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1115), .A4(new_n1120), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1058), .A2(new_n719), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n716), .B1(new_n788), .B2(G68), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n753), .A2(new_n345), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n938), .B(new_n1185), .C1(G97), .C2(new_n768), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n371), .B1(new_n754), .B2(new_n766), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G107), .B2(new_n792), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(new_n529), .C2(new_n773), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n533), .A2(new_n794), .B1(new_n761), .B2(new_n765), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1085), .A2(new_n761), .B1(new_n794), .B2(new_n1081), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n252), .A2(new_n738), .B1(new_n737), .B2(new_n742), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G50), .B2(new_n799), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n263), .B1(new_n755), .B2(new_n247), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G137), .B2(new_n778), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(new_n1092), .C2(new_n773), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1189), .A2(new_n1190), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1184), .B1(new_n1197), .B2(new_n722), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1178), .A2(new_n715), .B1(new_n1183), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1182), .A2(new_n1199), .ZN(G381));
  INV_X1    g1000(.A(G375), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1071), .A2(new_n1096), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1123), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1098), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1046), .B1(new_n966), .B2(new_n714), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1049), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1206), .B1(new_n1207), .B2(new_n1047), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n990), .A2(new_n663), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n710), .A2(new_n973), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n785), .B(new_n1025), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1208), .A2(new_n826), .A3(new_n1212), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(G387), .A2(G381), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1201), .A2(new_n1205), .A3(new_n1214), .ZN(G407));
  NAND2_X1  g1015(.A1(new_n636), .A2(G213), .ZN(new_n1216));
  OR3_X1    g1016(.A1(G375), .A2(G378), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(G407), .A3(G213), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT120), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1218), .B(new_n1219), .ZN(G409));
  INV_X1    g1020(.A(KEYINPUT123), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n785), .B1(new_n991), .B2(new_n1025), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1208), .B1(new_n1212), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(G390), .A3(new_n1211), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1223), .A2(new_n1225), .A3(new_n987), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n987), .B1(new_n1225), .B2(new_n1223), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1221), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(G387), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1223), .A2(new_n1225), .A3(new_n987), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(KEYINPUT123), .A3(new_n1231), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1228), .A2(new_n1232), .A3(KEYINPUT124), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT124), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(G378), .B(new_n1176), .C1(new_n1145), .C2(new_n1147), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1126), .A2(new_n1146), .A3(new_n1181), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1176), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1205), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1112), .A2(KEYINPUT60), .A3(new_n1114), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n663), .ZN(new_n1242));
  OAI21_X1  g1042(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1180), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1199), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n826), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1243), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(new_n1179), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G384), .B(new_n1199), .C1(new_n1248), .C2(new_n1242), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1240), .A2(new_n1216), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT121), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1240), .A2(KEYINPUT121), .A3(new_n1216), .A4(new_n1250), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT62), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1240), .A2(new_n1216), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n636), .A2(G213), .A3(G2897), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT122), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1246), .A2(new_n1258), .A3(new_n1249), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1257), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1246), .A2(new_n1258), .A3(new_n1249), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1257), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1256), .A2(new_n1261), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1251), .A2(KEYINPUT62), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1235), .B1(new_n1255), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1253), .A2(new_n1270), .A3(new_n1254), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1240), .A2(new_n1216), .B1(new_n1263), .B2(new_n1262), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT61), .B1(new_n1274), .B2(new_n1261), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1251), .A2(new_n1270), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1271), .A2(new_n1273), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1269), .A2(new_n1277), .ZN(G405));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1250), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(KEYINPUT126), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1250), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G375), .A2(new_n1205), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(new_n1236), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1236), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1228), .A2(new_n1232), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1286), .A2(new_n1288), .A3(new_n1232), .A4(new_n1228), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(G402));
endmodule


