

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(G2105), .A2(n518), .ZN(n987) );
  AND2_X2 U551 ( .A1(n769), .A2(n675), .ZN(n712) );
  AND2_X1 U552 ( .A1(n712), .A2(G1996), .ZN(n680) );
  NOR2_X1 U553 ( .A1(n683), .A2(n999), .ZN(n684) );
  XNOR2_X1 U554 ( .A(n698), .B(KEYINPUT92), .ZN(n699) );
  XNOR2_X1 U555 ( .A(n700), .B(n699), .ZN(n702) );
  NOR2_X1 U556 ( .A1(n723), .A2(n722), .ZN(n724) );
  INV_X1 U557 ( .A(n768), .ZN(n675) );
  INV_X1 U558 ( .A(KEYINPUT102), .ZN(n756) );
  NOR2_X1 U559 ( .A1(G2104), .A2(n517), .ZN(n981) );
  NOR2_X1 U560 ( .A1(G651), .A2(n634), .ZN(n640) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n643) );
  NOR2_X1 U562 ( .A1(n518), .A2(n517), .ZN(n982) );
  INV_X1 U563 ( .A(G2105), .ZN(n517) );
  NAND2_X1 U564 ( .A1(G126), .A2(n981), .ZN(n515) );
  XNOR2_X1 U565 ( .A(KEYINPUT83), .B(n515), .ZN(n525) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XOR2_X2 U567 ( .A(KEYINPUT17), .B(n516), .Z(n985) );
  NAND2_X1 U568 ( .A1(G138), .A2(n985), .ZN(n523) );
  INV_X1 U569 ( .A(G2104), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n982), .A2(G114), .ZN(n521) );
  NAND2_X1 U571 ( .A1(G102), .A2(n987), .ZN(n519) );
  XNOR2_X1 U572 ( .A(n519), .B(KEYINPUT84), .ZN(n520) );
  AND2_X1 U573 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U574 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n527) );
  INV_X1 U576 ( .A(KEYINPUT85), .ZN(n526) );
  XNOR2_X1 U577 ( .A(n527), .B(n526), .ZN(G164) );
  NAND2_X1 U578 ( .A1(G113), .A2(n982), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G137), .A2(n985), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U581 ( .A(KEYINPUT66), .B(n530), .ZN(n537) );
  NAND2_X1 U582 ( .A1(n987), .A2(G101), .ZN(n531) );
  XOR2_X1 U583 ( .A(KEYINPUT23), .B(n531), .Z(n533) );
  NAND2_X1 U584 ( .A1(n981), .A2(G125), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n535) );
  INV_X1 U586 ( .A(KEYINPUT65), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n535), .B(n534), .ZN(n536) );
  NOR2_X2 U588 ( .A1(n537), .A2(n536), .ZN(G160) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U590 ( .A1(G123), .A2(n981), .ZN(n538) );
  XNOR2_X1 U591 ( .A(n538), .B(KEYINPUT18), .ZN(n545) );
  NAND2_X1 U592 ( .A1(G111), .A2(n982), .ZN(n540) );
  NAND2_X1 U593 ( .A1(G135), .A2(n985), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n543) );
  NAND2_X1 U595 ( .A1(G99), .A2(n987), .ZN(n541) );
  XNOR2_X1 U596 ( .A(KEYINPUT75), .B(n541), .ZN(n542) );
  NOR2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n971) );
  XNOR2_X1 U599 ( .A(G2096), .B(n971), .ZN(n546) );
  OR2_X1 U600 ( .A1(G2100), .A2(n546), .ZN(G156) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  NAND2_X1 U603 ( .A1(G88), .A2(n643), .ZN(n548) );
  XOR2_X1 U604 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  INV_X1 U605 ( .A(G651), .ZN(n549) );
  NOR2_X1 U606 ( .A1(n634), .A2(n549), .ZN(n637) );
  NAND2_X1 U607 ( .A1(G75), .A2(n637), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n554) );
  NOR2_X1 U609 ( .A1(G543), .A2(n549), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT1), .B(n550), .Z(n639) );
  NAND2_X1 U611 ( .A1(G62), .A2(n639), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G50), .A2(n640), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U614 ( .A1(n554), .A2(n553), .ZN(G166) );
  NAND2_X1 U615 ( .A1(G64), .A2(n639), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G52), .A2(n640), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G90), .A2(n643), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G77), .A2(n637), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U622 ( .A1(n561), .A2(n560), .ZN(G171) );
  NAND2_X1 U623 ( .A1(G63), .A2(n639), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G51), .A2(n640), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(KEYINPUT6), .B(n564), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n643), .A2(G89), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G76), .A2(n637), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U631 ( .A(n568), .B(KEYINPUT5), .Z(n569) );
  NOR2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT72), .B(n571), .Z(n572) );
  XNOR2_X1 U634 ( .A(KEYINPUT7), .B(n572), .ZN(G168) );
  XOR2_X1 U635 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n573) );
  XOR2_X1 U637 ( .A(n573), .B(KEYINPUT10), .Z(n1021) );
  NAND2_X1 U638 ( .A1(n1021), .A2(G567), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U640 ( .A1(n643), .A2(G81), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G68), .A2(n637), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n578), .Z(n582) );
  NAND2_X1 U645 ( .A1(G56), .A2(n639), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(KEYINPUT69), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT14), .ZN(n581) );
  NOR2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n640), .A2(G43), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n999) );
  INV_X1 U651 ( .A(G860), .ZN(n605) );
  OR2_X1 U652 ( .A1(n999), .A2(n605), .ZN(G153) );
  INV_X1 U653 ( .A(G171), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G301), .A2(G868), .ZN(n585) );
  XNOR2_X1 U655 ( .A(n585), .B(KEYINPUT70), .ZN(n595) );
  NAND2_X1 U656 ( .A1(G79), .A2(n637), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G66), .A2(n639), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G92), .A2(n643), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G54), .A2(n640), .ZN(n588) );
  XNOR2_X1 U661 ( .A(KEYINPUT71), .B(n588), .ZN(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n593), .B(KEYINPUT15), .ZN(n1002) );
  OR2_X1 U665 ( .A1(G868), .A2(n1002), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G65), .A2(n639), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G53), .A2(n640), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G91), .A2(n643), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G78), .A2(n637), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n706) );
  INV_X1 U674 ( .A(n706), .ZN(G299) );
  INV_X1 U675 ( .A(G868), .ZN(n656) );
  XOR2_X1 U676 ( .A(KEYINPUT73), .B(n656), .Z(n602) );
  NOR2_X1 U677 ( .A1(G286), .A2(n602), .ZN(n604) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U679 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n606), .A2(n1002), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U683 ( .A1(n1002), .A2(G868), .ZN(n608) );
  XNOR2_X1 U684 ( .A(KEYINPUT74), .B(n608), .ZN(n609) );
  NOR2_X1 U685 ( .A1(G559), .A2(n609), .ZN(n611) );
  NOR2_X1 U686 ( .A1(G868), .A2(n999), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G559), .A2(n1002), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(n999), .ZN(n654) );
  NOR2_X1 U690 ( .A1(n654), .A2(G860), .ZN(n622) );
  NAND2_X1 U691 ( .A1(G93), .A2(n643), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT76), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G55), .A2(n640), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G80), .A2(n637), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G67), .A2(n639), .ZN(n616) );
  XNOR2_X1 U697 ( .A(KEYINPUT77), .B(n616), .ZN(n617) );
  NOR2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n657) );
  XOR2_X1 U700 ( .A(n657), .B(KEYINPUT78), .Z(n621) );
  XNOR2_X1 U701 ( .A(n622), .B(n621), .ZN(G145) );
  NAND2_X1 U702 ( .A1(G60), .A2(n639), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G47), .A2(n640), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U705 ( .A(KEYINPUT67), .B(n625), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G85), .A2(n643), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G72), .A2(n637), .ZN(n626) );
  AND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G290) );
  NAND2_X1 U710 ( .A1(G49), .A2(n640), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n639), .A2(n632), .ZN(n633) );
  XOR2_X1 U714 ( .A(KEYINPUT79), .B(n633), .Z(n636) );
  NAND2_X1 U715 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U717 ( .A1(G73), .A2(n637), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n638), .B(KEYINPUT2), .ZN(n648) );
  NAND2_X1 U719 ( .A1(G61), .A2(n639), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G48), .A2(n640), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n643), .A2(G86), .ZN(n644) );
  XOR2_X1 U723 ( .A(KEYINPUT80), .B(n644), .Z(n645) );
  NOR2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(G305) );
  XNOR2_X1 U726 ( .A(G290), .B(G288), .ZN(n653) );
  XOR2_X1 U727 ( .A(KEYINPUT19), .B(G166), .Z(n649) );
  XNOR2_X1 U728 ( .A(n649), .B(n657), .ZN(n650) );
  XOR2_X1 U729 ( .A(G299), .B(n650), .Z(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(G305), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n1000) );
  XNOR2_X1 U732 ( .A(n654), .B(n1000), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n655), .A2(G868), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XOR2_X1 U741 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U743 ( .A1(G219), .A2(G220), .ZN(n665) );
  XNOR2_X1 U744 ( .A(KEYINPUT22), .B(KEYINPUT81), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U746 ( .A1(n666), .A2(G218), .ZN(n667) );
  NAND2_X1 U747 ( .A1(G96), .A2(n667), .ZN(n949) );
  NAND2_X1 U748 ( .A1(G2106), .A2(n949), .ZN(n672) );
  NAND2_X1 U749 ( .A1(G120), .A2(G69), .ZN(n668) );
  NOR2_X1 U750 ( .A1(G237), .A2(n668), .ZN(n669) );
  XNOR2_X1 U751 ( .A(KEYINPUT82), .B(n669), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n670), .A2(G108), .ZN(n948) );
  NAND2_X1 U753 ( .A1(G567), .A2(n948), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(n950) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n673) );
  NOR2_X1 U756 ( .A1(n950), .A2(n673), .ZN(n831) );
  NAND2_X1 U757 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U758 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U759 ( .A(G1981), .B(KEYINPUT101), .ZN(n674) );
  XNOR2_X1 U760 ( .A(n674), .B(G305), .ZN(n910) );
  NOR2_X1 U761 ( .A1(G164), .A2(G1384), .ZN(n769) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n768) );
  INV_X1 U763 ( .A(n712), .ZN(n689) );
  NAND2_X1 U764 ( .A1(G8), .A2(n689), .ZN(n767) );
  NOR2_X1 U765 ( .A1(G288), .A2(G1976), .ZN(n676) );
  XOR2_X1 U766 ( .A(n676), .B(KEYINPUT99), .Z(n747) );
  INV_X1 U767 ( .A(n747), .ZN(n905) );
  NOR2_X1 U768 ( .A1(n767), .A2(n905), .ZN(n677) );
  NAND2_X1 U769 ( .A1(KEYINPUT33), .A2(n677), .ZN(n678) );
  NAND2_X1 U770 ( .A1(n910), .A2(n678), .ZN(n755) );
  XNOR2_X1 U771 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n679) );
  XNOR2_X1 U772 ( .A(n680), .B(n679), .ZN(n682) );
  NAND2_X1 U773 ( .A1(n689), .A2(G1341), .ZN(n681) );
  NAND2_X1 U774 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U775 ( .A(n684), .B(KEYINPUT64), .ZN(n687) );
  NOR2_X1 U776 ( .A1(n1002), .A2(n687), .ZN(n686) );
  INV_X1 U777 ( .A(KEYINPUT98), .ZN(n685) );
  XNOR2_X1 U778 ( .A(n686), .B(n685), .ZN(n696) );
  NAND2_X1 U779 ( .A1(n1002), .A2(n687), .ZN(n694) );
  NAND2_X1 U780 ( .A1(G2067), .A2(n712), .ZN(n688) );
  XNOR2_X1 U781 ( .A(n688), .B(KEYINPUT96), .ZN(n691) );
  NAND2_X1 U782 ( .A1(G1348), .A2(n689), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U784 ( .A(KEYINPUT97), .B(n692), .Z(n693) );
  NAND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n704) );
  NAND2_X1 U787 ( .A1(G2072), .A2(n712), .ZN(n697) );
  XNOR2_X1 U788 ( .A(KEYINPUT27), .B(n697), .ZN(n700) );
  INV_X1 U789 ( .A(KEYINPUT93), .ZN(n698) );
  XOR2_X1 U790 ( .A(G1956), .B(KEYINPUT94), .Z(n917) );
  NOR2_X1 U791 ( .A1(n712), .A2(n917), .ZN(n701) );
  NOR2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U793 ( .A1(n706), .A2(n705), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n709) );
  NOR2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U796 ( .A(n707), .B(KEYINPUT28), .Z(n708) );
  NAND2_X1 U797 ( .A1(n709), .A2(n708), .ZN(n711) );
  INV_X1 U798 ( .A(KEYINPUT29), .ZN(n710) );
  XNOR2_X1 U799 ( .A(n711), .B(n710), .ZN(n717) );
  INV_X1 U800 ( .A(G1961), .ZN(n965) );
  NAND2_X1 U801 ( .A1(n689), .A2(n965), .ZN(n714) );
  XNOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .ZN(n850) );
  NAND2_X1 U803 ( .A1(n712), .A2(n850), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n721) );
  AND2_X1 U805 ( .A1(n721), .A2(G171), .ZN(n715) );
  XNOR2_X1 U806 ( .A(KEYINPUT91), .B(n715), .ZN(n716) );
  NAND2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n738) );
  INV_X1 U808 ( .A(KEYINPUT31), .ZN(n725) );
  NOR2_X1 U809 ( .A1(G1966), .A2(n767), .ZN(n727) );
  NOR2_X1 U810 ( .A1(G2084), .A2(n689), .ZN(n726) );
  NOR2_X1 U811 ( .A1(n727), .A2(n726), .ZN(n718) );
  NAND2_X1 U812 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U813 ( .A(KEYINPUT30), .B(n719), .ZN(n720) );
  NOR2_X1 U814 ( .A1(G168), .A2(n720), .ZN(n723) );
  NOR2_X1 U815 ( .A1(G171), .A2(n721), .ZN(n722) );
  XNOR2_X1 U816 ( .A(n725), .B(n724), .ZN(n736) );
  AND2_X1 U817 ( .A1(n738), .A2(n736), .ZN(n730) );
  AND2_X1 U818 ( .A1(G8), .A2(n726), .ZN(n728) );
  OR2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n729) );
  OR2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n745) );
  INV_X1 U821 ( .A(G8), .ZN(n735) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n767), .ZN(n732) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n689), .ZN(n731) );
  NOR2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U825 ( .A1(n733), .A2(G303), .ZN(n734) );
  OR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n739) );
  AND2_X1 U827 ( .A1(n736), .A2(n739), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n742) );
  INV_X1 U829 ( .A(n739), .ZN(n740) );
  OR2_X1 U830 ( .A1(n740), .A2(G286), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U832 ( .A(n743), .B(KEYINPUT32), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n758) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n746) );
  NOR2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n758), .A2(n748), .ZN(n749) );
  XNOR2_X1 U837 ( .A(n749), .B(KEYINPUT100), .ZN(n752) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n896) );
  INV_X1 U839 ( .A(n896), .ZN(n750) );
  NOR2_X1 U840 ( .A1(n767), .A2(n750), .ZN(n751) );
  AND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n753), .A2(KEYINPUT33), .ZN(n754) );
  NOR2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n757) );
  XNOR2_X1 U844 ( .A(n757), .B(n756), .ZN(n815) );
  INV_X1 U845 ( .A(n758), .ZN(n761) );
  NAND2_X1 U846 ( .A1(G166), .A2(G8), .ZN(n759) );
  NOR2_X1 U847 ( .A1(G2090), .A2(n759), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U849 ( .A(KEYINPUT103), .B(n762), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n763), .A2(n767), .ZN(n813) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U852 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  XNOR2_X1 U853 ( .A(KEYINPUT90), .B(n765), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n811) );
  NOR2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n816) );
  NAND2_X1 U856 ( .A1(G140), .A2(n985), .ZN(n771) );
  NAND2_X1 U857 ( .A1(G104), .A2(n987), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(n772), .ZN(n777) );
  NAND2_X1 U860 ( .A1(G128), .A2(n981), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G116), .A2(n982), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U863 ( .A(n775), .B(KEYINPUT35), .Z(n776) );
  NOR2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U865 ( .A(KEYINPUT36), .B(n778), .Z(n779) );
  XOR2_X1 U866 ( .A(KEYINPUT86), .B(n779), .Z(n996) );
  XNOR2_X1 U867 ( .A(G2067), .B(KEYINPUT37), .ZN(n808) );
  OR2_X1 U868 ( .A1(n996), .A2(n808), .ZN(n780) );
  XNOR2_X1 U869 ( .A(n780), .B(KEYINPUT87), .ZN(n863) );
  NAND2_X1 U870 ( .A1(n816), .A2(n863), .ZN(n817) );
  NAND2_X1 U871 ( .A1(G129), .A2(n981), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G141), .A2(n985), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n987), .A2(G105), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n982), .A2(G117), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n970) );
  NOR2_X1 U879 ( .A1(G1996), .A2(n970), .ZN(n868) );
  XOR2_X1 U880 ( .A(KEYINPUT89), .B(n816), .Z(n797) );
  NAND2_X1 U881 ( .A1(G1996), .A2(n970), .ZN(n788) );
  XNOR2_X1 U882 ( .A(n788), .B(KEYINPUT88), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G119), .A2(n981), .ZN(n790) );
  NAND2_X1 U884 ( .A1(G107), .A2(n982), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U886 ( .A1(G131), .A2(n985), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G95), .A2(n987), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n793) );
  OR2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n974) );
  NAND2_X1 U890 ( .A1(G1991), .A2(n974), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n861) );
  NAND2_X1 U892 ( .A1(n797), .A2(n861), .ZN(n818) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n798) );
  XOR2_X1 U894 ( .A(n798), .B(KEYINPUT104), .Z(n800) );
  NOR2_X1 U895 ( .A1(G1991), .A2(n974), .ZN(n799) );
  XNOR2_X1 U896 ( .A(KEYINPUT105), .B(n799), .ZN(n859) );
  NAND2_X1 U897 ( .A1(n800), .A2(n859), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n818), .A2(n801), .ZN(n802) );
  XOR2_X1 U899 ( .A(KEYINPUT106), .B(n802), .Z(n803) );
  NOR2_X1 U900 ( .A1(n868), .A2(n803), .ZN(n804) );
  XOR2_X1 U901 ( .A(n804), .B(KEYINPUT107), .Z(n805) );
  XNOR2_X1 U902 ( .A(KEYINPUT39), .B(n805), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n817), .A2(n806), .ZN(n807) );
  XNOR2_X1 U904 ( .A(n807), .B(KEYINPUT108), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n996), .A2(n808), .ZN(n887) );
  NAND2_X1 U906 ( .A1(n809), .A2(n887), .ZN(n810) );
  AND2_X1 U907 ( .A1(n810), .A2(n816), .ZN(n822) );
  NOR2_X1 U908 ( .A1(n811), .A2(n822), .ZN(n812) );
  AND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n824) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n895) );
  AND2_X1 U912 ( .A1(n895), .A2(n816), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  OR2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U917 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n1021), .ZN(G217) );
  NAND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n826) );
  XNOR2_X1 U920 ( .A(KEYINPUT109), .B(n826), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n827), .A2(G661), .ZN(n828) );
  XNOR2_X1 U922 ( .A(KEYINPUT110), .B(n828), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n829) );
  XOR2_X1 U924 ( .A(KEYINPUT111), .B(n829), .Z(n830) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(G188) );
  NAND2_X1 U927 ( .A1(G112), .A2(n982), .ZN(n833) );
  NAND2_X1 U928 ( .A1(G100), .A2(n987), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n833), .A2(n832), .ZN(n839) );
  NAND2_X1 U930 ( .A1(G136), .A2(n985), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(KEYINPUT114), .ZN(n837) );
  NAND2_X1 U932 ( .A1(G124), .A2(n981), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n835), .B(KEYINPUT44), .ZN(n836) );
  NAND2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G162) );
  XOR2_X1 U936 ( .A(G2090), .B(G35), .Z(n842) );
  XOR2_X1 U937 ( .A(G34), .B(KEYINPUT54), .Z(n840) );
  XNOR2_X1 U938 ( .A(G2084), .B(n840), .ZN(n841) );
  NAND2_X1 U939 ( .A1(n842), .A2(n841), .ZN(n855) );
  XNOR2_X1 U940 ( .A(G1996), .B(G32), .ZN(n844) );
  XNOR2_X1 U941 ( .A(G33), .B(G2072), .ZN(n843) );
  NOR2_X1 U942 ( .A1(n844), .A2(n843), .ZN(n849) );
  XOR2_X1 U943 ( .A(G1991), .B(G25), .Z(n845) );
  NAND2_X1 U944 ( .A1(n845), .A2(G28), .ZN(n847) );
  XNOR2_X1 U945 ( .A(G26), .B(G2067), .ZN(n846) );
  NOR2_X1 U946 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n852) );
  XOR2_X1 U948 ( .A(G27), .B(n850), .Z(n851) );
  NOR2_X1 U949 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n853), .B(KEYINPUT53), .ZN(n854) );
  NOR2_X1 U951 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U952 ( .A(KEYINPUT122), .B(n856), .ZN(n857) );
  NOR2_X1 U953 ( .A1(G29), .A2(n857), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n858), .B(KEYINPUT55), .ZN(n893) );
  XOR2_X1 U955 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n890) );
  NAND2_X1 U956 ( .A1(n859), .A2(n971), .ZN(n860) );
  NOR2_X1 U957 ( .A1(n861), .A2(n860), .ZN(n865) );
  XOR2_X1 U958 ( .A(G160), .B(G2084), .Z(n862) );
  NOR2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n864) );
  NAND2_X1 U960 ( .A1(n865), .A2(n864), .ZN(n872) );
  XOR2_X1 U961 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n870) );
  XOR2_X1 U962 ( .A(G2090), .B(G162), .Z(n866) );
  XNOR2_X1 U963 ( .A(KEYINPUT118), .B(n866), .ZN(n867) );
  NOR2_X1 U964 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U965 ( .A(n870), .B(n869), .ZN(n871) );
  NOR2_X1 U966 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U967 ( .A(KEYINPUT120), .B(n873), .Z(n886) );
  NAND2_X1 U968 ( .A1(G139), .A2(n985), .ZN(n875) );
  NAND2_X1 U969 ( .A1(G103), .A2(n987), .ZN(n874) );
  NAND2_X1 U970 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U971 ( .A1(n981), .A2(G127), .ZN(n876) );
  XNOR2_X1 U972 ( .A(n876), .B(KEYINPUT116), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G115), .A2(n982), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U976 ( .A1(n881), .A2(n880), .ZN(n977) );
  XOR2_X1 U977 ( .A(G2072), .B(n977), .Z(n883) );
  XOR2_X1 U978 ( .A(G164), .B(G2078), .Z(n882) );
  NOR2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U980 ( .A(KEYINPUT50), .B(n884), .Z(n885) );
  NOR2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n888) );
  NAND2_X1 U982 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U983 ( .A(n890), .B(n889), .ZN(n891) );
  NAND2_X1 U984 ( .A1(G29), .A2(n891), .ZN(n892) );
  NAND2_X1 U985 ( .A1(n893), .A2(n892), .ZN(n945) );
  INV_X1 U986 ( .A(G16), .ZN(n940) );
  XOR2_X1 U987 ( .A(n940), .B(KEYINPUT56), .Z(n916) );
  XNOR2_X1 U988 ( .A(G1341), .B(n999), .ZN(n894) );
  NOR2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n901) );
  XOR2_X1 U990 ( .A(G299), .B(G1956), .Z(n897) );
  NAND2_X1 U991 ( .A1(n897), .A2(n896), .ZN(n899) );
  XOR2_X1 U992 ( .A(n1002), .B(G1348), .Z(n898) );
  NOR2_X1 U993 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U994 ( .A1(n901), .A2(n900), .ZN(n908) );
  XOR2_X1 U995 ( .A(G303), .B(G1971), .Z(n902) );
  XNOR2_X1 U996 ( .A(n902), .B(KEYINPUT123), .ZN(n904) );
  XOR2_X1 U997 ( .A(n965), .B(G301), .Z(n903) );
  NOR2_X1 U998 ( .A1(n904), .A2(n903), .ZN(n906) );
  NAND2_X1 U999 ( .A1(n906), .A2(n905), .ZN(n907) );
  NOR2_X1 U1000 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(KEYINPUT124), .B(n909), .ZN(n914) );
  XNOR2_X1 U1002 ( .A(G1966), .B(G168), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1004 ( .A(KEYINPUT57), .B(n912), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1006 ( .A1(n916), .A2(n915), .ZN(n942) );
  XOR2_X1 U1007 ( .A(G5), .B(G1961), .Z(n937) );
  XNOR2_X1 U1008 ( .A(n917), .B(G20), .ZN(n921) );
  XNOR2_X1 U1009 ( .A(G1341), .B(G19), .ZN(n919) );
  XNOR2_X1 U1010 ( .A(G6), .B(G1981), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1012 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1013 ( .A(KEYINPUT59), .B(G1348), .Z(n922) );
  XNOR2_X1 U1014 ( .A(G4), .B(n922), .ZN(n923) );
  NOR2_X1 U1015 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1016 ( .A(KEYINPUT60), .B(n925), .Z(n927) );
  XNOR2_X1 U1017 ( .A(G1966), .B(G21), .ZN(n926) );
  NOR2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(KEYINPUT125), .B(n928), .ZN(n935) );
  XNOR2_X1 U1020 ( .A(G1971), .B(G22), .ZN(n930) );
  XNOR2_X1 U1021 ( .A(G23), .B(G1976), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n932) );
  XOR2_X1 U1023 ( .A(G1986), .B(G24), .Z(n931) );
  NAND2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(KEYINPUT58), .B(n933), .ZN(n934) );
  NOR2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1028 ( .A(KEYINPUT61), .B(n938), .Z(n939) );
  NAND2_X1 U1029 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1030 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1031 ( .A(n943), .B(KEYINPUT126), .ZN(n944) );
  NOR2_X1 U1032 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1033 ( .A1(n946), .A2(G11), .ZN(n947) );
  XOR2_X1 U1034 ( .A(KEYINPUT62), .B(n947), .Z(G311) );
  XNOR2_X1 U1035 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1036 ( .A(G120), .ZN(G236) );
  INV_X1 U1037 ( .A(G108), .ZN(G238) );
  INV_X1 U1038 ( .A(G96), .ZN(G221) );
  INV_X1 U1039 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(G325) );
  INV_X1 U1041 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1042 ( .A(KEYINPUT112), .B(n950), .Z(G319) );
  XOR2_X1 U1043 ( .A(KEYINPUT113), .B(G2678), .Z(n952) );
  XNOR2_X1 U1044 ( .A(G2078), .B(G2084), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(n952), .B(n951), .ZN(n953) );
  XOR2_X1 U1046 ( .A(n953), .B(KEYINPUT42), .Z(n955) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G2072), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(n955), .B(n954), .ZN(n959) );
  XOR2_X1 U1049 ( .A(G2100), .B(G2096), .Z(n957) );
  XNOR2_X1 U1050 ( .A(G2090), .B(KEYINPUT43), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n957), .B(n956), .ZN(n958) );
  XOR2_X1 U1052 ( .A(n959), .B(n958), .Z(G227) );
  XOR2_X1 U1053 ( .A(KEYINPUT41), .B(G1971), .Z(n961) );
  XNOR2_X1 U1054 ( .A(G1986), .B(G1966), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n961), .B(n960), .ZN(n962) );
  XOR2_X1 U1056 ( .A(n962), .B(G1976), .Z(n964) );
  XNOR2_X1 U1057 ( .A(G1991), .B(G1996), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n964), .B(n963), .ZN(n969) );
  XOR2_X1 U1059 ( .A(G2474), .B(G1981), .Z(n967) );
  XOR2_X1 U1060 ( .A(G1956), .B(n965), .Z(n966) );
  XNOR2_X1 U1061 ( .A(n967), .B(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(n969), .B(n968), .ZN(G229) );
  XNOR2_X1 U1063 ( .A(G162), .B(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n972), .B(n971), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(KEYINPUT48), .B(n973), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n974), .B(KEYINPUT46), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n976), .B(n975), .ZN(n978) );
  XOR2_X1 U1068 ( .A(n978), .B(n977), .Z(n980) );
  XNOR2_X1 U1069 ( .A(G164), .B(G160), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n980), .B(n979), .ZN(n994) );
  NAND2_X1 U1071 ( .A1(G130), .A2(n981), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(G118), .A2(n982), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n992) );
  NAND2_X1 U1074 ( .A1(n985), .A2(G142), .ZN(n986) );
  XOR2_X1 U1075 ( .A(KEYINPUT115), .B(n986), .Z(n989) );
  NAND2_X1 U1076 ( .A1(n987), .A2(G106), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1078 ( .A(n990), .B(KEYINPUT45), .Z(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1080 ( .A(n994), .B(n993), .Z(n995) );
  XOR2_X1 U1081 ( .A(n996), .B(n995), .Z(n997) );
  NOR2_X1 U1082 ( .A1(G37), .A2(n997), .ZN(n998) );
  XOR2_X1 U1083 ( .A(KEYINPUT117), .B(n998), .Z(G395) );
  XOR2_X1 U1084 ( .A(G301), .B(n999), .Z(n1001) );
  XNOR2_X1 U1085 ( .A(n1001), .B(n1000), .ZN(n1004) );
  XOR2_X1 U1086 ( .A(G286), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1087 ( .A(n1004), .B(n1003), .ZN(n1005) );
  NOR2_X1 U1088 ( .A1(G37), .A2(n1005), .ZN(G397) );
  XOR2_X1 U1089 ( .A(G2446), .B(G2451), .Z(n1007) );
  XNOR2_X1 U1090 ( .A(G1348), .B(G2430), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(n1007), .B(n1006), .ZN(n1013) );
  XOR2_X1 U1092 ( .A(G2443), .B(G2438), .Z(n1009) );
  XNOR2_X1 U1093 ( .A(G2454), .B(G2435), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(n1009), .B(n1008), .ZN(n1011) );
  XOR2_X1 U1095 ( .A(G1341), .B(G2427), .Z(n1010) );
  XNOR2_X1 U1096 ( .A(n1011), .B(n1010), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(n1013), .B(n1012), .Z(n1014) );
  NAND2_X1 U1098 ( .A1(G14), .A2(n1014), .ZN(n1020) );
  NAND2_X1 U1099 ( .A1(n1020), .A2(G319), .ZN(n1017) );
  NOR2_X1 U1100 ( .A1(G227), .A2(G229), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT49), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NOR2_X1 U1103 ( .A1(G395), .A2(G397), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(G225) );
  INV_X1 U1105 ( .A(G225), .ZN(G308) );
  INV_X1 U1106 ( .A(n1020), .ZN(G401) );
  INV_X1 U1107 ( .A(n1021), .ZN(G223) );
endmodule

