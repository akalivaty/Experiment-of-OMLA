//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g0008(.A(new_n208), .B1(G68), .B2(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n203), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n205), .B(new_n225), .C1(new_n207), .C2(new_n211), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(G58), .A2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n233), .A2(G50), .A3(new_n234), .ZN(new_n235));
  OAI22_X1  g0035(.A1(new_n226), .A2(KEYINPUT0), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT0), .B2(new_n226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n223), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n220), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT66), .B(G250), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G257), .ZN(new_n245));
  XOR2_X1   g0045(.A(G264), .B(G270), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n243), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT72), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n256), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G50), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n227), .B1(new_n203), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n259), .B2(new_n260), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G1), .B2(new_n228), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n214), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  XOR2_X1   g0069(.A(KEYINPUT8), .B(G58), .Z(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n264), .B2(G20), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n228), .A2(KEYINPUT69), .A3(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G150), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT70), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT70), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n274), .A2(new_n279), .A3(new_n276), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n232), .A2(G50), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n278), .B(new_n280), .C1(new_n228), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT71), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(new_n265), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n283), .B1(new_n282), .B2(new_n265), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n263), .B(new_n269), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n264), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G222), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT68), .B(G223), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n291), .B(new_n293), .C1(new_n294), .C2(new_n292), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n295), .B(new_n296), .C1(G77), .C2(new_n291), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G1), .A3(G13), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT67), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n302), .B(new_n256), .C1(G41), .C2(G45), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n299), .A2(G274), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n298), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G226), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n297), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G179), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n308), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n287), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n282), .A2(new_n265), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT71), .ZN(new_n314));
  AOI211_X1 g0114(.A(new_n262), .B(new_n268), .C1(new_n314), .C2(new_n284), .ZN(new_n315));
  INV_X1    g0115(.A(new_n308), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n315), .A2(KEYINPUT9), .B1(G190), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT9), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n287), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n308), .A2(G200), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n317), .A2(new_n318), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n320), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n316), .A2(G190), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n321), .B(new_n324), .C1(new_n287), .C2(new_n319), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT10), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n312), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT82), .ZN(new_n328));
  INV_X1    g0128(.A(new_n261), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n270), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n267), .B2(new_n270), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT16), .ZN(new_n332));
  INV_X1    g0132(.A(G68), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n289), .A2(new_n228), .A3(new_n290), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT7), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT80), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(KEYINPUT80), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT79), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n288), .A2(KEYINPUT79), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n264), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n344), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n290), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n333), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n219), .A2(new_n333), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n347), .B2(new_n231), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n275), .A2(G159), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n332), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n265), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n288), .A2(KEYINPUT79), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n354), .A3(G33), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(new_n228), .A3(new_n289), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n333), .B1(new_n356), .B2(KEYINPUT7), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n355), .A2(new_n335), .A3(new_n228), .A4(new_n289), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n350), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n352), .B1(new_n359), .B2(KEYINPUT16), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n331), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n303), .A2(new_n301), .A3(G274), .ZN(new_n363));
  INV_X1    g0163(.A(G41), .ZN(new_n364));
  INV_X1    g0164(.A(G45), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n302), .B1(new_n366), .B2(new_n256), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n363), .A2(new_n367), .B1(new_n305), .B2(new_n220), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT81), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n304), .B(KEYINPUT81), .C1(new_n220), .C2(new_n305), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n355), .A2(new_n289), .ZN(new_n373));
  OR2_X1    g0173(.A1(G223), .A2(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n215), .A2(G1698), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n264), .A2(new_n204), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n301), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n362), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(new_n378), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n296), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(new_n370), .A4(new_n371), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n361), .A2(KEYINPUT17), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT17), .B1(new_n361), .B2(new_n385), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n328), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(G169), .B1(new_n372), .B2(new_n379), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n382), .A2(G179), .A3(new_n370), .A4(new_n371), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n361), .A2(new_n391), .A3(KEYINPUT18), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n356), .A2(KEYINPUT7), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(G68), .A3(new_n358), .ZN(new_n395));
  INV_X1    g0195(.A(new_n350), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n334), .A2(KEYINPUT80), .A3(new_n335), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT80), .B1(new_n334), .B2(new_n335), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n345), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n350), .B1(new_n400), .B2(G68), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n265), .B(new_n397), .C1(new_n401), .C2(KEYINPUT16), .ZN(new_n402));
  INV_X1    g0202(.A(new_n331), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n389), .A2(new_n390), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n393), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n392), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n380), .A2(new_n384), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n361), .A2(KEYINPUT17), .A3(new_n385), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(KEYINPUT82), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n388), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n306), .A2(G238), .ZN(new_n414));
  NOR2_X1   g0214(.A1(G226), .A2(G1698), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n220), .B2(G1698), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(new_n291), .B1(G33), .B2(G97), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n414), .B(new_n304), .C1(new_n417), .C2(new_n301), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT13), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n418), .A2(KEYINPUT13), .ZN(new_n421));
  OAI21_X1  g0221(.A(G169), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(KEYINPUT78), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n418), .B(KEYINPUT13), .ZN(new_n426));
  INV_X1    g0226(.A(new_n424), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(G169), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n420), .A2(new_n421), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G179), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n425), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n272), .A2(G77), .A3(new_n273), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT75), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n333), .A2(G20), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n432), .B2(new_n434), .ZN(new_n436));
  INV_X1    g0236(.A(new_n275), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(new_n214), .ZN(new_n438));
  OR3_X1    g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g0239(.A(KEYINPUT76), .B(KEYINPUT11), .Z(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n265), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n440), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(new_n352), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n259), .A2(new_n333), .A3(new_n260), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n447), .A2(KEYINPUT12), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(KEYINPUT12), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n333), .B2(new_n267), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n446), .B1(new_n445), .B2(new_n452), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n431), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n426), .A2(G200), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n429), .A2(G190), .ZN(new_n458));
  AOI211_X1 g0258(.A(KEYINPUT77), .B(new_n451), .C1(new_n441), .C2(new_n444), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(new_n454), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n413), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n291), .A2(G232), .A3(new_n292), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT73), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n291), .A2(G238), .A3(G1698), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n465), .B(new_n466), .C1(new_n210), .C2(new_n291), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n296), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n306), .A2(G244), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n468), .A2(new_n304), .A3(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n470), .A2(new_n362), .ZN(new_n471));
  OR3_X1    g0271(.A1(new_n261), .A2(KEYINPUT74), .A3(G77), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT74), .B1(new_n261), .B2(G77), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n272), .A2(new_n273), .ZN(new_n475));
  XOR2_X1   g0275(.A(KEYINPUT15), .B(G87), .Z(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n270), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n475), .A2(new_n477), .B1(new_n478), .B2(new_n437), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(G20), .B2(G77), .ZN(new_n480));
  OAI221_X1 g0280(.A(new_n474), .B1(new_n216), .B2(new_n267), .C1(new_n480), .C2(new_n352), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n470), .B2(G190), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n471), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G179), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n468), .A2(new_n484), .A3(new_n304), .A4(new_n469), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n481), .B(new_n485), .C1(new_n470), .C2(G169), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n327), .A2(new_n462), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n329), .A2(new_n206), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n256), .A2(G33), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n261), .A2(new_n352), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n206), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT83), .B1(new_n275), .B2(G77), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n275), .A2(KEYINPUT83), .A3(G77), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n210), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  XNOR2_X1  g0296(.A(G97), .B(G107), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n494), .B(new_n495), .C1(new_n499), .C2(new_n228), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n400), .B2(G107), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n488), .B(new_n492), .C1(new_n501), .C2(new_n352), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n292), .A2(G244), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n355), .B2(new_n289), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT84), .B1(new_n505), .B2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT4), .ZN(new_n508));
  NOR2_X1   g0308(.A1(KEYINPUT3), .A2(G33), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(G33), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n507), .B(new_n508), .C1(new_n511), .C2(new_n504), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n504), .A2(new_n508), .B1(new_n205), .B2(new_n292), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n513), .A2(new_n291), .B1(G33), .B2(G283), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n506), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n296), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n364), .A3(KEYINPUT5), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT5), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(KEYINPUT85), .B2(G41), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n365), .A2(G1), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G274), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n522), .A2(new_n301), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G257), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n516), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G200), .ZN(new_n528));
  INV_X1    g0328(.A(new_n526), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n515), .B2(new_n296), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G190), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n503), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n373), .A2(new_n228), .A3(G68), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n204), .A2(new_n206), .A3(new_n210), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n535), .A2(new_n264), .A3(new_n206), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n534), .B1(new_n536), .B2(G20), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n475), .B2(new_n206), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n533), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n265), .ZN(new_n540));
  INV_X1    g0340(.A(new_n490), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n476), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n261), .A2(new_n476), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n301), .B1(G250), .B2(new_n521), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n365), .A2(G1), .A3(G274), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G116), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n264), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G238), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n355), .A2(new_n289), .B1(new_n552), .B2(new_n292), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n217), .A2(G1698), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n484), .B(new_n549), .C1(new_n555), .C2(new_n301), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n292), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n373), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n551), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n301), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n310), .B1(new_n560), .B2(new_n548), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n545), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(G200), .B1(new_n560), .B2(new_n548), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n543), .B1(new_n539), .B2(new_n265), .ZN(new_n564));
  OAI211_X1 g0364(.A(G190), .B(new_n549), .C1(new_n555), .C2(new_n301), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT86), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n490), .B2(new_n204), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n266), .A2(KEYINPUT86), .A3(G87), .A4(new_n489), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n563), .A2(new_n564), .A3(new_n565), .A4(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n516), .A2(new_n484), .A3(new_n526), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n502), .B(new_n572), .C1(G169), .C2(new_n530), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n522), .A2(G270), .A3(new_n301), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT87), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n524), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G257), .A2(G1698), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n292), .A2(G264), .ZN(new_n579));
  AOI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n355), .C2(new_n289), .ZN(new_n580));
  INV_X1    g0380(.A(G303), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n291), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n296), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n261), .A2(G116), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n490), .A2(new_n550), .ZN(new_n587));
  AOI21_X1  g0387(.A(G20), .B1(G33), .B2(G283), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G33), .B2(new_n206), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n550), .A2(G20), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n265), .A2(KEYINPUT88), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT88), .B1(new_n265), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT20), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(KEYINPUT20), .B(new_n589), .C1(new_n592), .C2(new_n593), .ZN(new_n597));
  AOI211_X1 g0397(.A(new_n586), .B(new_n587), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n585), .B(new_n598), .C1(new_n383), .C2(new_n584), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n532), .A2(new_n571), .A3(new_n573), .A4(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n579), .B1(new_n355), .B2(new_n289), .ZN(new_n601));
  INV_X1    g0401(.A(new_n578), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n582), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n577), .B1(new_n603), .B2(new_n301), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n574), .B(KEYINPUT87), .ZN(new_n605));
  OAI21_X1  g0405(.A(G169), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n598), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n579), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n373), .A2(new_n602), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n582), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n524), .B1(new_n612), .B2(new_n296), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n310), .B1(new_n613), .B2(new_n576), .ZN(new_n614));
  INV_X1    g0414(.A(new_n587), .ZN(new_n615));
  INV_X1    g0415(.A(new_n586), .ZN(new_n616));
  INV_X1    g0416(.A(new_n593), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n591), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT20), .B1(new_n618), .B2(new_n589), .ZN(new_n619));
  INV_X1    g0419(.A(new_n597), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n615), .B(new_n616), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT21), .B1(new_n614), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n608), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT23), .B1(new_n228), .B2(G107), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT23), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n210), .A3(G20), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n228), .A2(G33), .A3(G116), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT89), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n624), .A2(new_n626), .A3(new_n627), .A4(KEYINPUT89), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n204), .A2(G20), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n373), .A2(KEYINPUT22), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n291), .A2(new_n633), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT22), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n632), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT24), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n630), .A2(new_n631), .B1(new_n635), .B2(new_n636), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT24), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n634), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n352), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n490), .A2(new_n210), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT25), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n261), .B2(G107), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(KEYINPUT90), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n205), .A2(new_n292), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n292), .A2(G257), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n373), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G294), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n264), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n656), .A2(new_n296), .B1(G264), .B2(new_n525), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT91), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n657), .A2(new_n658), .A3(new_n383), .A4(new_n577), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n525), .A2(G264), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n650), .B1(new_n355), .B2(new_n289), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n654), .B1(new_n661), .B2(new_n649), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n577), .B(new_n660), .C1(new_n662), .C2(new_n301), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT91), .B1(new_n663), .B2(G190), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n362), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n659), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n329), .A2(KEYINPUT25), .A3(new_n210), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(KEYINPUT90), .A3(new_n646), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n648), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n584), .A2(new_n484), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n621), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n641), .A2(new_n632), .A3(new_n637), .A4(new_n634), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n641), .B1(new_n640), .B2(new_n634), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n265), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n644), .ZN(new_n675));
  INV_X1    g0475(.A(new_n647), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n674), .A2(new_n668), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n663), .A2(G179), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n310), .B2(new_n663), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n623), .A2(new_n669), .A3(new_n671), .A4(new_n680), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n487), .A2(new_n600), .A3(new_n681), .ZN(G372));
  NAND2_X1  g0482(.A1(new_n456), .A2(new_n486), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n460), .A3(new_n388), .A4(new_n412), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT92), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n392), .B2(new_n406), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT18), .B1(new_n361), .B2(new_n391), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n404), .A2(new_n393), .A3(new_n405), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(KEYINPUT92), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n322), .A2(new_n326), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(new_n312), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n573), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n570), .A2(KEYINPUT26), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n532), .A2(new_n570), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n677), .A2(new_n679), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n607), .B1(new_n598), .B2(new_n606), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n614), .A2(KEYINPUT21), .A3(new_n621), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n671), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n669), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n699), .B1(new_n704), .B2(new_n573), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n698), .B1(new_n705), .B2(KEYINPUT26), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n562), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n695), .B1(new_n487), .B2(new_n708), .ZN(G369));
  NAND2_X1  g0509(.A1(new_n228), .A2(G13), .ZN(new_n710));
  OR3_X1    g0510(.A1(new_n710), .A2(KEYINPUT27), .A3(G1), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT27), .B1(new_n710), .B2(G1), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G343), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n677), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n700), .B1(new_n669), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n680), .A2(new_n715), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n715), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n703), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n621), .A2(new_n715), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n703), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n703), .A2(new_n724), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n599), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G330), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n722), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n718), .B1(new_n719), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(G399));
  NOR2_X1   g0533(.A1(new_n225), .A2(G41), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n534), .A2(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G1), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n235), .B2(new_n735), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n400), .A2(G107), .ZN(new_n740));
  INV_X1    g0540(.A(new_n500), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n491), .B1(new_n742), .B2(new_n265), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n743), .A2(new_n488), .B1(new_n527), .B2(new_n310), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT93), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n697), .A3(new_n745), .A4(new_n572), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT26), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n562), .A2(new_n570), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n573), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n570), .A2(KEYINPUT26), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT93), .B1(new_n573), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n746), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n752), .A2(KEYINPUT94), .A3(new_n562), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT94), .B1(new_n752), .B2(new_n562), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n532), .A2(new_n571), .A3(new_n573), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n704), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(KEYINPUT29), .B1(new_n757), .B2(new_n715), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT29), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n707), .A2(new_n759), .A3(new_n721), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n560), .A2(new_n548), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n670), .A2(new_n530), .A3(new_n762), .A4(new_n657), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT30), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n527), .A2(new_n484), .A3(new_n584), .A4(new_n663), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(new_n762), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT31), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(new_n770), .A3(new_n715), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n681), .A2(new_n600), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(new_n773), .B2(new_n721), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n769), .A2(new_n715), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n772), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G330), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n761), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n739), .B1(new_n779), .B2(G1), .ZN(G364));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n727), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n291), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n228), .A2(new_n383), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n362), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n785), .B1(new_n788), .B2(new_n581), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G179), .A2(G200), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n228), .B1(new_n790), .B2(G190), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT98), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(KEYINPUT98), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n789), .B1(new_n795), .B2(G294), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n228), .A2(G190), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n787), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n484), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n786), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n797), .A2(new_n790), .ZN(new_n804));
  INV_X1    g0604(.A(G329), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n484), .A2(new_n362), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n797), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT33), .B(G317), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n800), .B(new_n806), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n807), .A2(new_n786), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G326), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n797), .A2(new_n801), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G311), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n796), .A2(new_n811), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n788), .A2(new_n204), .B1(new_n815), .B2(new_n216), .ZN(new_n819));
  INV_X1    g0619(.A(G159), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n804), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT97), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(KEYINPUT32), .ZN(new_n823));
  INV_X1    g0623(.A(new_n798), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n819), .B(new_n823), .C1(G107), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n802), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G58), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n794), .A2(new_n206), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n785), .B(new_n828), .C1(G50), .C2(new_n813), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n822), .A2(KEYINPUT32), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n825), .A2(new_n827), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n808), .A2(new_n333), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n818), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n227), .B1(G20), .B2(new_n310), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n710), .B(KEYINPUT95), .Z(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G45), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G1), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n735), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT96), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n783), .A2(new_n834), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n785), .A2(new_n225), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G355), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n251), .A2(new_n365), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n373), .A2(new_n225), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n235), .B2(G45), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n845), .B1(G116), .B2(new_n224), .C1(new_n846), .C2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n842), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n784), .A2(new_n835), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT99), .ZN(new_n852));
  INV_X1    g0652(.A(new_n729), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n842), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n728), .B2(new_n727), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(G396));
  AOI21_X1  g0657(.A(new_n715), .B1(new_n706), .B2(new_n562), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n486), .A2(new_n715), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n481), .A2(new_n715), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n483), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n859), .B1(new_n861), .B2(new_n486), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n859), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n471), .A2(new_n482), .B1(new_n481), .B2(new_n715), .ZN(new_n865));
  INV_X1    g0665(.A(new_n486), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n715), .B(new_n867), .C1(new_n706), .C2(new_n562), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(new_n777), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n842), .ZN(new_n871));
  INV_X1    g0671(.A(new_n834), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n798), .A2(new_n204), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n873), .B(new_n828), .C1(G294), .C2(new_n826), .ZN(new_n874));
  INV_X1    g0674(.A(G311), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n815), .A2(new_n550), .B1(new_n804), .B2(new_n875), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n291), .B(new_n876), .C1(G283), .C2(new_n809), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n878), .B1(new_n210), .B2(new_n788), .C1(new_n581), .C2(new_n812), .ZN(new_n879));
  INV_X1    g0679(.A(G132), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n804), .A2(new_n880), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n373), .B1(new_n333), .B2(new_n798), .C1(new_n794), .C2(new_n219), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT34), .ZN(new_n883));
  AOI22_X1  g0683(.A1(G143), .A2(new_n826), .B1(new_n816), .B2(G159), .ZN(new_n884));
  INV_X1    g0684(.A(G137), .ZN(new_n885));
  INV_X1    g0685(.A(G150), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n884), .B1(new_n885), .B2(new_n812), .C1(new_n886), .C2(new_n808), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n887), .ZN(new_n888));
  OAI221_X1 g0688(.A(new_n888), .B1(new_n883), .B2(new_n887), .C1(new_n214), .C2(new_n788), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n872), .B1(new_n879), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n834), .A2(new_n781), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT100), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n842), .B(new_n890), .C1(new_n216), .C2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n862), .B2(new_n782), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n871), .A2(new_n894), .ZN(G384));
  NAND2_X1  g0695(.A1(new_n410), .A2(new_n411), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n686), .B2(new_n689), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n361), .A2(new_n713), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT107), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n404), .A2(new_n405), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(new_n685), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n404), .A2(new_n409), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(new_n898), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n901), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n902), .A2(KEYINPUT105), .ZN(new_n908));
  INV_X1    g0708(.A(new_n901), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n902), .A2(KEYINPUT105), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n908), .A2(new_n905), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n896), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n687), .A2(KEYINPUT92), .A3(new_n688), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT92), .B1(new_n687), .B2(new_n688), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT107), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(new_n898), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n900), .A2(new_n912), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n359), .A2(KEYINPUT16), .ZN(new_n922));
  OR3_X1    g0722(.A1(new_n922), .A2(KEYINPUT103), .A3(new_n352), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT103), .B1(new_n922), .B2(new_n352), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n397), .A3(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n925), .A2(new_n403), .B1(new_n391), .B2(new_n713), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT37), .B1(new_n926), .B2(new_n904), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n911), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n713), .B1(new_n925), .B2(new_n403), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n413), .A2(KEYINPUT104), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT104), .B1(new_n413), .B2(new_n929), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT38), .B(new_n928), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n921), .A2(new_n932), .ZN(new_n933));
  AND4_X1   g0733(.A1(new_n573), .A2(new_n532), .A3(new_n571), .A4(new_n599), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n700), .A2(new_n703), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(new_n669), .A4(new_n721), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(KEYINPUT31), .A3(new_n775), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n771), .A3(new_n862), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n455), .A2(new_n453), .A3(new_n715), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n456), .A2(new_n460), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n431), .A2(new_n453), .A3(new_n455), .A4(new_n715), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT102), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(new_n940), .B2(new_n941), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n933), .A2(KEYINPUT40), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n920), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n932), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT40), .B1(new_n951), .B2(new_n946), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n948), .A2(new_n952), .A3(new_n487), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n951), .A2(new_n946), .ZN(new_n954));
  OAI211_X1 g0754(.A(G330), .B(new_n947), .C1(new_n954), .C2(KEYINPUT40), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n777), .A2(new_n487), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n776), .A2(new_n953), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n950), .A2(KEYINPUT39), .A3(new_n932), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n456), .A2(new_n715), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT39), .B1(new_n921), .B2(new_n932), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n950), .A2(new_n932), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n940), .A2(new_n941), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT102), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n940), .A2(new_n942), .A3(new_n941), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n868), .B2(new_n859), .ZN(new_n969));
  INV_X1    g0769(.A(new_n713), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n964), .A2(new_n969), .B1(new_n690), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n963), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n958), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n487), .B1(new_n758), .B2(new_n760), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n694), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n973), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n256), .B2(new_n836), .ZN(new_n977));
  OAI21_X1  g0777(.A(G77), .B1(new_n219), .B2(new_n333), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n235), .A2(new_n978), .B1(G50), .B2(new_n333), .ZN(new_n979));
  INV_X1    g0779(.A(G13), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(G1), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT35), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n230), .B1(new_n499), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n983), .B(G116), .C1(new_n982), .C2(new_n499), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT101), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT36), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n977), .A2(new_n981), .A3(new_n986), .ZN(G367));
  AOI21_X1  g0787(.A(new_n721), .B1(new_n564), .B2(new_n569), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n562), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n571), .B2(new_n988), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT108), .Z(new_n991));
  INV_X1    g0791(.A(KEYINPUT43), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n532), .B(new_n573), .C1(new_n503), .C2(new_n721), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n696), .A2(new_n715), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT109), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT109), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n719), .A2(new_n731), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT42), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n999), .A2(new_n700), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n715), .B1(new_n1004), .B2(new_n573), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n993), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n991), .A2(new_n992), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n730), .A2(new_n1000), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1003), .A2(new_n992), .A3(new_n991), .A4(new_n1006), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n730), .B2(new_n1000), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n734), .B(KEYINPUT41), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n999), .A2(new_n732), .A3(KEYINPUT44), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT44), .B1(new_n999), .B2(new_n732), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n999), .A2(KEYINPUT45), .A3(new_n732), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT45), .B1(new_n999), .B2(new_n732), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(new_n730), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n730), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1019), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n853), .A2(new_n720), .A3(new_n722), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1028), .A2(new_n730), .A3(new_n1001), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1029), .A2(new_n777), .A3(new_n758), .A4(new_n760), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1030), .A2(KEYINPUT110), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(KEYINPUT110), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1027), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1016), .B1(new_n1033), .B2(new_n779), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1012), .B(new_n1014), .C1(new_n1034), .C2(new_n838), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n842), .B1(new_n991), .B2(new_n783), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n847), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n843), .B1(new_n224), .B2(new_n477), .C1(new_n247), .C2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n291), .B1(new_n788), .B2(new_n219), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G159), .A2(new_n809), .B1(new_n824), .B2(G77), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n214), .B2(new_n815), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n813), .A2(G143), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n886), .B2(new_n802), .C1(new_n794), .C2(new_n333), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1039), .B(new_n1041), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n885), .B2(new_n804), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT112), .Z(new_n1048));
  INV_X1    g0848(.A(G317), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n798), .A2(new_n206), .B1(new_n804), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n788), .A2(new_n550), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1051), .A2(KEYINPUT46), .B1(new_n581), .B2(new_n802), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1051), .A2(KEYINPUT46), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n808), .A2(new_n653), .ZN(new_n1054));
  OR4_X1    g0854(.A1(new_n373), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1050), .B(new_n1055), .C1(G311), .C2(new_n813), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n210), .B2(new_n794), .C1(new_n799), .C2(new_n815), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1048), .A2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT47), .Z(new_n1059));
  OAI211_X1 g0859(.A(new_n1036), .B(new_n1038), .C1(new_n1059), .C2(new_n872), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1035), .A2(new_n1060), .ZN(G387));
  AOI21_X1  g0861(.A(new_n1037), .B1(new_n243), .B2(G45), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n736), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1062), .B1(new_n1063), .B2(new_n844), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n270), .A2(new_n214), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT50), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n333), .A2(new_n216), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1066), .A2(G45), .A3(new_n1067), .A4(new_n1063), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1064), .A2(new_n1068), .B1(G107), .B2(new_n224), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n842), .B1(new_n1069), .B2(new_n843), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n783), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1070), .B1(new_n719), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n795), .A2(new_n476), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n214), .B2(new_n802), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT113), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n804), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G68), .A2(new_n816), .B1(new_n1076), .B2(G150), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n216), .B2(new_n788), .C1(new_n478), .C2(new_n808), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n511), .B(new_n1078), .C1(G97), .C2(new_n824), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1075), .B(new_n1079), .C1(new_n820), .C2(new_n812), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n788), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n795), .A2(G283), .B1(G294), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n813), .A2(G322), .B1(new_n809), .B2(G311), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n581), .B2(new_n815), .C1(new_n1049), .C2(new_n802), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT114), .Z(new_n1085));
  INV_X1    g0885(.A(KEYINPUT48), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1082), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT115), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT49), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1076), .A2(G326), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n824), .A2(G116), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1090), .A2(new_n511), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1089), .A2(KEYINPUT49), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1080), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1072), .B1(new_n1095), .B2(new_n834), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n838), .B2(new_n1029), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n779), .B2(new_n1029), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1099), .B2(new_n735), .ZN(G393));
  OAI21_X1  g0900(.A(new_n843), .B1(new_n206), .B2(new_n224), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n254), .B2(new_n847), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n794), .A2(new_n216), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G150), .A2(new_n813), .B1(new_n826), .B2(G159), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1103), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n816), .A2(new_n270), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1104), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n873), .B1(new_n1109), .B2(new_n1105), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n214), .A2(new_n808), .B1(new_n788), .B2(new_n333), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n511), .B(new_n1111), .C1(G143), .C2(new_n1076), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n812), .A2(new_n1049), .B1(new_n802), .B2(new_n875), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT52), .Z(new_n1115));
  NOR2_X1   g0915(.A1(new_n788), .A2(new_n799), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n210), .A2(new_n798), .B1(new_n815), .B2(new_n653), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1115), .A2(new_n291), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n550), .B2(new_n794), .C1(new_n581), .C2(new_n808), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n804), .A2(new_n803), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1113), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n842), .B(new_n1102), .C1(new_n1121), .C2(new_n834), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n999), .B2(new_n1071), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n839), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n735), .B1(new_n1124), .B2(new_n1098), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n1033), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(G390));
  INV_X1    g0928(.A(KEYINPUT39), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n933), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n950), .A2(KEYINPUT39), .A3(new_n932), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1130), .A2(new_n1131), .B1(new_n969), .B2(new_n961), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n933), .A2(new_n961), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n861), .A2(new_n486), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n752), .A2(new_n562), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT94), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n752), .A2(KEYINPUT94), .A3(new_n562), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n721), .B(new_n1134), .C1(new_n1139), .C2(new_n756), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n945), .B1(new_n1140), .B2(new_n864), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1133), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n776), .A2(G330), .A3(new_n968), .A4(new_n862), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1132), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n707), .A2(new_n721), .A3(new_n862), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n945), .B1(new_n1146), .B2(new_n864), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n959), .A2(new_n962), .B1(new_n960), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1140), .A2(new_n864), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n961), .B(new_n933), .C1(new_n1149), .C2(new_n945), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1143), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1145), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n937), .A2(G330), .A3(new_n771), .A4(new_n862), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n945), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1143), .A2(new_n864), .A3(new_n1154), .A4(new_n1140), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n946), .A2(G330), .B1(new_n945), .B2(new_n1153), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n859), .B1(new_n858), .B2(new_n862), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n974), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n695), .A3(new_n957), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT117), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n974), .A2(new_n694), .A3(new_n956), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT117), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1158), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1152), .A2(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1163), .A2(new_n1158), .A3(new_n1164), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1164), .B1(new_n1163), .B2(new_n1158), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1144), .B1(new_n1132), .B2(new_n1142), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1148), .A2(new_n1150), .A3(new_n1143), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1167), .A2(new_n1174), .A3(new_n734), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n781), .B1(new_n959), .B2(new_n962), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n892), .A2(new_n478), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n291), .B1(new_n813), .B2(G283), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n206), .B2(new_n815), .C1(new_n210), .C2(new_n808), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1103), .B(new_n1179), .C1(G116), .C2(new_n826), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G87), .A2(new_n1081), .B1(new_n824), .B2(G68), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n653), .C2(new_n804), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n802), .A2(new_n880), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n785), .B1(new_n809), .B2(G137), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT54), .B(G143), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1185), .B1(new_n214), .B2(new_n798), .C1(new_n815), .C2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1184), .B(new_n1187), .C1(G128), .C2(new_n813), .ZN(new_n1188));
  INV_X1    g0988(.A(G125), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1188), .B1(new_n1189), .B2(new_n804), .C1(new_n820), .C2(new_n794), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n788), .A2(new_n886), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n842), .B(new_n1177), .C1(new_n1194), .C2(new_n834), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1152), .A2(new_n838), .B1(new_n1176), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1175), .A2(new_n1196), .ZN(G378));
  INV_X1    g0997(.A(KEYINPUT57), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1161), .B1(new_n1152), .B2(new_n1166), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1130), .A2(new_n960), .A3(new_n1131), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n690), .A2(new_n970), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1147), .B2(new_n951), .ZN(new_n1202));
  XOR2_X1   g1002(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n327), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n327), .A2(new_n1204), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n315), .A2(new_n713), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OR3_X1    g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1200), .A2(new_n1202), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n955), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1211), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n963), .B2(new_n971), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n948), .A2(new_n952), .A3(new_n728), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1200), .A2(new_n1202), .A3(new_n1211), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1214), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1198), .B1(new_n1199), .B2(new_n1220), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1212), .A2(new_n1213), .A3(new_n955), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1217), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1163), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(KEYINPUT57), .A3(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1221), .A2(new_n1226), .A3(new_n734), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n794), .A2(new_n886), .B1(new_n885), .B2(new_n815), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n812), .A2(new_n1189), .B1(new_n808), .B2(new_n880), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n826), .A2(G128), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n788), .C2(new_n1186), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n824), .A2(G159), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G41), .B1(new_n1076), .B2(G124), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1233), .A2(new_n264), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1237));
  AOI21_X1  g1037(.A(G41), .B1(new_n510), .B2(G33), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n1236), .A2(new_n1237), .B1(G50), .B2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n788), .A2(new_n216), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n511), .B(new_n364), .C1(new_n206), .C2(new_n808), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(G283), .C2(new_n1076), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n794), .A2(new_n333), .B1(new_n477), .B2(new_n815), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n812), .A2(new_n550), .B1(new_n798), .B2(new_n219), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1242), .B(new_n1245), .C1(new_n210), .C2(new_n802), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT58), .Z(new_n1247));
  OAI21_X1  g1047(.A(new_n834), .B1(new_n1239), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n842), .B1(new_n214), .B2(new_n891), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1211), .B2(new_n781), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1224), .B2(new_n838), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1227), .A2(new_n1252), .ZN(G375));
  NAND2_X1  g1053(.A1(new_n945), .A2(new_n781), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n892), .A2(new_n333), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n815), .A2(new_n886), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n812), .A2(new_n880), .B1(new_n808), .B2(new_n1186), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G137), .B2(new_n826), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT121), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n788), .A2(new_n820), .B1(new_n798), .B2(new_n219), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G128), .B2(new_n1076), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n373), .A3(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1256), .B(new_n1262), .C1(G50), .C2(new_n795), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1073), .B1(new_n206), .B2(new_n788), .C1(new_n799), .C2(new_n802), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n813), .A2(G294), .B1(new_n816), .B2(G107), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n550), .B2(new_n808), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT120), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1266), .A2(new_n1267), .B1(G77), .B2(new_n824), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1268), .B(new_n785), .C1(new_n1267), .C2(new_n1266), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1264), .B(new_n1269), .C1(G303), .C2(new_n1076), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n834), .B1(new_n1263), .B2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1254), .A2(new_n841), .A3(new_n1255), .A4(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1159), .B2(new_n839), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1015), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1166), .B2(new_n1276), .ZN(G381));
  NOR2_X1   g1077(.A1(G375), .A2(G378), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(G381), .A2(G384), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1035), .A2(new_n1060), .A3(new_n1127), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1280), .A2(G396), .A3(G393), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1278), .A2(new_n1279), .A3(new_n1281), .ZN(G407));
  NAND2_X1  g1082(.A1(new_n714), .A2(G213), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1278), .A2(KEYINPUT122), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G407), .A2(new_n1285), .A3(G213), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT122), .B1(new_n1278), .B2(new_n1284), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1286), .A2(new_n1287), .ZN(G409));
  NAND2_X1  g1088(.A1(G375), .A2(G378), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n839), .A2(KEYINPUT123), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1199), .B2(new_n1016), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1251), .B1(new_n1291), .B2(new_n1224), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1220), .A2(KEYINPUT123), .A3(new_n838), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1293), .A2(new_n1175), .A3(new_n1196), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1284), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1289), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1284), .A2(G2897), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1275), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1275), .A2(KEYINPUT124), .A3(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT124), .B1(new_n1163), .B2(new_n1158), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n735), .B1(new_n1302), .B2(KEYINPUT60), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1299), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1299), .A2(new_n1303), .A3(KEYINPUT125), .A4(new_n1301), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(G384), .B1(new_n1308), .B2(new_n1274), .ZN(new_n1309));
  INV_X1    g1109(.A(G384), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n1310), .B(new_n1273), .C1(new_n1306), .C2(new_n1307), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1284), .A2(KEYINPUT126), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1298), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1313), .ZN(new_n1315));
  NOR4_X1   g1115(.A1(new_n1309), .A2(new_n1311), .A3(new_n1297), .A4(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1296), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1289), .A2(new_n1312), .A3(new_n1295), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT61), .B1(new_n1318), .B2(KEYINPUT62), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1289), .A2(new_n1312), .A3(new_n1295), .A4(new_n1320), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1317), .A2(new_n1319), .A3(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(G393), .B(new_n856), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1280), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1127), .B1(new_n1035), .B2(new_n1060), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1325), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G387), .A2(G390), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT127), .B1(new_n1329), .B2(new_n1280), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1324), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1327), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1323), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1318), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1335), .B1(new_n1317), .B2(KEYINPUT63), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT61), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1289), .A2(new_n1312), .A3(new_n1295), .A4(KEYINPUT63), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1334), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  OAI22_X1  g1139(.A1(new_n1322), .A2(new_n1334), .B1(new_n1336), .B2(new_n1339), .ZN(G405));
  XNOR2_X1  g1140(.A(G375), .B(G378), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1341), .B(new_n1312), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1334), .ZN(new_n1343));
  OR2_X1    g1143(.A1(new_n1341), .A2(new_n1312), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1341), .A2(new_n1312), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1344), .A2(new_n1331), .A3(new_n1333), .A4(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1343), .A2(new_n1346), .ZN(G402));
endmodule


