//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n207), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n213), .B(new_n227), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n222), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G97), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n228), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT6), .ZN(new_n250));
  NOR3_X1   g0050(.A1(new_n250), .A2(new_n223), .A3(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G97), .B(G107), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n251), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n207), .A2(new_n255), .A3(KEYINPUT66), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT66), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G20), .B2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n253), .A2(new_n207), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G107), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT7), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n255), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n263), .B1(new_n267), .B2(G20), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n262), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n249), .B1(new_n261), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n223), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n249), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G1), .B2(new_n255), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G97), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n274), .A2(new_n277), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n206), .A2(G45), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT5), .A2(G41), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT5), .A2(G41), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  INV_X1    g0088(.A(new_n228), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G1), .ZN(new_n294));
  AND2_X1   g0094(.A1(KEYINPUT5), .A2(G41), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(new_n284), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(new_n290), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(G257), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT4), .ZN(new_n300));
  OR2_X1    g0100(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n301), .B(new_n302), .C1(new_n269), .C2(new_n270), .ZN(new_n303));
  INV_X1    g0103(.A(G244), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G1698), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n265), .B2(new_n266), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT65), .B(G1698), .Z(new_n309));
  NAND4_X1  g0109(.A1(new_n309), .A2(KEYINPUT4), .A3(G244), .A4(new_n267), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n299), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n282), .B(new_n315), .C1(G169), .C2(new_n313), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(G190), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n277), .B1(new_n279), .B2(new_n223), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n254), .B1(new_n256), .B2(new_n258), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n252), .A2(new_n250), .ZN(new_n320));
  INV_X1    g0120(.A(new_n251), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n319), .B1(new_n322), .B2(G20), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n267), .A2(new_n263), .A3(G20), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT7), .B1(new_n271), .B2(new_n207), .ZN(new_n325));
  OAI21_X1  g0125(.A(G107), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n318), .B1(new_n327), .B2(new_n249), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n317), .B(new_n328), .C1(new_n329), .C2(new_n313), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT76), .ZN(new_n333));
  OAI211_X1 g0133(.A(G244), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n267), .A2(KEYINPUT75), .A3(G244), .A4(G1698), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G116), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n303), .A2(new_n216), .B1(new_n255), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n333), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n255), .A2(new_n339), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT65), .B(G1698), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n271), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n344), .B2(G238), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n336), .A2(new_n337), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(KEYINPUT76), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n297), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n312), .A2(new_n218), .A3(new_n294), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n350), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n351), .A2(new_n352), .B1(new_n291), .B2(new_n294), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n332), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n345), .A2(KEYINPUT76), .A3(new_n346), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT76), .B1(new_n345), .B2(new_n346), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n312), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(new_n314), .A3(new_n353), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n255), .A2(G20), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT19), .B1(new_n360), .B2(G97), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n271), .A2(G20), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(G68), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G97), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT69), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(G20), .B1(new_n366), .B2(KEYINPUT19), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT77), .B(G87), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(new_n223), .A3(new_n262), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n363), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n249), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT68), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n275), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n206), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n372), .B(new_n379), .C1(new_n378), .C2(new_n279), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n355), .A2(new_n359), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(G200), .B1(new_n348), .B2(new_n354), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n358), .A2(G190), .A3(new_n353), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n280), .A2(G87), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n372), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n331), .A2(new_n381), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(G20), .B1(G33), .B2(G283), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G33), .B2(new_n223), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n339), .A2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n249), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT20), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n391), .B(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n249), .B1(new_n374), .B2(new_n375), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n339), .B1(new_n206), .B2(G33), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n377), .A2(new_n339), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n332), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT78), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n224), .B1(new_n265), .B2(new_n266), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n309), .B1(G303), .B2(new_n271), .ZN(new_n400));
  OAI211_X1 g0200(.A(G264), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n297), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n296), .A2(new_n297), .ZN(new_n403));
  INV_X1    g0203(.A(G270), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n292), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n398), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n265), .A2(G303), .A3(new_n266), .ZN(new_n407));
  OAI21_X1  g0207(.A(G257), .B1(new_n269), .B2(new_n270), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n401), .B(new_n407), .C1(new_n408), .C2(new_n343), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n312), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT5), .B(G41), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(new_n294), .B1(new_n289), .B2(new_n290), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(G270), .B1(new_n291), .B2(new_n287), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(new_n413), .A3(KEYINPUT78), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n397), .A2(new_n406), .A3(KEYINPUT21), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n393), .A2(new_n396), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n416), .A2(G179), .A3(new_n410), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n410), .A2(new_n413), .A3(KEYINPUT78), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT78), .B1(new_n410), .B2(new_n413), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT21), .B1(new_n421), .B2(new_n397), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n296), .A2(G264), .A3(new_n297), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT80), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT80), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n296), .A2(new_n426), .A3(G264), .A4(new_n297), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G294), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(new_n430), .C1(new_n303), .C2(new_n218), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n312), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n428), .A2(new_n292), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(KEYINPUT81), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT81), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n428), .A2(new_n292), .A3(new_n432), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(new_n329), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(G190), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n279), .A2(new_n262), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n276), .A2(new_n262), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT25), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n207), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT22), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT22), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n267), .A2(new_n448), .A3(new_n207), .A4(G87), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT23), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n207), .B2(G107), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n262), .A2(KEYINPUT23), .A3(G20), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n452), .A2(new_n453), .B1(new_n342), .B2(new_n207), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT79), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n450), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(KEYINPUT24), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n249), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n457), .B1(new_n450), .B2(new_n454), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT24), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n445), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n440), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n421), .A2(G200), .ZN(new_n466));
  INV_X1    g0266(.A(new_n416), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n466), .B(new_n467), .C1(new_n434), .C2(new_n421), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n459), .A2(new_n463), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n444), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n437), .A2(new_n332), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n437), .A2(G179), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n423), .A2(new_n465), .A3(new_n468), .A4(new_n474), .ZN(new_n475));
  XOR2_X1   g0275(.A(KEYINPUT8), .B(G58), .Z(new_n476));
  AOI22_X1  g0276(.A1(new_n476), .A2(new_n360), .B1(G20), .B2(new_n203), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n259), .A2(G150), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n460), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n278), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n206), .A2(G20), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G50), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n480), .A2(new_n482), .B1(G50), .B2(new_n275), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n484), .A2(KEYINPUT9), .ZN(new_n485));
  INV_X1    g0285(.A(G223), .ZN(new_n486));
  INV_X1    g0286(.A(G222), .ZN(new_n487));
  OAI221_X1 g0287(.A(new_n267), .B1(new_n486), .B2(new_n306), .C1(new_n343), .C2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(new_n312), .C1(G77), .C2(new_n267), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n312), .A2(new_n288), .A3(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n297), .A2(new_n490), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(G226), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(G190), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n484), .A2(KEYINPUT9), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n489), .A2(new_n493), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n485), .A2(new_n494), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT10), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n484), .B1(new_n496), .B2(new_n332), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(G179), .B2(new_n496), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI221_X1 g0302(.A(new_n267), .B1(new_n216), .B2(new_n306), .C1(new_n343), .C2(new_n222), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n312), .C1(G107), .C2(new_n267), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n491), .B1(G244), .B2(new_n492), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G179), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n332), .B2(new_n506), .ZN(new_n508));
  INV_X1    g0308(.A(new_n378), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n360), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT67), .ZN(new_n511));
  INV_X1    g0311(.A(new_n476), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n512), .A2(new_n260), .B1(new_n207), .B2(new_n254), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n249), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n254), .B1(new_n206), .B2(G20), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n377), .A2(new_n254), .B1(new_n394), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n506), .A2(G200), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n434), .B2(new_n506), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n502), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n309), .A2(G226), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G232), .A2(G1698), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n271), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n312), .B1(new_n525), .B2(new_n366), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n491), .B1(G238), .B2(new_n492), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT13), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(KEYINPUT70), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT70), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n526), .A2(new_n531), .A3(KEYINPUT13), .A4(new_n527), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G190), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT71), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n529), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n526), .A2(KEYINPUT13), .A3(new_n527), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(G200), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n259), .A2(G50), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n360), .A2(G77), .B1(G20), .B2(new_n215), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n460), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n541), .A2(KEYINPUT11), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n394), .A2(G68), .A3(new_n481), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(KEYINPUT11), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT12), .B1(new_n376), .B2(G68), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n207), .A2(KEYINPUT12), .A3(G68), .ZN(new_n546));
  INV_X1    g0346(.A(G13), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(G1), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n534), .A2(new_n535), .A3(new_n538), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n538), .A2(new_n552), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n434), .B1(new_n530), .B2(new_n532), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT71), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n476), .A2(new_n481), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n278), .B1(new_n276), .B2(new_n512), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n215), .B1(new_n268), .B2(new_n272), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G58), .B(G68), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n259), .A2(G159), .B1(new_n562), .B2(G20), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n460), .B1(new_n565), .B2(KEYINPUT16), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT16), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n561), .B2(new_n564), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n560), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G226), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G87), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n570), .B(new_n571), .C1(new_n303), .C2(new_n486), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n312), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n491), .B1(G232), .B2(new_n492), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n332), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n575), .B1(G179), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT18), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n573), .A2(new_n574), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G169), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n314), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g0381(.A(G68), .B1(new_n324), .B2(new_n325), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(KEYINPUT16), .A3(new_n563), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n568), .A2(new_n583), .A3(new_n249), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n559), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT18), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n579), .A2(G200), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n573), .A2(new_n574), .A3(G190), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n584), .A2(new_n559), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT17), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n329), .B1(new_n573), .B2(new_n574), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(G190), .B2(new_n576), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n594), .A2(KEYINPUT17), .A3(new_n584), .A4(new_n559), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n578), .A2(new_n587), .A3(new_n592), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n536), .A2(G169), .A3(new_n537), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT72), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT14), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n533), .A2(G179), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(KEYINPUT14), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n536), .A2(G169), .A3(new_n537), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n596), .B1(new_n551), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n522), .A2(new_n557), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT73), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n522), .A2(KEYINPUT73), .A3(new_n557), .A4(new_n604), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n387), .B(new_n475), .C1(new_n607), .C2(new_n608), .ZN(G372));
  NAND2_X1  g0409(.A1(new_n592), .A2(new_n595), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(new_n551), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n534), .A2(new_n538), .A3(new_n552), .ZN(new_n612));
  INV_X1    g0412(.A(new_n518), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n610), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n578), .A2(new_n587), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n499), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n501), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n607), .A2(new_n608), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n381), .A2(new_n386), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT26), .B1(new_n621), .B2(new_n316), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT82), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n460), .B1(new_n323), .B2(new_n326), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n313), .A2(G169), .B1(new_n624), .B2(new_n318), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n313), .A2(new_n314), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n313), .A2(G169), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(KEYINPUT82), .A3(new_n315), .A4(new_n282), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n381), .A4(new_n386), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n622), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n406), .A2(new_n416), .A3(G169), .A4(new_n414), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n417), .A3(new_n415), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n437), .A2(new_n332), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(G179), .B2(new_n437), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n464), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n465), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n381), .B1(new_n387), .B2(new_n641), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n619), .B1(new_n620), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g0444(.A(new_n644), .B(KEYINPUT83), .Z(G369));
  AND2_X1   g0445(.A1(new_n423), .A2(new_n468), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n548), .A2(new_n207), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n416), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n423), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n470), .A2(new_n652), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n465), .A2(new_n474), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n640), .A2(new_n652), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT84), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT84), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n659), .A2(new_n663), .A3(new_n660), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n423), .A2(new_n652), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n662), .B2(new_n664), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n474), .A2(new_n652), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n210), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n206), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n369), .A2(G116), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n675), .A2(new_n676), .B1(new_n231), .B2(new_n674), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT28), .Z(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  INV_X1    g0479(.A(new_n652), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n643), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n627), .A2(new_n629), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT26), .B1(new_n621), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n316), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n381), .A2(new_n386), .A3(new_n631), .A4(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n680), .B1(new_n686), .B2(new_n642), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n428), .A2(new_n432), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n410), .A2(new_n413), .A3(G179), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n358), .A2(new_n693), .A3(new_n313), .A4(new_n353), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n433), .A2(new_n313), .A3(G179), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n358), .A2(new_n353), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n421), .ZN(new_n699));
  AOI211_X1 g0499(.A(new_n695), .B(new_n299), .C1(new_n311), .C2(new_n312), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n358), .A2(new_n693), .A3(new_n700), .A4(new_n353), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT31), .B1(new_n702), .B2(new_n652), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n387), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n640), .B1(new_n464), .B2(new_n440), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n646), .A4(new_n680), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n690), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT85), .B1(new_n689), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n709), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT85), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n681), .A2(new_n711), .A3(new_n712), .A4(new_n688), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n678), .B1(new_n714), .B2(G1), .ZN(G364));
  NOR2_X1   g0515(.A1(new_n547), .A2(G20), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G45), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT86), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n674), .A2(new_n718), .A3(new_n206), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n657), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G330), .B2(new_n655), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n210), .A2(new_n267), .ZN(new_n722));
  INV_X1    g0522(.A(G355), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n722), .A2(new_n723), .B1(G116), .B2(new_n210), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n673), .A2(new_n267), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n293), .B2(new_n231), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n243), .A2(new_n293), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n547), .A2(new_n255), .A3(KEYINPUT87), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT87), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G13), .B2(G33), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n207), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT88), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n228), .B1(G20), .B2(new_n332), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n719), .B1(new_n729), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n207), .A2(new_n314), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n741), .A2(new_n329), .A3(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n215), .B1(new_n744), .B2(new_n202), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n271), .B(new_n745), .C1(G77), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n207), .A2(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n434), .A3(new_n329), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G159), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(new_n434), .A3(G200), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n751), .A2(KEYINPUT32), .B1(new_n262), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n368), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n748), .A2(G190), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n740), .A2(G190), .A3(new_n329), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT89), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G58), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n434), .A2(G179), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n207), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n223), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n751), .B2(KEYINPUT32), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n747), .A2(new_n757), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n763), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G294), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n744), .B(KEYINPUT90), .ZN(new_n769));
  INV_X1    g0569(.A(G326), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n771), .A2(KEYINPUT91), .B1(G311), .B2(new_n746), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(KEYINPUT91), .B2(new_n771), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT92), .Z(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT33), .B(G317), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n750), .A2(G329), .B1(new_n742), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n758), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n267), .B1(new_n777), .B2(G322), .ZN(new_n778));
  INV_X1    g0578(.A(new_n752), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n756), .A2(G303), .B1(new_n779), .B2(G283), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n776), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n766), .B1(new_n774), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n739), .B1(new_n782), .B2(new_n736), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n655), .B2(new_n735), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n721), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n643), .A2(new_n680), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n613), .A2(new_n680), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n520), .A2(new_n517), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n680), .B1(new_n514), .B2(new_n516), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n518), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n792), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n680), .B(new_n794), .C1(new_n633), .C2(new_n642), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n719), .B1(new_n796), .B2(new_n711), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n711), .B2(new_n796), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n792), .A2(new_n733), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n267), .B(new_n764), .C1(G294), .C2(new_n777), .ZN(new_n800));
  INV_X1    g0600(.A(new_n744), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G303), .A2(new_n801), .B1(new_n750), .B2(G311), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G116), .A2(new_n746), .B1(new_n742), .B2(G283), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n752), .A2(new_n217), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G107), .B2(new_n756), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n800), .A2(new_n802), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n746), .A2(G159), .B1(new_n801), .B2(G137), .ZN(new_n807));
  INV_X1    g0607(.A(G150), .ZN(new_n808));
  INV_X1    g0608(.A(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n743), .C1(new_n759), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n267), .B1(new_n749), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT93), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n763), .A2(new_n221), .B1(new_n755), .B2(new_n202), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n752), .A2(new_n215), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n812), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n810), .A2(new_n811), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n806), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n736), .ZN(new_n822));
  INV_X1    g0622(.A(new_n719), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n733), .A2(new_n736), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n254), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n799), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n798), .A2(new_n826), .ZN(G384));
  NAND2_X1  g0627(.A1(new_n322), .A2(KEYINPUT35), .ZN(new_n828));
  OAI211_X1 g0628(.A(G116), .B(new_n229), .C1(new_n322), .C2(KEYINPUT35), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT94), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT36), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n231), .B(G77), .C1(new_n221), .C2(new_n215), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n202), .A2(G68), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n206), .B(G13), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT40), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT95), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n561), .B2(new_n564), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n582), .A2(KEYINPUT95), .A3(new_n563), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n840), .A2(new_n841), .A3(new_n567), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n560), .B1(new_n842), .B2(new_n566), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n590), .B1(new_n843), .B2(new_n577), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n650), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT37), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n581), .A2(new_n585), .ZN(new_n847));
  INV_X1    g0647(.A(new_n650), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n585), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n847), .A2(new_n849), .A3(new_n850), .A4(new_n590), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n596), .A2(new_n845), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n705), .A2(new_n708), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n551), .A2(new_n652), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n612), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n611), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n603), .B1(new_n553), .B2(new_n556), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n858), .A2(new_n859), .A3(new_n794), .A4(new_n864), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n859), .A2(new_n864), .A3(new_n794), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n847), .A2(new_n849), .A3(new_n590), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n851), .ZN(new_n869));
  INV_X1    g0669(.A(new_n849), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n596), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n855), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n838), .B1(new_n873), .B2(new_n857), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n838), .A2(new_n865), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n875), .A2(new_n620), .A3(new_n859), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n620), .B2(new_n859), .ZN(new_n877));
  OR3_X1    g0677(.A1(new_n876), .A2(new_n877), .A3(new_n690), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT96), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n872), .B2(new_n855), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT39), .B1(new_n858), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(KEYINPUT96), .A2(KEYINPUT39), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n873), .A2(new_n857), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n611), .A2(new_n652), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n884), .A2(new_n885), .B1(new_n617), .B2(new_n650), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n599), .A2(new_n602), .A3(new_n600), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n557), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n860), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(new_n889), .B1(new_n611), .B2(new_n861), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n795), .B2(new_n788), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n858), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n689), .A2(new_n620), .ZN(new_n894));
  INV_X1    g0694(.A(new_n619), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n893), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n878), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n206), .B2(new_n716), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n878), .A2(new_n897), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n837), .B1(new_n899), .B2(new_n900), .ZN(G367));
  OAI21_X1  g0701(.A(new_n331), .B1(new_n328), .B2(new_n680), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n684), .A2(new_n652), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n669), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n316), .B1(new_n902), .B2(new_n474), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n905), .A2(KEYINPUT42), .B1(new_n680), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(KEYINPUT42), .B2(new_n905), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT43), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n385), .A2(new_n680), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n381), .A3(new_n386), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(KEYINPUT97), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n910), .A2(new_n381), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(KEYINPUT97), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n908), .B1(new_n909), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n909), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT98), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n666), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n904), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n674), .B(KEYINPUT41), .Z(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT99), .B1(new_n671), .B2(new_n904), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n659), .A2(new_n663), .A3(new_n660), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n663), .B1(new_n659), .B2(new_n660), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n667), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n670), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT99), .ZN(new_n931));
  INV_X1    g0731(.A(new_n904), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n925), .A2(KEYINPUT44), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT44), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n931), .B1(new_n930), .B2(new_n932), .ZN(new_n936));
  AOI211_X1 g0736(.A(KEYINPUT99), .B(new_n904), .C1(new_n928), .C2(new_n929), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n928), .A2(new_n929), .A3(new_n904), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT45), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n921), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n665), .A2(new_n667), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n944), .A2(new_n656), .A3(new_n669), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n656), .B1(new_n944), .B2(new_n669), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n710), .B2(new_n713), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n934), .A2(new_n938), .A3(new_n666), .A4(new_n941), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n943), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT100), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT100), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n943), .A2(new_n952), .A3(new_n948), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n924), .B1(new_n954), .B2(new_n714), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n718), .A2(new_n206), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n923), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n726), .A2(new_n239), .B1(new_n210), .B2(new_n378), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n719), .B1(new_n959), .B2(new_n738), .ZN(new_n960));
  INV_X1    g0760(.A(G159), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n267), .B1(new_n755), .B2(new_n221), .C1(new_n743), .C2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n752), .A2(new_n254), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n763), .A2(new_n215), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n746), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n966), .A2(new_n202), .B1(new_n758), .B2(new_n808), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G137), .B2(new_n750), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n965), .B(new_n968), .C1(new_n809), .C2(new_n769), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n756), .A2(G116), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT46), .ZN(new_n971));
  INV_X1    g0771(.A(G303), .ZN(new_n972));
  INV_X1    g0772(.A(G311), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n971), .B1(new_n972), .B2(new_n759), .C1(new_n973), .C2(new_n769), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n742), .A2(G294), .B1(G317), .B2(new_n750), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n752), .A2(new_n223), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G107), .B2(new_n767), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n267), .B1(new_n746), .B2(G283), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n969), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n960), .B1(new_n981), .B2(new_n736), .ZN(new_n982));
  INV_X1    g0782(.A(new_n916), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(new_n735), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n958), .A2(new_n984), .ZN(G387));
  NAND3_X1  g0785(.A1(new_n710), .A2(new_n947), .A3(new_n713), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT105), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n948), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(new_n987), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n988), .A2(new_n674), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n676), .A2(new_n722), .B1(G107), .B2(new_n210), .ZN(new_n992));
  INV_X1    g0792(.A(new_n236), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n726), .B1(new_n993), .B2(G45), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n676), .B(new_n293), .C1(new_n215), .C2(new_n254), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT101), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(KEYINPUT101), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n512), .A2(KEYINPUT50), .A3(G50), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT50), .B1(new_n512), .B2(G50), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n992), .B1(new_n994), .B2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT102), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n738), .B1(new_n1001), .B2(KEYINPUT102), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n823), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n758), .A2(new_n202), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n744), .A2(new_n961), .B1(new_n749), .B2(new_n808), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G68), .C2(new_n746), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n271), .B(new_n976), .C1(new_n476), .C2(new_n742), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n767), .A2(new_n509), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n756), .A2(G77), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n767), .A2(G283), .B1(new_n756), .B2(G294), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G303), .A2(new_n746), .B1(new_n742), .B2(G311), .ZN(new_n1013));
  INV_X1    g0813(.A(G322), .ZN(new_n1014));
  INV_X1    g0814(.A(G317), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1013), .B1(new_n769), .B2(new_n1014), .C1(new_n1015), .C2(new_n759), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT103), .Z(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(KEYINPUT49), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n267), .B1(new_n750), .B2(G326), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n339), .C2(new_n752), .ZN(new_n1023));
  AOI21_X1  g0823(.A(KEYINPUT49), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1011), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT104), .Z(new_n1026));
  OAI221_X1 g0826(.A(new_n1004), .B1(new_n665), .B2(new_n735), .C1(new_n1026), .C2(new_n737), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n945), .A2(new_n946), .A3(new_n957), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n991), .A2(new_n1029), .ZN(G393));
  NAND2_X1  g0830(.A1(new_n725), .A2(new_n246), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n223), .B2(new_n210), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n719), .B1(new_n1032), .B2(new_n738), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n743), .A2(new_n972), .B1(new_n749), .B2(new_n1014), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n267), .B(new_n1034), .C1(G294), .C2(new_n746), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n758), .A2(new_n973), .B1(new_n744), .B2(new_n1015), .ZN(new_n1036));
  XOR2_X1   g0836(.A(KEYINPUT107), .B(KEYINPUT52), .Z(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n767), .A2(G116), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n756), .A2(G283), .B1(new_n779), .B2(G107), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n758), .A2(new_n961), .B1(new_n744), .B2(new_n808), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT51), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n271), .B1(new_n742), .B2(G50), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n746), .A2(new_n476), .B1(G143), .B2(new_n750), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n755), .A2(new_n215), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n804), .B(new_n1046), .C1(G77), .C2(new_n767), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT106), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1041), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1033), .B1(new_n1052), .B2(new_n736), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT108), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n735), .B2(new_n904), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n943), .A2(new_n949), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1056), .B2(new_n956), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n674), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1056), .B2(new_n989), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1057), .B1(new_n954), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1060), .A2(KEYINPUT109), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT109), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1062), .B(new_n1057), .C1(new_n954), .C2(new_n1059), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G390));
  NAND3_X1  g0865(.A1(new_n709), .A2(new_n794), .A3(new_n864), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n881), .B(new_n883), .C1(new_n891), .C2(new_n885), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n680), .B(new_n791), .C1(new_n686), .C2(new_n642), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n788), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n864), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n885), .B1(new_n873), .B2(new_n857), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1066), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n694), .A2(new_n695), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n311), .A2(new_n312), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n299), .ZN(new_n1077));
  AOI21_X1  g0877(.A(G179), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n421), .A2(new_n437), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n348), .A2(new_n354), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n701), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n652), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT31), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n475), .A2(new_n387), .A3(new_n652), .ZN(new_n1087));
  OAI211_X1 g0887(.A(G330), .B(new_n794), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(KEYINPUT110), .B1(new_n1088), .B2(new_n890), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT110), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n709), .A2(new_n1090), .A3(new_n794), .A4(new_n864), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1073), .B1(new_n1074), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n881), .A2(new_n733), .A3(new_n883), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n824), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n719), .B1(new_n476), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n267), .B(new_n817), .C1(G283), .C2(new_n801), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n254), .B2(new_n763), .C1(new_n217), .C2(new_n755), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n746), .A2(G97), .B1(G294), .B2(new_n750), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n262), .B2(new_n743), .C1(new_n339), .C2(new_n758), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n271), .B1(new_n746), .B2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n202), .B2(new_n752), .C1(new_n961), .C2(new_n763), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n742), .A2(G137), .B1(new_n777), .B2(G132), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G128), .A2(new_n801), .B1(new_n750), .B2(G125), .ZN(new_n1107));
  OR3_X1    g0907(.A1(new_n755), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT53), .B1(new_n755), .B2(new_n808), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1099), .A2(new_n1101), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1111), .A2(KEYINPUT115), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n737), .B1(new_n1111), .B2(KEYINPUT115), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1097), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1094), .A2(new_n957), .B1(new_n1095), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT112), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1088), .A2(new_n890), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n788), .A3(new_n1068), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1092), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1069), .B1(new_n890), .B2(new_n1088), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1120), .A2(KEYINPUT112), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT111), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1088), .A2(new_n1123), .A3(new_n890), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n795), .A2(new_n788), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1066), .A2(new_n1117), .A3(KEYINPUT111), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n620), .A2(new_n709), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n894), .A2(new_n1130), .A3(new_n895), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1094), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(KEYINPUT113), .A3(new_n674), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT114), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1135), .A3(new_n1132), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1119), .A2(new_n1121), .B1(new_n1127), .B2(new_n1126), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT114), .B1(new_n1137), .B2(new_n1131), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1093), .A2(new_n1067), .A3(new_n1072), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1074), .B2(new_n1066), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1134), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT113), .B1(new_n1133), .B2(new_n674), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1115), .B1(new_n1142), .B2(new_n1143), .ZN(G378));
  INV_X1    g0944(.A(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1131), .A2(KEYINPUT120), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT120), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n894), .A2(new_n1130), .A3(new_n1147), .A4(new_n895), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1131), .B1(new_n1122), .B2(new_n1128), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n1094), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n484), .A2(new_n650), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n502), .B(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1153), .B(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n875), .B2(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n865), .A2(new_n838), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n866), .A2(new_n874), .ZN(new_n1159));
  AND4_X1   g0959(.A1(G330), .A2(new_n1158), .A3(new_n1156), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n893), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(G330), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1156), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1158), .A2(new_n1156), .A3(new_n1159), .A4(G330), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1164), .A2(new_n892), .A3(new_n886), .A4(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1145), .B1(new_n1151), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1140), .A2(new_n1137), .A3(new_n1131), .ZN(new_n1170));
  OAI211_X1 g0970(.A(KEYINPUT57), .B(new_n1169), .C1(new_n1170), .C2(new_n1149), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n1171), .A3(new_n674), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1163), .A2(new_n733), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n719), .B1(G50), .B2(new_n1096), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G97), .A2(new_n742), .B1(new_n746), .B2(new_n509), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT117), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G41), .B(new_n267), .C1(new_n750), .C2(G283), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n777), .A2(G107), .B1(new_n801), .B2(G116), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1010), .B1(new_n215), .B2(new_n763), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G58), .B2(new_n779), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1180), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1182));
  INV_X1    g0982(.A(G41), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n255), .A2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT116), .ZN(new_n1185));
  AOI21_X1  g0985(.A(G50), .B1(new_n271), .B2(new_n1183), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1181), .A2(new_n1182), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1185), .B1(G124), .B2(new_n750), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n746), .A2(G137), .B1(new_n777), .B2(G128), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n813), .B2(new_n743), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G150), .A2(new_n767), .B1(new_n801), .B2(G125), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT119), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n756), .C2(new_n1103), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT59), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1188), .B1(new_n961), .B2(new_n752), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1187), .B1(new_n1182), .B2(new_n1181), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1174), .B1(new_n1197), .B2(new_n736), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1169), .A2(new_n957), .B1(new_n1173), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1172), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT121), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT121), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1172), .A2(new_n1202), .A3(new_n1199), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(G375));
  INV_X1    g1005(.A(new_n924), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1137), .A2(new_n1131), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1136), .A2(new_n1138), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n890), .A2(new_n733), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n221), .A2(new_n752), .B1(new_n755), .B2(new_n961), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n750), .A2(G128), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(new_n267), .C1(new_n808), .C2(new_n966), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(G50), .C2(new_n767), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT122), .Z(new_n1214));
  OAI22_X1  g1014(.A1(new_n743), .A2(new_n1102), .B1(new_n744), .B2(new_n813), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n760), .B2(G137), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n267), .B(new_n963), .C1(G294), .C2(new_n801), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n746), .A2(G107), .B1(new_n777), .B2(G283), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n742), .A2(G116), .B1(G303), .B2(new_n750), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n767), .A2(new_n509), .B1(new_n756), .B2(G97), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n737), .B1(new_n1217), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n823), .B(new_n1223), .C1(new_n215), .C2(new_n824), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1129), .A2(new_n957), .B1(new_n1209), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1208), .A2(new_n1225), .ZN(G381));
  NOR2_X1   g1026(.A1(G393), .A2(G396), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n798), .A3(new_n826), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(G390), .A2(G387), .A3(G381), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G378), .A2(KEYINPUT123), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT123), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1231), .B(new_n1115), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1229), .A2(new_n1204), .A3(new_n1233), .ZN(G407));
  NAND2_X1  g1034(.A1(new_n651), .A2(G213), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT124), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1204), .A2(new_n1233), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(G407), .A2(G213), .A3(new_n1237), .ZN(G409));
  INV_X1    g1038(.A(KEYINPUT61), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1169), .B1(new_n1170), .B2(new_n1149), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1199), .B1(new_n1240), .B2(new_n924), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1230), .A2(new_n1232), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G378), .A2(new_n1199), .A3(new_n1172), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1236), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1150), .A2(new_n1058), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1207), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT60), .B1(new_n1207), .B2(KEYINPUT125), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1225), .B1(G384), .B2(KEYINPUT126), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1245), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1249), .A2(new_n1245), .A3(new_n1251), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(G2897), .A3(new_n1236), .A4(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1254), .ZN(new_n1256));
  INV_X1    g1056(.A(G2897), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1236), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1256), .A2(new_n1252), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1239), .B1(new_n1244), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1258), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1256), .A2(new_n1252), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1263), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(new_n1064), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n785), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n958), .B(new_n984), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1266), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1244), .A2(KEYINPUT63), .A3(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1262), .A2(new_n1267), .A3(new_n1273), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1244), .A2(new_n1277), .A3(new_n1274), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1244), .B2(new_n1274), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1278), .A2(new_n1261), .A3(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1276), .B1(new_n1280), .B2(new_n1273), .ZN(G405));
  INV_X1    g1081(.A(KEYINPUT127), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1201), .A2(new_n1203), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1283), .A2(new_n1243), .A3(new_n1266), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1266), .B1(new_n1283), .B2(new_n1243), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1282), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1243), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1274), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1283), .A2(new_n1243), .A3(new_n1266), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(KEYINPUT127), .A3(new_n1289), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1286), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1273), .A2(KEYINPUT127), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(G402));
endmodule


