

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772;

  AND2_X1 U370 ( .A1(n418), .A2(n415), .ZN(n360) );
  XNOR2_X2 U371 ( .A(n441), .B(n440), .ZN(n553) );
  INV_X2 U372 ( .A(G953), .ZN(n763) );
  NAND2_X1 U373 ( .A1(n483), .A2(n431), .ZN(n365) );
  XNOR2_X2 U374 ( .A(n589), .B(KEYINPUT38), .ZN(n624) );
  INV_X2 U375 ( .A(n493), .ZN(n589) );
  INV_X2 U376 ( .A(G125), .ZN(n430) );
  AND2_X1 U377 ( .A1(n411), .A2(n581), .ZN(n410) );
  NAND2_X1 U378 ( .A1(n592), .A2(n591), .ZN(n593) );
  AND2_X1 U379 ( .A1(n401), .A2(n400), .ZN(n399) );
  OR2_X1 U380 ( .A1(n639), .A2(n455), .ZN(n348) );
  XNOR2_X1 U381 ( .A(n588), .B(KEYINPUT82), .ZN(n545) );
  XNOR2_X1 U382 ( .A(n395), .B(n393), .ZN(n548) );
  XOR2_X1 U383 ( .A(KEYINPUT59), .B(n707), .Z(n708) );
  XOR2_X1 U384 ( .A(G134), .B(G131), .Z(n462) );
  NOR2_X1 U385 ( .A1(n639), .A2(n455), .ZN(n569) );
  AND2_X1 U386 ( .A1(n575), .A2(n349), .ZN(n689) );
  AND2_X1 U387 ( .A1(n640), .A2(n561), .ZN(n349) );
  NOR2_X1 U388 ( .A1(n553), .A2(n521), .ZN(n522) );
  NAND2_X2 U389 ( .A1(n606), .A2(n362), .ZN(n732) );
  XNOR2_X2 U390 ( .A(n386), .B(KEYINPUT115), .ZN(n606) );
  XNOR2_X2 U391 ( .A(n370), .B(KEYINPUT79), .ZN(n592) );
  NOR2_X1 U392 ( .A1(n639), .A2(n640), .ZN(n564) );
  XNOR2_X1 U393 ( .A(KEYINPUT67), .B(G101), .ZN(n445) );
  XOR2_X1 U394 ( .A(KEYINPUT8), .B(n427), .Z(n513) );
  NOR2_X1 U395 ( .A1(n743), .A2(n582), .ZN(n669) );
  INV_X1 U396 ( .A(G146), .ZN(n449) );
  NAND2_X1 U397 ( .A1(n522), .A2(n634), .ZN(n384) );
  INV_X1 U398 ( .A(KEYINPUT30), .ZN(n372) );
  INV_X1 U399 ( .A(KEYINPUT28), .ZN(n596) );
  INV_X1 U400 ( .A(KEYINPUT0), .ZN(n542) );
  XNOR2_X1 U401 ( .A(G107), .B(G104), .ZN(n448) );
  XOR2_X1 U402 ( .A(G140), .B(G131), .Z(n499) );
  XNOR2_X1 U403 ( .A(n391), .B(n387), .ZN(n502) );
  XNOR2_X1 U404 ( .A(n500), .B(n501), .ZN(n391) );
  XNOR2_X1 U405 ( .A(n389), .B(n388), .ZN(n387) );
  XNOR2_X1 U406 ( .A(G143), .B(G104), .ZN(n500) );
  XNOR2_X1 U407 ( .A(n530), .B(n529), .ZN(n656) );
  NAND2_X1 U408 ( .A1(n564), .A2(n555), .ZN(n530) );
  XNOR2_X1 U409 ( .A(n738), .B(KEYINPUT107), .ZN(n571) );
  INV_X1 U410 ( .A(KEYINPUT1), .ZN(n406) );
  XNOR2_X1 U411 ( .A(n506), .B(n394), .ZN(n393) );
  OR2_X1 U412 ( .A1(n707), .A2(G902), .ZN(n395) );
  INV_X1 U413 ( .A(G475), .ZN(n394) );
  OR2_X1 U414 ( .A1(n422), .A2(n417), .ZN(n416) );
  INV_X1 U415 ( .A(n571), .ZN(n392) );
  XNOR2_X1 U416 ( .A(G146), .B(G137), .ZN(n468) );
  XOR2_X1 U417 ( .A(KEYINPUT77), .B(KEYINPUT99), .Z(n469) );
  INV_X1 U418 ( .A(KEYINPUT70), .ZN(n374) );
  XNOR2_X1 U419 ( .A(n390), .B(G113), .ZN(n389) );
  INV_X1 U420 ( .A(G122), .ZN(n390) );
  XNOR2_X1 U421 ( .A(KEYINPUT12), .B(KEYINPUT101), .ZN(n388) );
  XNOR2_X1 U422 ( .A(KEYINPUT102), .B(KEYINPUT11), .ZN(n501) );
  INV_X1 U423 ( .A(KEYINPUT45), .ZN(n412) );
  NAND2_X1 U424 ( .A1(n410), .A2(n408), .ZN(n407) );
  XNOR2_X1 U425 ( .A(G107), .B(G134), .ZN(n507) );
  XOR2_X1 U426 ( .A(G122), .B(G116), .Z(n508) );
  XNOR2_X1 U427 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U428 ( .A(KEYINPUT90), .ZN(n533) );
  NAND2_X1 U429 ( .A1(n399), .A2(n396), .ZN(n404) );
  NAND2_X1 U430 ( .A1(n398), .A2(n397), .ZN(n396) );
  NAND2_X1 U431 ( .A1(n656), .A2(n402), .ZN(n400) );
  XNOR2_X1 U432 ( .A(n479), .B(n372), .ZN(n371) );
  AND2_X1 U433 ( .A1(n569), .A2(n414), .ZN(n373) );
  INV_X1 U434 ( .A(n640), .ZN(n405) );
  XNOR2_X1 U435 ( .A(KEYINPUT24), .B(G128), .ZN(n428) );
  XNOR2_X1 U436 ( .A(n504), .B(n505), .ZN(n707) );
  NOR2_X1 U437 ( .A1(n763), .A2(G952), .ZN(n718) );
  NOR2_X1 U438 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U439 ( .A(n610), .B(KEYINPUT40), .ZN(n772) );
  XNOR2_X1 U440 ( .A(n567), .B(n566), .ZN(n737) );
  XNOR2_X1 U441 ( .A(n520), .B(KEYINPUT106), .ZN(n738) );
  XNOR2_X1 U442 ( .A(G140), .B(G137), .ZN(n350) );
  INV_X1 U443 ( .A(n609), .ZN(n423) );
  AND2_X1 U444 ( .A1(n425), .A2(n424), .ZN(n351) );
  AND2_X1 U445 ( .A1(n674), .A2(n673), .ZN(n352) );
  NAND2_X1 U446 ( .A1(n392), .A2(n423), .ZN(n425) );
  AND2_X1 U447 ( .A1(n563), .A2(n379), .ZN(n353) );
  XOR2_X1 U448 ( .A(KEYINPUT16), .B(G122), .Z(n354) );
  XOR2_X1 U449 ( .A(KEYINPUT95), .B(KEYINPUT3), .Z(n355) );
  NOR2_X1 U450 ( .A1(n526), .A2(n405), .ZN(n356) );
  NOR2_X1 U451 ( .A1(n574), .A2(n405), .ZN(n357) );
  OR2_X1 U452 ( .A1(KEYINPUT89), .A2(KEYINPUT44), .ZN(n358) );
  BUF_X1 U453 ( .A(n676), .Z(n359) );
  NAND2_X1 U454 ( .A1(n599), .A2(n600), .ZN(n386) );
  NAND2_X1 U455 ( .A1(n404), .A2(n545), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n605), .B(n604), .ZN(n658) );
  AND2_X2 U457 ( .A1(n678), .A2(n677), .ZN(n361) );
  AND2_X2 U458 ( .A1(n678), .A2(n677), .ZN(n712) );
  BUF_X1 U459 ( .A(n601), .Z(n362) );
  XNOR2_X1 U460 ( .A(n583), .B(n535), .ZN(n601) );
  NAND2_X1 U461 ( .A1(n568), .A2(n550), .ZN(n552) );
  NAND2_X1 U462 ( .A1(n363), .A2(n364), .ZN(n366) );
  NAND2_X1 U463 ( .A1(n365), .A2(n366), .ZN(n496) );
  INV_X1 U464 ( .A(n483), .ZN(n363) );
  INV_X1 U465 ( .A(n431), .ZN(n364) );
  XNOR2_X1 U466 ( .A(KEYINPUT69), .B(KEYINPUT10), .ZN(n431) );
  XNOR2_X1 U467 ( .A(n758), .B(n433), .ZN(n434) );
  XNOR2_X1 U468 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X2 U469 ( .A(KEYINPUT42), .B(n607), .ZN(n771) );
  XNOR2_X1 U470 ( .A(n378), .B(KEYINPUT75), .ZN(n377) );
  XNOR2_X1 U471 ( .A(n375), .B(n374), .ZN(n615) );
  NOR2_X2 U472 ( .A1(n367), .A2(n743), .ZN(n676) );
  NAND2_X1 U473 ( .A1(n756), .A2(n757), .ZN(n367) );
  BUF_X1 U474 ( .A(n475), .Z(n368) );
  BUF_X1 U475 ( .A(n715), .Z(n369) );
  NAND2_X1 U476 ( .A1(n373), .A2(n371), .ZN(n370) );
  NAND2_X1 U477 ( .A1(n377), .A2(n376), .ZN(n375) );
  INV_X1 U478 ( .A(n740), .ZN(n376) );
  NAND2_X1 U479 ( .A1(n385), .A2(n426), .ZN(n378) );
  INV_X1 U480 ( .A(n379), .ZN(n380) );
  NAND2_X1 U481 ( .A1(n577), .A2(n379), .ZN(n578) );
  XNOR2_X2 U482 ( .A(n559), .B(KEYINPUT32), .ZN(n379) );
  XNOR2_X1 U483 ( .A(n380), .B(n690), .ZN(G21) );
  NAND2_X1 U484 ( .A1(n353), .A2(n381), .ZN(n409) );
  NAND2_X1 U485 ( .A1(n383), .A2(n382), .ZN(n381) );
  INV_X1 U486 ( .A(KEYINPUT89), .ZN(n382) );
  INV_X1 U487 ( .A(n579), .ZN(n383) );
  BUF_X1 U488 ( .A(n579), .Z(n691) );
  XNOR2_X2 U489 ( .A(n384), .B(KEYINPUT71), .ZN(n595) );
  NAND2_X1 U490 ( .A1(n421), .A2(n351), .ZN(n420) );
  XNOR2_X2 U491 ( .A(n444), .B(KEYINPUT68), .ZN(n639) );
  NAND2_X1 U492 ( .A1(n360), .A2(n420), .ZN(n385) );
  NOR2_X1 U493 ( .A1(n656), .A2(n402), .ZN(n397) );
  INV_X1 U494 ( .A(n565), .ZN(n398) );
  NAND2_X1 U495 ( .A1(n565), .A2(n402), .ZN(n401) );
  INV_X1 U496 ( .A(KEYINPUT34), .ZN(n402) );
  XNOR2_X2 U497 ( .A(n403), .B(n546), .ZN(n579) );
  XNOR2_X2 U498 ( .A(n599), .B(n406), .ZN(n640) );
  XNOR2_X2 U499 ( .A(n407), .B(n412), .ZN(n743) );
  NAND2_X1 U500 ( .A1(n409), .A2(n358), .ZN(n408) );
  NAND2_X1 U501 ( .A1(n580), .A2(n579), .ZN(n411) );
  XNOR2_X2 U502 ( .A(n413), .B(G143), .ZN(n514) );
  XNOR2_X2 U503 ( .A(G128), .B(KEYINPUT65), .ZN(n413) );
  XNOR2_X1 U504 ( .A(n471), .B(n354), .ZN(n751) );
  XNOR2_X1 U505 ( .A(n467), .B(n355), .ZN(n471) );
  INV_X1 U506 ( .A(n521), .ZN(n414) );
  NOR2_X1 U507 ( .A1(n732), .A2(n417), .ZN(n421) );
  OR2_X1 U508 ( .A1(n571), .A2(n416), .ZN(n415) );
  INV_X1 U509 ( .A(n594), .ZN(n417) );
  NAND2_X1 U510 ( .A1(n732), .A2(n419), .ZN(n418) );
  AND2_X1 U511 ( .A1(n603), .A2(n594), .ZN(n419) );
  XNOR2_X1 U512 ( .A(n770), .B(KEYINPUT85), .ZN(n426) );
  XNOR2_X2 U513 ( .A(n593), .B(KEYINPUT113), .ZN(n770) );
  NAND2_X1 U514 ( .A1(n423), .A2(n603), .ZN(n422) );
  INV_X1 U515 ( .A(n603), .ZN(n424) );
  INV_X1 U516 ( .A(n425), .ZN(n628) );
  XNOR2_X2 U517 ( .A(n475), .B(n749), .ZN(n486) );
  XNOR2_X2 U518 ( .A(G119), .B(G116), .ZN(n466) );
  XNOR2_X2 U519 ( .A(G113), .B(KEYINPUT72), .ZN(n465) );
  XNOR2_X2 U520 ( .A(n761), .B(n446), .ZN(n475) );
  XNOR2_X2 U521 ( .A(n514), .B(KEYINPUT4), .ZN(n761) );
  XNOR2_X2 U522 ( .A(n617), .B(n616), .ZN(n756) );
  XNOR2_X1 U523 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n611) );
  XNOR2_X1 U524 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U525 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U526 ( .A(n432), .B(G119), .ZN(n433) );
  XNOR2_X1 U527 ( .A(n759), .B(n451), .ZN(n452) );
  XNOR2_X1 U528 ( .A(n596), .B(KEYINPUT114), .ZN(n597) );
  XNOR2_X1 U529 ( .A(n473), .B(n472), .ZN(n474) );
  INV_X1 U530 ( .A(KEYINPUT41), .ZN(n604) );
  INV_X1 U531 ( .A(n692), .ZN(n693) );
  XNOR2_X1 U532 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n566) );
  XNOR2_X1 U533 ( .A(n665), .B(n664), .ZN(G75) );
  NAND2_X1 U534 ( .A1(G234), .A2(n763), .ZN(n427) );
  NAND2_X1 U535 ( .A1(G221), .A2(n513), .ZN(n429) );
  XNOR2_X1 U536 ( .A(n429), .B(n428), .ZN(n435) );
  XNOR2_X2 U537 ( .A(n430), .B(G146), .ZN(n483) );
  XNOR2_X2 U538 ( .A(n496), .B(n350), .ZN(n758) );
  XOR2_X1 U539 ( .A(G110), .B(KEYINPUT23), .Z(n432) );
  XNOR2_X1 U540 ( .A(n434), .B(n435), .ZN(n692) );
  INV_X1 U541 ( .A(G902), .ZN(n518) );
  NAND2_X1 U542 ( .A1(n692), .A2(n518), .ZN(n441) );
  XOR2_X1 U543 ( .A(KEYINPUT25), .B(KEYINPUT98), .Z(n439) );
  XNOR2_X1 U544 ( .A(KEYINPUT94), .B(KEYINPUT15), .ZN(n436) );
  XNOR2_X1 U545 ( .A(n436), .B(G902), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n487), .A2(G234), .ZN(n437) );
  XNOR2_X1 U547 ( .A(n437), .B(KEYINPUT20), .ZN(n442) );
  NAND2_X1 U548 ( .A1(n442), .A2(G217), .ZN(n438) );
  XNOR2_X1 U549 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U550 ( .A1(n442), .A2(G221), .ZN(n443) );
  XNOR2_X1 U551 ( .A(n443), .B(KEYINPUT21), .ZN(n549) );
  INV_X1 U552 ( .A(n549), .ZN(n634) );
  NAND2_X1 U553 ( .A1(n553), .A2(n634), .ZN(n444) );
  XNOR2_X1 U554 ( .A(n445), .B(KEYINPUT66), .ZN(n446) );
  XNOR2_X1 U555 ( .A(KEYINPUT78), .B(G110), .ZN(n447) );
  XNOR2_X1 U556 ( .A(n448), .B(n447), .ZN(n749) );
  XOR2_X1 U557 ( .A(KEYINPUT97), .B(n462), .Z(n759) );
  NAND2_X1 U558 ( .A1(G227), .A2(n763), .ZN(n450) );
  XNOR2_X1 U559 ( .A(n452), .B(n350), .ZN(n453) );
  XNOR2_X1 U560 ( .A(n486), .B(n453), .ZN(n682) );
  NAND2_X1 U561 ( .A1(n682), .A2(n518), .ZN(n454) );
  XNOR2_X2 U562 ( .A(n454), .B(G469), .ZN(n599) );
  INV_X1 U563 ( .A(n599), .ZN(n455) );
  NAND2_X1 U564 ( .A1(G237), .A2(G234), .ZN(n457) );
  INV_X1 U565 ( .A(KEYINPUT14), .ZN(n456) );
  XNOR2_X1 U566 ( .A(n457), .B(n456), .ZN(n652) );
  NAND2_X1 U567 ( .A1(G953), .A2(G902), .ZN(n536) );
  NOR2_X1 U568 ( .A1(n652), .A2(n536), .ZN(n458) );
  XNOR2_X1 U569 ( .A(n458), .B(KEYINPUT111), .ZN(n459) );
  NOR2_X1 U570 ( .A1(G900), .A2(n459), .ZN(n461) );
  NAND2_X1 U571 ( .A1(G952), .A2(n763), .ZN(n537) );
  NOR2_X1 U572 ( .A1(n652), .A2(n537), .ZN(n460) );
  NOR2_X1 U573 ( .A1(n461), .A2(n460), .ZN(n521) );
  XOR2_X1 U574 ( .A(n462), .B(KEYINPUT5), .Z(n464) );
  NOR2_X1 U575 ( .A1(G953), .A2(G237), .ZN(n497) );
  NAND2_X1 U576 ( .A1(n497), .A2(G210), .ZN(n463) );
  XNOR2_X1 U577 ( .A(n464), .B(n463), .ZN(n473) );
  XNOR2_X1 U578 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U579 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U580 ( .A(n368), .B(n474), .ZN(n698) );
  NAND2_X1 U581 ( .A1(n698), .A2(n518), .ZN(n477) );
  XOR2_X1 U582 ( .A(KEYINPUT73), .B(G472), .Z(n476) );
  XNOR2_X2 U583 ( .A(n477), .B(n476), .ZN(n637) );
  INV_X1 U584 ( .A(G237), .ZN(n478) );
  NAND2_X1 U585 ( .A1(n518), .A2(n478), .ZN(n489) );
  NAND2_X1 U586 ( .A1(n489), .A2(G214), .ZN(n623) );
  NAND2_X1 U587 ( .A1(n637), .A2(n623), .ZN(n479) );
  XNOR2_X1 U588 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n481) );
  NAND2_X1 U589 ( .A1(n763), .A2(G224), .ZN(n480) );
  XNOR2_X1 U590 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U591 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U592 ( .A(n751), .B(n484), .ZN(n485) );
  XNOR2_X1 U593 ( .A(n486), .B(n485), .ZN(n715) );
  INV_X1 U594 ( .A(n487), .ZN(n671) );
  NOR2_X1 U595 ( .A1(n715), .A2(n671), .ZN(n488) );
  INV_X1 U596 ( .A(n488), .ZN(n492) );
  NAND2_X1 U597 ( .A1(n489), .A2(G210), .ZN(n490) );
  XNOR2_X1 U598 ( .A(n490), .B(KEYINPUT96), .ZN(n491) );
  XNOR2_X1 U599 ( .A(n492), .B(n491), .ZN(n532) );
  INV_X1 U600 ( .A(n532), .ZN(n493) );
  NAND2_X1 U601 ( .A1(n592), .A2(n624), .ZN(n495) );
  XNOR2_X1 U602 ( .A(KEYINPUT88), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U603 ( .A(n495), .B(n494), .ZN(n608) );
  XNOR2_X1 U604 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n506) );
  BUF_X1 U605 ( .A(n496), .Z(n505) );
  NAND2_X1 U606 ( .A1(n497), .A2(G214), .ZN(n498) );
  XNOR2_X1 U607 ( .A(n499), .B(n498), .ZN(n503) );
  XNOR2_X1 U608 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U609 ( .A(n508), .B(n507), .ZN(n512) );
  XOR2_X1 U610 ( .A(KEYINPUT105), .B(KEYINPUT9), .Z(n510) );
  XNOR2_X1 U611 ( .A(KEYINPUT7), .B(KEYINPUT104), .ZN(n509) );
  XNOR2_X1 U612 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U613 ( .A(n512), .B(n511), .Z(n517) );
  NAND2_X1 U614 ( .A1(G217), .A2(n513), .ZN(n515) );
  XNOR2_X1 U615 ( .A(n514), .B(n515), .ZN(n516) );
  XNOR2_X1 U616 ( .A(n517), .B(n516), .ZN(n705) );
  NAND2_X1 U617 ( .A1(n705), .A2(n518), .ZN(n519) );
  XNOR2_X1 U618 ( .A(n519), .B(G478), .ZN(n544) );
  NAND2_X1 U619 ( .A1(n548), .A2(n544), .ZN(n520) );
  NAND2_X1 U620 ( .A1(n608), .A2(n571), .ZN(n742) );
  NOR2_X1 U621 ( .A1(n544), .A2(n548), .ZN(n609) );
  XOR2_X1 U622 ( .A(n609), .B(KEYINPUT110), .Z(n735) );
  INV_X1 U623 ( .A(n735), .ZN(n523) );
  NAND2_X1 U624 ( .A1(n595), .A2(n523), .ZN(n525) );
  INV_X1 U625 ( .A(KEYINPUT6), .ZN(n524) );
  XNOR2_X1 U626 ( .A(n637), .B(n524), .ZN(n555) );
  INV_X1 U627 ( .A(n555), .ZN(n573) );
  NOR2_X1 U628 ( .A1(n525), .A2(n573), .ZN(n585) );
  NAND2_X1 U629 ( .A1(n585), .A2(n623), .ZN(n526) );
  XNOR2_X1 U630 ( .A(KEYINPUT43), .B(KEYINPUT112), .ZN(n527) );
  XOR2_X1 U631 ( .A(n356), .B(n527), .Z(n528) );
  NAND2_X1 U632 ( .A1(n528), .A2(n589), .ZN(n688) );
  AND2_X1 U633 ( .A1(n742), .A2(n688), .ZN(n757) );
  INV_X1 U634 ( .A(n757), .ZN(n582) );
  INV_X1 U635 ( .A(KEYINPUT33), .ZN(n529) );
  INV_X1 U636 ( .A(n623), .ZN(n531) );
  NOR2_X2 U637 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X2 U638 ( .A(n534), .B(n533), .ZN(n583) );
  XNOR2_X1 U639 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n535) );
  NOR2_X1 U640 ( .A1(G898), .A2(n536), .ZN(n539) );
  INV_X1 U641 ( .A(n537), .ZN(n538) );
  NOR2_X1 U642 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U643 ( .A1(n540), .A2(n652), .ZN(n541) );
  NAND2_X1 U644 ( .A1(n601), .A2(n541), .ZN(n543) );
  XNOR2_X2 U645 ( .A(n543), .B(n542), .ZN(n568) );
  INV_X1 U646 ( .A(n568), .ZN(n565) );
  INV_X1 U647 ( .A(n544), .ZN(n547) );
  NOR2_X1 U648 ( .A1(n548), .A2(n547), .ZN(n588) );
  XNOR2_X1 U649 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n546) );
  NAND2_X1 U650 ( .A1(n548), .A2(n547), .ZN(n626) );
  NOR2_X1 U651 ( .A1(n626), .A2(n549), .ZN(n550) );
  XOR2_X1 U652 ( .A(KEYINPUT74), .B(KEYINPUT22), .Z(n551) );
  XNOR2_X2 U653 ( .A(n552), .B(n551), .ZN(n575) );
  BUF_X1 U654 ( .A(n553), .Z(n560) );
  XNOR2_X1 U655 ( .A(n560), .B(KEYINPUT108), .ZN(n633) );
  NOR2_X1 U656 ( .A1(n640), .A2(n633), .ZN(n554) );
  XNOR2_X1 U657 ( .A(n554), .B(KEYINPUT109), .ZN(n557) );
  XOR2_X1 U658 ( .A(KEYINPUT83), .B(n555), .Z(n556) );
  NOR2_X1 U659 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U660 ( .A1(n575), .A2(n558), .ZN(n559) );
  NOR2_X1 U661 ( .A1(n637), .A2(n560), .ZN(n561) );
  INV_X1 U662 ( .A(KEYINPUT44), .ZN(n562) );
  NOR2_X1 U663 ( .A1(n689), .A2(n562), .ZN(n563) );
  NAND2_X1 U664 ( .A1(n564), .A2(n637), .ZN(n645) );
  NOR2_X1 U665 ( .A1(n565), .A2(n645), .ZN(n567) );
  NOR2_X1 U666 ( .A1(n348), .A2(n637), .ZN(n570) );
  NAND2_X1 U667 ( .A1(n398), .A2(n570), .ZN(n724) );
  NAND2_X1 U668 ( .A1(n737), .A2(n724), .ZN(n572) );
  NAND2_X1 U669 ( .A1(n572), .A2(n425), .ZN(n576) );
  NAND2_X1 U670 ( .A1(n573), .A2(n633), .ZN(n574) );
  NAND2_X1 U671 ( .A1(n575), .A2(n357), .ZN(n721) );
  AND2_X1 U672 ( .A1(n576), .A2(n721), .ZN(n581) );
  NOR2_X1 U673 ( .A1(n689), .A2(KEYINPUT44), .ZN(n577) );
  NAND2_X1 U674 ( .A1(n578), .A2(n382), .ZN(n580) );
  INV_X1 U675 ( .A(n583), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U677 ( .A(n586), .B(KEYINPUT36), .ZN(n587) );
  NOR2_X1 U678 ( .A1(n640), .A2(n587), .ZN(n740) );
  INV_X1 U679 ( .A(n588), .ZN(n590) );
  NOR2_X1 U680 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U681 ( .A(KEYINPUT76), .ZN(n602) );
  NAND2_X1 U682 ( .A1(KEYINPUT47), .A2(n602), .ZN(n594) );
  NAND2_X1 U683 ( .A1(n595), .A2(n637), .ZN(n598) );
  XNOR2_X1 U684 ( .A(n598), .B(n597), .ZN(n600) );
  NOR2_X1 U685 ( .A1(KEYINPUT47), .A2(n602), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n624), .A2(n623), .ZN(n627) );
  NOR2_X1 U687 ( .A1(n626), .A2(n627), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n606), .A2(n658), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n771), .A2(n772), .ZN(n612) );
  INV_X1 U691 ( .A(n613), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n617) );
  INV_X1 U693 ( .A(KEYINPUT48), .ZN(n616) );
  INV_X1 U694 ( .A(n676), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n619), .A2(KEYINPUT84), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n618), .B(KEYINPUT2), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n619), .A2(KEYINPUT84), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n622), .B(KEYINPUT87), .ZN(n663) );
  NOR2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n630) );
  NOR2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U702 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U703 ( .A1(n631), .A2(n656), .ZN(n632) );
  XOR2_X1 U704 ( .A(KEYINPUT122), .B(n632), .Z(n650) );
  NOR2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U706 ( .A(KEYINPUT49), .B(n635), .Z(n636) );
  NOR2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U708 ( .A(n638), .B(KEYINPUT120), .ZN(n644) );
  XOR2_X1 U709 ( .A(KEYINPUT121), .B(KEYINPUT50), .Z(n642) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n642), .B(n641), .ZN(n643) );
  NAND2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U714 ( .A(KEYINPUT51), .B(n647), .Z(n648) );
  NAND2_X1 U715 ( .A1(n658), .A2(n648), .ZN(n649) );
  NAND2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U717 ( .A(KEYINPUT52), .B(n651), .Z(n655) );
  INV_X1 U718 ( .A(n652), .ZN(n653) );
  NAND2_X1 U719 ( .A1(n653), .A2(G952), .ZN(n654) );
  NOR2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n661) );
  INV_X1 U721 ( .A(n656), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U723 ( .A1(n659), .A2(n763), .ZN(n660) );
  NOR2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n665) );
  INV_X1 U726 ( .A(KEYINPUT53), .ZN(n664) );
  NAND2_X1 U727 ( .A1(n676), .A2(n671), .ZN(n667) );
  INV_X1 U728 ( .A(KEYINPUT86), .ZN(n666) );
  NAND2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n675) );
  AND2_X1 U730 ( .A1(KEYINPUT86), .A2(n671), .ZN(n668) );
  AND2_X1 U731 ( .A1(n756), .A2(n668), .ZN(n670) );
  NAND2_X1 U732 ( .A1(n669), .A2(n670), .ZN(n674) );
  INV_X1 U733 ( .A(KEYINPUT2), .ZN(n672) );
  OR2_X1 U734 ( .A1(n487), .A2(n672), .ZN(n673) );
  NAND2_X1 U735 ( .A1(n675), .A2(n352), .ZN(n678) );
  NAND2_X1 U736 ( .A1(n359), .A2(KEYINPUT2), .ZN(n677) );
  NAND2_X1 U737 ( .A1(n712), .A2(G469), .ZN(n684) );
  XOR2_X1 U738 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n680) );
  XNOR2_X1 U739 ( .A(KEYINPUT124), .B(KEYINPUT123), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U741 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U742 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X2 U743 ( .A1(n685), .A2(n718), .ZN(n687) );
  INV_X1 U744 ( .A(KEYINPUT125), .ZN(n686) );
  XNOR2_X1 U745 ( .A(n687), .B(n686), .ZN(G54) );
  XNOR2_X1 U746 ( .A(n688), .B(G140), .ZN(G42) );
  XOR2_X1 U747 ( .A(G110), .B(n689), .Z(G12) );
  XNOR2_X1 U748 ( .A(G119), .B(KEYINPUT127), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n691), .B(G122), .ZN(G24) );
  NAND2_X1 U750 ( .A1(n361), .A2(G217), .ZN(n694) );
  XNOR2_X1 U751 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X2 U752 ( .A1(n695), .A2(n718), .ZN(n696) );
  XNOR2_X1 U753 ( .A(n696), .B(KEYINPUT126), .ZN(G66) );
  NAND2_X1 U754 ( .A1(n712), .A2(G472), .ZN(n700) );
  XNOR2_X1 U755 ( .A(KEYINPUT93), .B(KEYINPUT62), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X2 U757 ( .A1(n701), .A2(n718), .ZN(n703) );
  XNOR2_X1 U758 ( .A(KEYINPUT91), .B(KEYINPUT63), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n703), .B(n702), .ZN(G57) );
  NAND2_X1 U760 ( .A1(n361), .A2(G478), .ZN(n704) );
  XOR2_X1 U761 ( .A(n705), .B(n704), .Z(n706) );
  NOR2_X1 U762 ( .A1(n706), .A2(n718), .ZN(G63) );
  NAND2_X1 U763 ( .A1(n361), .A2(G475), .ZN(n709) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X2 U765 ( .A1(n710), .A2(n718), .ZN(n711) );
  XNOR2_X1 U766 ( .A(n711), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U767 ( .A1(n712), .A2(G210), .ZN(n717) );
  XOR2_X1 U768 ( .A(KEYINPUT92), .B(KEYINPUT54), .Z(n713) );
  XNOR2_X1 U769 ( .A(n713), .B(KEYINPUT55), .ZN(n714) );
  XNOR2_X1 U770 ( .A(n369), .B(n714), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(n719) );
  NOR2_X2 U772 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n720), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U774 ( .A(G101), .B(n721), .ZN(G3) );
  NOR2_X1 U775 ( .A1(n735), .A2(n724), .ZN(n722) );
  XOR2_X1 U776 ( .A(KEYINPUT116), .B(n722), .Z(n723) );
  XNOR2_X1 U777 ( .A(G104), .B(n723), .ZN(G6) );
  NOR2_X1 U778 ( .A1(n724), .A2(n738), .ZN(n728) );
  XOR2_X1 U779 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n726) );
  XNOR2_X1 U780 ( .A(G107), .B(KEYINPUT117), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U782 ( .A(n728), .B(n727), .ZN(G9) );
  NOR2_X1 U783 ( .A1(n732), .A2(n738), .ZN(n730) );
  XNOR2_X1 U784 ( .A(KEYINPUT118), .B(KEYINPUT29), .ZN(n729) );
  XNOR2_X1 U785 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U786 ( .A(G128), .B(n731), .ZN(G30) );
  NOR2_X1 U787 ( .A1(n732), .A2(n735), .ZN(n734) );
  XNOR2_X1 U788 ( .A(G146), .B(KEYINPUT119), .ZN(n733) );
  XNOR2_X1 U789 ( .A(n734), .B(n733), .ZN(G48) );
  NOR2_X1 U790 ( .A1(n735), .A2(n737), .ZN(n736) );
  XOR2_X1 U791 ( .A(G113), .B(n736), .Z(G15) );
  NOR2_X1 U792 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U793 ( .A(G116), .B(n739), .Z(G18) );
  XNOR2_X1 U794 ( .A(G125), .B(n740), .ZN(n741) );
  XNOR2_X1 U795 ( .A(n741), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U796 ( .A(G134), .B(n742), .ZN(G36) );
  NOR2_X1 U797 ( .A1(n743), .A2(G953), .ZN(n748) );
  INV_X1 U798 ( .A(G898), .ZN(n746) );
  NAND2_X1 U799 ( .A1(G953), .A2(G224), .ZN(n744) );
  XOR2_X1 U800 ( .A(KEYINPUT61), .B(n744), .Z(n745) );
  NOR2_X1 U801 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U802 ( .A1(n748), .A2(n747), .ZN(n755) );
  XOR2_X1 U803 ( .A(G101), .B(n749), .Z(n750) );
  XNOR2_X1 U804 ( .A(n751), .B(n750), .ZN(n753) );
  NOR2_X1 U805 ( .A1(G898), .A2(n763), .ZN(n752) );
  NOR2_X1 U806 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U807 ( .A(n755), .B(n754), .Z(G69) );
  NAND2_X1 U808 ( .A1(n756), .A2(n757), .ZN(n762) );
  XNOR2_X1 U809 ( .A(n758), .B(n759), .ZN(n760) );
  XOR2_X1 U810 ( .A(n761), .B(n760), .Z(n765) );
  XNOR2_X1 U811 ( .A(n762), .B(n765), .ZN(n764) );
  NAND2_X1 U812 ( .A1(n764), .A2(n763), .ZN(n769) );
  XNOR2_X1 U813 ( .A(G227), .B(n765), .ZN(n766) );
  NAND2_X1 U814 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U815 ( .A1(n767), .A2(G953), .ZN(n768) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(G72) );
  XOR2_X1 U817 ( .A(n770), .B(G143), .Z(G45) );
  XNOR2_X1 U818 ( .A(G137), .B(n771), .ZN(G39) );
  XNOR2_X1 U819 ( .A(G131), .B(n772), .ZN(G33) );
endmodule

