//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT35), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT23), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n207), .A2(new_n209), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n214), .A2(new_n215), .A3(new_n210), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n204), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n207), .A2(new_n209), .ZN(new_n218));
  INV_X1    g017(.A(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT24), .A3(new_n220), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n214), .A2(new_n210), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n218), .A2(new_n221), .A3(KEYINPUT25), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT27), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G183gat), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(G183gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT65), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT28), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(G190gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n230), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n231), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n234), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n205), .A3(new_n206), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n241), .A2(new_n205), .A3(new_n206), .A4(KEYINPUT66), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n212), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n205), .A2(new_n206), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(KEYINPUT26), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n214), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n224), .A2(KEYINPUT64), .B1(new_n240), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n217), .A2(new_n223), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT71), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n250), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n253), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT29), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(new_n255), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n224), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n256), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n257), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT70), .B(G218gat), .Z(new_n270));
  AOI21_X1  g069(.A(KEYINPUT22), .B1(new_n270), .B2(G211gat), .ZN(new_n271));
  XOR2_X1   g070(.A(G197gat), .B(G204gat), .Z(new_n272));
  OAI21_X1  g071(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT22), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT70), .B(G218gat), .ZN(new_n275));
  INV_X1    g074(.A(G211gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n272), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n268), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n267), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n251), .A2(new_n256), .A3(new_n253), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n261), .A3(new_n255), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(G36gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT72), .B(G8gat), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n285), .B1(new_n267), .B2(new_n281), .ZN(new_n293));
  INV_X1    g092(.A(new_n291), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(KEYINPUT30), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n282), .A2(new_n286), .A3(new_n294), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n293), .A2(new_n299), .A3(new_n294), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT74), .B(KEYINPUT30), .Z(new_n302));
  AOI21_X1  g101(.A(new_n296), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G228gat), .ZN(new_n304));
  INV_X1    g103(.A(G233gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G141gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n313), .B2(G148gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317));
  NOR2_X1   g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n307), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(G148gat), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n309), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n318), .A2(new_n317), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n315), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(KEYINPUT77), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G141gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G148gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT2), .B1(new_n309), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G155gat), .B(G162gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT75), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n318), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n334));
  XNOR2_X1  g133(.A(G141gat), .B(G148gat), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(KEYINPUT2), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n320), .A2(new_n327), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n279), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n268), .B1(new_n277), .B2(new_n278), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n261), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n332), .A2(new_n336), .ZN(new_n343));
  AOI221_X4 g142(.A(new_n307), .B1(new_n325), .B2(new_n315), .C1(new_n323), .C2(new_n309), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT77), .B1(new_n324), .B2(new_n326), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n341), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n280), .B1(new_n346), .B2(new_n261), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n306), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G218gat), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n349), .A2(KEYINPUT70), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(KEYINPUT70), .ZN(new_n351));
  OAI21_X1  g150(.A(G211gat), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n272), .B1(new_n352), .B2(new_n274), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT86), .B1(new_n353), .B2(new_n268), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT85), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n279), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n357), .B(new_n269), .C1(new_n271), .C2(new_n272), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT85), .A4(new_n268), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n354), .A2(new_n356), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n261), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n337), .B1(new_n361), .B2(new_n341), .ZN(new_n362));
  INV_X1    g161(.A(new_n306), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n337), .B2(new_n341), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n280), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n348), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G22gat), .ZN(new_n367));
  INV_X1    g166(.A(G22gat), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n348), .B(new_n368), .C1(new_n362), .C2(new_n365), .ZN(new_n369));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT31), .ZN(new_n371));
  INV_X1    g170(.A(G50gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n367), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n375), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n367), .A2(new_n369), .ZN(new_n378));
  INV_X1    g177(.A(new_n373), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT88), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381));
  AOI211_X1 g180(.A(new_n381), .B(new_n373), .C1(new_n367), .C2(new_n369), .ZN(new_n382));
  OAI22_X1  g181(.A1(new_n376), .A2(new_n377), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G113gat), .B(G120gat), .Z(new_n384));
  INV_X1    g183(.A(KEYINPUT1), .ZN(new_n385));
  AND2_X1   g184(.A1(G127gat), .A2(G134gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(G127gat), .A2(G134gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n384), .B(new_n385), .C1(KEYINPUT67), .C2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G113gat), .ZN(new_n390));
  INV_X1    g189(.A(G120gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G113gat), .A2(G120gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n385), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(KEYINPUT67), .A3(new_n393), .ZN(new_n395));
  XNOR2_X1  g194(.A(G127gat), .B(G134gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n260), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n398), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n251), .A2(new_n400), .A3(new_n253), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n399), .A2(G227gat), .A3(new_n401), .A4(G233gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(KEYINPUT32), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT32), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n407), .A3(new_n403), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G15gat), .B(G43gat), .Z(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n413), .B1(new_n411), .B2(new_n416), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n409), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n411), .A2(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n412), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n422), .A2(new_n408), .A3(new_n406), .A4(new_n417), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n303), .A2(new_n383), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G57gat), .ZN(new_n428));
  INV_X1    g227(.A(G85gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT5), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n398), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT82), .B1(new_n433), .B2(KEYINPUT4), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n337), .A2(new_n435), .A3(new_n436), .A4(new_n398), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n433), .A2(new_n440), .A3(KEYINPUT4), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n433), .B2(KEYINPUT4), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n432), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(G225gat), .A2(G233gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT78), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n389), .A2(new_n397), .A3(KEYINPUT78), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n337), .B2(new_n341), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT79), .ZN(new_n453));
  INV_X1    g252(.A(new_n346), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n456), .A2(KEYINPUT3), .B1(new_n450), .B2(new_n449), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT79), .B1(new_n457), .B2(new_n346), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n445), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n444), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n449), .A2(new_n450), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n433), .B1(new_n461), .B2(new_n337), .ZN(new_n462));
  INV_X1    g261(.A(new_n445), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT5), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n453), .B1(new_n452), .B2(new_n454), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n457), .A2(KEYINPUT79), .A3(new_n346), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n433), .A2(KEYINPUT4), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT80), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n337), .A2(KEYINPUT81), .A3(new_n436), .A4(new_n398), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT81), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n433), .B2(KEYINPUT4), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT80), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n433), .A2(new_n474), .A3(KEYINPUT4), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n470), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n465), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT6), .B(new_n431), .C1(new_n460), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n479));
  INV_X1    g278(.A(new_n465), .ZN(new_n480));
  INV_X1    g279(.A(new_n476), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n459), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n441), .A2(new_n442), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT5), .B1(new_n483), .B2(new_n438), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n468), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT6), .A4(new_n431), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n468), .A2(new_n476), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n489), .A2(new_n480), .B1(new_n484), .B2(new_n468), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT6), .B1(new_n490), .B2(new_n430), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n431), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n479), .A2(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n203), .B1(new_n425), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n420), .A2(new_n423), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n378), .A2(new_n379), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n381), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n378), .A2(KEYINPUT88), .A3(new_n379), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n374), .B(new_n375), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n479), .A2(new_n488), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n491), .A2(new_n492), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n501), .A2(KEYINPUT35), .A3(new_n504), .A4(new_n303), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n494), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n283), .A2(new_n284), .A3(new_n281), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n507), .A2(KEYINPUT37), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n267), .B2(new_n281), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n293), .B2(KEYINPUT37), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n294), .A2(KEYINPUT38), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n298), .A2(new_n300), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n502), .A2(new_n512), .A3(new_n503), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n493), .A2(KEYINPUT90), .A3(new_n512), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT38), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n293), .B(KEYINPUT37), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n291), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT40), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n483), .A2(new_n438), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n466), .A2(new_n467), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n445), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT39), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n445), .B(new_n433), .C1(new_n461), .C2(new_n337), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT39), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n430), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n522), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n525), .A2(new_n532), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n535), .A2(KEYINPUT40), .A3(new_n430), .A4(new_n527), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n536), .A3(new_n492), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n383), .B1(new_n537), .B2(new_n303), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n383), .ZN(new_n541));
  INV_X1    g340(.A(new_n300), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n299), .B1(new_n293), .B2(new_n294), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n302), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n296), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n541), .B1(new_n493), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n424), .B2(KEYINPUT36), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n495), .A2(KEYINPUT69), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n424), .A2(KEYINPUT36), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n506), .B1(new_n540), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n372), .A2(G43gat), .ZN(new_n557));
  INV_X1    g356(.A(G43gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G50gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT94), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(KEYINPUT15), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n372), .A2(KEYINPUT95), .A3(G43gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n559), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT15), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G29gat), .ZN(new_n571));
  INV_X1    g370(.A(G36gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT14), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT14), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(G29gat), .B2(G36gat), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n573), .B(new_n575), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n564), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n564), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT17), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT96), .ZN(new_n581));
  XNOR2_X1  g380(.A(G15gat), .B(G22gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT16), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(G1gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(G1gat), .B2(new_n582), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(G8gat), .Z(new_n586));
  OR2_X1    g385(.A1(new_n579), .A2(KEYINPUT17), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n581), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n586), .A2(new_n579), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT97), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(KEYINPUT18), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n586), .A2(new_n579), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n592), .B(KEYINPUT13), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(new_n592), .A3(new_n590), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT18), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT93), .ZN(new_n602));
  XOR2_X1   g401(.A(G113gat), .B(G141gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT92), .ZN(new_n604));
  XOR2_X1   g403(.A(G169gat), .B(G197gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n601), .A2(KEYINPUT93), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n202), .B1(new_n556), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n519), .B1(new_n513), .B2(new_n514), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n538), .B1(new_n616), .B2(new_n516), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(new_n554), .ZN(new_n618));
  OAI211_X1 g417(.A(KEYINPUT98), .B(new_n613), .C1(new_n618), .C2(new_n506), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621));
  INV_X1    g420(.A(G92gat), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n621), .B1(new_n429), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(KEYINPUT7), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT7), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n621), .B(new_n626), .C1(new_n429), .C2(new_n622), .ZN(new_n627));
  NAND2_X1  g426(.A1(G99gat), .A2(G106gat), .ZN(new_n628));
  AOI22_X1  g427(.A1(KEYINPUT8), .A2(new_n628), .B1(new_n429), .B2(new_n622), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G99gat), .ZN(new_n631));
  INV_X1    g430(.A(G106gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n630), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n628), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n625), .A2(new_n635), .A3(new_n627), .A4(new_n629), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n581), .A2(new_n587), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n579), .A2(new_n637), .ZN(new_n640));
  AND2_X1   g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(KEYINPUT41), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OR3_X1    g442(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n645));
  XNOR2_X1  g444(.A(G190gat), .B(G218gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n639), .B1(new_n638), .B2(new_n643), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n644), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n644), .B2(new_n648), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT21), .ZN(new_n653));
  XOR2_X1   g452(.A(G57gat), .B(G64gat), .Z(new_n654));
  AOI21_X1  g453(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G71gat), .B(G78gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n586), .B1(new_n653), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n228), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n662));
  NAND2_X1  g461(.A1(G231gat), .A2(G233gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n661), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n653), .ZN(new_n666));
  XOR2_X1   g465(.A(G127gat), .B(G155gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n276), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n669), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(G230gat), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n305), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n637), .B(new_n659), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(KEYINPUT10), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n637), .A2(new_n659), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT10), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n676), .B2(new_n675), .ZN(new_n681));
  XNOR2_X1  g480(.A(G120gat), .B(G148gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G176gat), .ZN(new_n683));
  INV_X1    g482(.A(G204gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n652), .A2(new_n673), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n620), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n493), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g492(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n546), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT16), .B(G8gat), .Z(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT102), .Z(new_n697));
  OAI21_X1  g496(.A(new_n694), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(G8gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(KEYINPUT42), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n698), .B(new_n699), .C1(new_n695), .C2(new_n700), .ZN(G1325gat));
  NAND3_X1  g500(.A1(new_n620), .A2(new_n424), .A3(new_n689), .ZN(new_n702));
  INV_X1    g501(.A(G15gat), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n702), .A2(KEYINPUT103), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT103), .B1(new_n702), .B2(new_n703), .ZN(new_n705));
  INV_X1    g504(.A(new_n553), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  OAI22_X1  g506(.A1(new_n704), .A2(new_n705), .B1(new_n690), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1326gat));
  NOR2_X1   g509(.A1(new_n690), .A2(new_n383), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NOR2_X1   g512(.A1(new_n672), .A2(new_n688), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n620), .A2(new_n652), .A3(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G29gat), .A3(new_n504), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT45), .Z(new_n717));
  NAND2_X1  g516(.A1(new_n613), .A2(new_n714), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n540), .A2(new_n555), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT105), .B1(new_n617), .B2(new_n554), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n506), .A2(KEYINPUT106), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n494), .A2(new_n505), .A3(new_n723), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n651), .A2(KEYINPUT44), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT107), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n722), .A2(new_n724), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n719), .B1(new_n540), .B2(new_n555), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n617), .A2(KEYINPUT105), .A3(new_n554), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n726), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT44), .B1(new_n556), .B2(new_n651), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n718), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n504), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n717), .A2(new_n739), .ZN(G1328gat));
  NAND2_X1  g539(.A1(new_n546), .A2(new_n572), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n715), .A2(KEYINPUT108), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n715), .B2(new_n741), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n742), .B(new_n743), .C1(KEYINPUT109), .C2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(KEYINPUT46), .ZN(new_n747));
  OAI21_X1  g546(.A(G36gat), .B1(new_n738), .B2(new_n303), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n742), .A2(KEYINPUT109), .A3(new_n744), .A4(new_n743), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(G1329gat));
  NAND2_X1  g549(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n558), .B1(new_n737), .B2(new_n706), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n424), .A2(new_n558), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n715), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n751), .B(new_n754), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n725), .A2(KEYINPUT107), .A3(new_n727), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n733), .B1(new_n732), .B2(new_n726), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n736), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n718), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(new_n706), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G43gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n757), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n764), .A2(new_n752), .A3(new_n753), .A4(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n758), .A2(new_n766), .ZN(G1330gat));
  AOI21_X1  g566(.A(new_n372), .B1(new_n737), .B2(new_n541), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT48), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n715), .A2(G50gat), .A3(new_n383), .ZN(new_n770));
  OR3_X1    g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1331gat));
  NAND3_X1  g572(.A1(new_n651), .A2(new_n672), .A3(new_n688), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n725), .A2(new_n613), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n493), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g576(.A(new_n303), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT111), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n780), .B(new_n781), .Z(G1333gat));
  NAND2_X1  g581(.A1(new_n775), .A2(new_n706), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n495), .A2(G71gat), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n783), .A2(G71gat), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n775), .A2(new_n541), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g587(.A1(new_n613), .A2(new_n672), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n688), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n735), .B2(new_n736), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n493), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n652), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n725), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT51), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n493), .A2(new_n429), .A3(new_n688), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT112), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n792), .A2(new_n429), .B1(new_n796), .B2(new_n798), .ZN(G1336gat));
  NAND4_X1  g598(.A1(new_n795), .A2(new_n622), .A3(new_n546), .A4(new_n688), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n622), .B1(new_n791), .B2(new_n546), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n791), .A2(new_n546), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n804), .B(new_n800), .C1(new_n805), .C2(new_n622), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(G1337gat));
  AND2_X1   g606(.A1(new_n791), .A2(new_n706), .ZN(new_n808));
  OAI21_X1  g607(.A(G99gat), .B1(new_n808), .B2(KEYINPUT113), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n791), .A2(KEYINPUT113), .A3(new_n706), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n688), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n424), .A2(new_n631), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(G1338gat));
  NAND4_X1  g612(.A1(new_n795), .A2(new_n632), .A3(new_n541), .A4(new_n688), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n632), .B1(new_n791), .B2(new_n541), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT53), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n791), .A2(new_n541), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n818), .B(new_n814), .C1(new_n819), .C2(new_n632), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(G1339gat));
  NAND2_X1  g620(.A1(new_n689), .A2(new_n614), .ZN(new_n822));
  INV_X1    g621(.A(new_n680), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n677), .A2(new_n679), .A3(new_n675), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(KEYINPUT54), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n685), .B1(new_n680), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(KEYINPUT55), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n687), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT55), .B1(new_n825), .B2(new_n827), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n828), .A2(KEYINPUT114), .A3(new_n687), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n831), .A2(new_n834), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n593), .A2(new_n597), .A3(new_n600), .A4(new_n609), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n591), .A2(new_n592), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n595), .A2(new_n596), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n608), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n838), .A2(new_n651), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n688), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n614), .B2(new_n838), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n844), .B1(new_n848), .B2(new_n651), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n822), .B1(new_n849), .B2(new_n672), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n383), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n493), .A2(new_n303), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n495), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n614), .ZN(new_n858));
  INV_X1    g657(.A(new_n822), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n848), .A2(new_n651), .ZN(new_n860));
  INV_X1    g659(.A(new_n844), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n859), .B1(new_n862), .B2(new_n673), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n504), .A3(new_n425), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT117), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n390), .A3(new_n613), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n858), .A2(new_n866), .ZN(G1340gat));
  OAI21_X1  g666(.A(G120gat), .B1(new_n857), .B2(new_n845), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n391), .A3(new_n688), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1341gat));
  NAND4_X1  g669(.A1(new_n854), .A2(G127gat), .A3(new_n672), .A4(new_n856), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g672(.A(G127gat), .B1(new_n864), .B2(new_n672), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1342gat));
  INV_X1    g674(.A(G134gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n864), .A2(new_n876), .A3(new_n652), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n854), .A2(new_n652), .A3(new_n856), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n883), .A2(new_n884), .A3(G134gat), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n883), .B2(G134gat), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n880), .B(new_n882), .C1(new_n885), .C2(new_n886), .ZN(G1343gat));
  NOR2_X1   g686(.A1(new_n706), .A2(new_n383), .ZN(new_n888));
  AND4_X1   g687(.A1(new_n493), .A2(new_n850), .A3(new_n303), .A4(new_n888), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n889), .A2(new_n328), .A3(new_n613), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(KEYINPUT58), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n833), .A2(new_n687), .A3(new_n828), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n610), .B2(new_n612), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n651), .B1(new_n894), .B2(new_n846), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT122), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n861), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n895), .A2(KEYINPUT122), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n673), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n822), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n892), .B1(new_n900), .B2(new_n541), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n383), .A2(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n850), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n706), .A2(new_n855), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT121), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n901), .A2(new_n614), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n891), .B1(new_n907), .B2(new_n313), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n909), .B1(new_n901), .B2(new_n906), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n844), .B1(new_n895), .B2(KEYINPUT122), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(KEYINPUT122), .B2(new_n895), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n859), .B1(new_n912), .B2(new_n673), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT57), .B1(new_n913), .B2(new_n383), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n914), .A2(KEYINPUT123), .A3(new_n903), .A4(new_n905), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n915), .A3(new_n613), .ZN(new_n916));
  INV_X1    g715(.A(new_n313), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n890), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n908), .B1(new_n918), .B2(new_n919), .ZN(G1344gat));
  NAND3_X1  g719(.A1(new_n910), .A2(new_n915), .A3(new_n688), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n308), .A2(KEYINPUT59), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924));
  INV_X1    g723(.A(new_n893), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n613), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n652), .B1(new_n926), .B2(new_n847), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n927), .B2(new_n844), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n861), .A2(KEYINPUT124), .A3(new_n895), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n929), .A3(new_n673), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n822), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n850), .A2(new_n541), .ZN(new_n932));
  AOI22_X1  g731(.A1(new_n902), .A2(new_n931), .B1(new_n932), .B2(KEYINPUT57), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n933), .A2(new_n688), .A3(new_n905), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT59), .B1(new_n934), .B2(new_n308), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n923), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n889), .A2(new_n308), .A3(new_n688), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1345gat));
  AOI21_X1  g737(.A(G155gat), .B1(new_n889), .B2(new_n672), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n910), .A2(new_n915), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n672), .A2(G155gat), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT125), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(G1346gat));
  NAND3_X1  g742(.A1(new_n910), .A2(new_n915), .A3(new_n652), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G162gat), .ZN(new_n945));
  INV_X1    g744(.A(G162gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n889), .A2(new_n946), .A3(new_n652), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1347gat));
  NOR2_X1   g747(.A1(new_n863), .A2(new_n493), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n541), .A2(new_n303), .A3(new_n495), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n613), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n493), .A2(new_n303), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT126), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(new_n495), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n958), .B1(new_n852), .B2(new_n853), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n614), .A2(new_n205), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n953), .B1(new_n959), .B2(new_n960), .ZN(G1348gat));
  NAND3_X1  g760(.A1(new_n952), .A2(new_n206), .A3(new_n688), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n959), .A2(new_n688), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n206), .ZN(G1349gat));
  INV_X1    g763(.A(KEYINPUT60), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n952), .A2(new_n230), .A3(new_n233), .A4(new_n672), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n959), .A2(new_n672), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n965), .B(new_n966), .C1(new_n967), .C2(new_n228), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n228), .B1(new_n959), .B2(new_n672), .ZN(new_n969));
  AND4_X1   g768(.A1(new_n230), .A2(new_n952), .A3(new_n233), .A4(new_n672), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT60), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(G1350gat));
  NAND3_X1  g771(.A1(new_n952), .A2(new_n237), .A3(new_n652), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n652), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(G190gat), .ZN(new_n976));
  AOI211_X1 g775(.A(KEYINPUT61), .B(new_n237), .C1(new_n959), .C2(new_n652), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(G1351gat));
  AND3_X1   g777(.A1(new_n949), .A2(new_n546), .A3(new_n888), .ZN(new_n979));
  AOI21_X1  g778(.A(G197gat), .B1(new_n979), .B2(new_n613), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n956), .A2(new_n706), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n933), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n613), .A2(G197gat), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1352gat));
  NAND3_X1  g783(.A1(new_n979), .A2(new_n684), .A3(new_n688), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n982), .A2(new_n688), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n986), .B(new_n987), .C1(new_n988), .C2(new_n684), .ZN(G1353gat));
  NAND3_X1  g788(.A1(new_n979), .A2(new_n276), .A3(new_n672), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n931), .A2(new_n902), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n932), .A2(KEYINPUT57), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n991), .A2(new_n992), .A3(new_n672), .A4(new_n981), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n276), .B1(new_n993), .B2(KEYINPUT127), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n933), .A2(new_n995), .A3(new_n672), .A4(new_n981), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n994), .A2(KEYINPUT63), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n994), .B2(new_n996), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n990), .B1(new_n997), .B2(new_n998), .ZN(G1354gat));
  AOI21_X1  g798(.A(G218gat), .B1(new_n979), .B2(new_n652), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n651), .A2(new_n275), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n1000), .B1(new_n982), .B2(new_n1001), .ZN(G1355gat));
endmodule


