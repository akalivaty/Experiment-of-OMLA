//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318;
  INV_X1    g0000(.A(KEYINPUT65), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(KEYINPUT64), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n205), .B1(G58), .B2(G68), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  AOI21_X1  g0008(.A(new_n201), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI211_X1 g0009(.A(KEYINPUT65), .B(G50), .C1(new_n204), .C2(new_n206), .ZN(new_n210));
  NOR3_X1   g0010(.A1(new_n209), .A2(new_n210), .A3(G77), .ZN(G353));
  OAI21_X1  g0011(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  NAND2_X1  g0016(.A1(KEYINPUT67), .A2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(KEYINPUT67), .A2(G68), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT66), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G50), .A2(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G116), .ZN(new_n223));
  INV_X1    g0023(.A(G270), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n220), .A2(G238), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n221), .B2(new_n225), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G77), .A2(G244), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n213), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(G20), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n207), .A2(new_n208), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n216), .B(new_n233), .C1(new_n236), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT69), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G50), .B(G68), .Z(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n234), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n235), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n235), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n259), .A2(new_n208), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT67), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n203), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n235), .B1(new_n264), .B2(new_n217), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n257), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT11), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT11), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n268), .B(new_n257), .C1(new_n262), .C2(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT12), .B1(new_n220), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT76), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT76), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n275), .B(KEYINPUT12), .C1(new_n220), .C2(new_n272), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n272), .A2(KEYINPUT12), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n270), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n257), .B1(new_n271), .B2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n203), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G232), .A3(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n286), .A2(new_n288), .A3(G226), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G97), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n285), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G1), .A3(G13), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT73), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT73), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n293), .A2(new_n296), .A3(G1), .A4(G13), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT13), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n294), .A2(new_n301), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(new_n305), .B2(G238), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n299), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n300), .B1(new_n299), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g0108(.A(G200), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n299), .A2(new_n306), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n299), .A2(new_n300), .A3(new_n306), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(G190), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n283), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT77), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT77), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n283), .A2(new_n309), .A3(new_n313), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n307), .A2(new_n308), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(G169), .B1(new_n307), .B2(new_n308), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(KEYINPUT14), .B2(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n321), .A2(KEYINPUT14), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n283), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT8), .B(G58), .Z(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(new_n259), .B1(new_n235), .B2(new_n261), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT15), .B(G87), .Z(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n260), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n257), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n280), .A2(G77), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n334), .C1(G77), .C2(new_n272), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n284), .A2(G1698), .ZN(new_n336));
  INV_X1    g0136(.A(G238), .ZN(new_n337));
  INV_X1    g0137(.A(G107), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n336), .A2(new_n337), .B1(new_n338), .B2(new_n284), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n286), .A2(new_n288), .ZN(new_n340));
  INV_X1    g0140(.A(G232), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n340), .A2(new_n341), .A3(G1698), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n298), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n303), .B1(new_n305), .B2(G244), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n335), .B1(new_n346), .B2(G190), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(G200), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n351), .B(new_n335), .C1(G179), .C2(new_n345), .ZN(new_n352));
  AND4_X1   g0152(.A1(new_n318), .A2(new_n326), .A3(new_n349), .A4(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n340), .A2(new_n289), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(G223), .B1(G77), .B2(new_n340), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n286), .A2(new_n288), .A3(G222), .A4(new_n289), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT71), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT71), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n284), .A2(new_n359), .A3(G222), .A4(new_n289), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n356), .A2(KEYINPUT72), .A3(new_n361), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n298), .ZN(new_n366));
  INV_X1    g0166(.A(G41), .ZN(new_n367));
  INV_X1    g0167(.A(G45), .ZN(new_n368));
  AOI21_X1  g0168(.A(G1), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G274), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT70), .B(G226), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n304), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n354), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n366), .A2(new_n354), .A3(new_n373), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(G200), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n366), .A2(new_n354), .A3(new_n373), .ZN(new_n378));
  OAI21_X1  g0178(.A(G190), .B1(new_n378), .B2(new_n374), .ZN(new_n379));
  INV_X1    g0179(.A(new_n257), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n209), .B2(new_n210), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n258), .A2(G20), .ZN(new_n382));
  NOR2_X1   g0182(.A1(G20), .A2(G33), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n327), .A2(new_n382), .B1(G150), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n380), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n280), .A2(G50), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G50), .B2(new_n272), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g0188(.A(new_n388), .B(KEYINPUT9), .Z(new_n389));
  NAND3_X1  g0189(.A1(new_n377), .A2(new_n379), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT10), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT10), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n377), .A2(new_n379), .A3(new_n389), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n218), .A2(new_n219), .A3(new_n202), .ZN(new_n396));
  OAI21_X1  g0196(.A(G20), .B1(new_n396), .B2(new_n207), .ZN(new_n397));
  INV_X1    g0197(.A(G159), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT78), .B1(new_n259), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT78), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n383), .A2(new_n400), .A3(G159), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n220), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n284), .B2(G20), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n340), .A2(KEYINPUT7), .A3(new_n235), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n395), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT7), .B1(new_n340), .B2(new_n235), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n405), .B(G20), .C1(new_n286), .C2(new_n288), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n264), .A2(G58), .A3(new_n217), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n206), .A3(new_n204), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(G20), .B1(new_n399), .B2(new_n401), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n415), .A3(KEYINPUT16), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n409), .A2(new_n416), .A3(new_n257), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n328), .A2(new_n272), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n280), .B2(new_n328), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n370), .B1(new_n304), .B2(new_n341), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n286), .A2(new_n288), .A3(G226), .A4(G1698), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n286), .A2(new_n288), .A3(G223), .A4(new_n289), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n421), .B1(new_n298), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G179), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n350), .B2(new_n426), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n420), .A2(KEYINPUT18), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT18), .B1(new_n420), .B2(new_n428), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(new_n298), .ZN(new_n432));
  INV_X1    g0232(.A(new_n421), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G200), .B2(new_n426), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n417), .A2(new_n419), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT17), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n417), .A2(new_n439), .A3(new_n419), .A4(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n431), .A2(KEYINPUT79), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT79), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n429), .A2(new_n430), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n438), .A2(new_n440), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n353), .A2(new_n394), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n375), .A2(new_n376), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n319), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n375), .A2(new_n376), .A3(new_n350), .ZN(new_n451));
  INV_X1    g0251(.A(new_n388), .ZN(new_n452));
  AND4_X1   g0252(.A1(KEYINPUT75), .A2(new_n450), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n388), .B1(new_n449), .B2(new_n319), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT75), .B1(new_n454), .B2(new_n451), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n272), .ZN(new_n458));
  INV_X1    g0258(.A(G97), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n380), .B(new_n272), .C1(G1), .C2(new_n258), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(new_n459), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(G107), .B1(new_n410), .B2(new_n411), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(KEYINPUT80), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT80), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G97), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT6), .A4(new_n338), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT6), .ZN(new_n469));
  AND2_X1   g0269(.A1(G97), .A2(G107), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G97), .A2(G107), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(G20), .B1(G77), .B2(new_n383), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n464), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n463), .B1(new_n475), .B2(new_n380), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n271), .B(G45), .C1(new_n367), .C2(KEYINPUT5), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n367), .A2(KEYINPUT5), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G274), .ZN(new_n480));
  OAI211_X1 g0280(.A(G257), .B(new_n294), .C1(new_n477), .C2(new_n478), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n286), .A2(new_n288), .A3(G244), .A4(new_n289), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n289), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n482), .B1(new_n489), .B2(new_n298), .ZN(new_n490));
  INV_X1    g0290(.A(G200), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI211_X1 g0292(.A(new_n434), .B(new_n482), .C1(new_n489), .C2(new_n298), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n476), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n298), .ZN(new_n495));
  INV_X1    g0295(.A(new_n482), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n380), .B1(new_n464), .B2(new_n474), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n497), .A2(G179), .B1(new_n498), .B2(new_n462), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n490), .A2(G169), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT81), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n350), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n490), .A2(new_n319), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n476), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n494), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n258), .A2(new_n223), .A3(G20), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n235), .B2(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n338), .A2(KEYINPUT23), .A3(G20), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(KEYINPUT84), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(new_n286), .A3(new_n288), .A4(new_n235), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n284), .A2(KEYINPUT22), .A3(new_n235), .A4(new_n513), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n511), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT24), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n511), .A2(new_n516), .A3(KEYINPUT24), .A4(new_n517), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n257), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n461), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT25), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n272), .B2(G107), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n458), .A2(KEYINPUT25), .A3(new_n338), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n523), .A2(G107), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n286), .A2(new_n288), .A3(G250), .A4(new_n289), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n286), .A2(new_n288), .A3(G257), .A4(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n298), .ZN(new_n533));
  OAI211_X1 g0333(.A(G264), .B(new_n294), .C1(new_n477), .C2(new_n478), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n480), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n491), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT85), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n533), .A2(new_n480), .A3(new_n534), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n434), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(KEYINPUT85), .A3(new_n491), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n528), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n330), .A2(new_n272), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n461), .A2(new_n331), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n235), .B1(new_n291), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n465), .A2(new_n467), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n512), .A2(new_n338), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n544), .B(new_n546), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n286), .A2(new_n288), .A3(new_n235), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n382), .A2(new_n465), .A3(new_n467), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n551), .A2(G68), .B1(new_n552), .B2(new_n545), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n549), .B1(new_n465), .B2(new_n467), .ZN(new_n554));
  INV_X1    g0354(.A(new_n546), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT82), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n550), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n542), .B(new_n543), .C1(new_n557), .C2(new_n257), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n234), .B1(G33), .B2(G41), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n271), .A2(G45), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G250), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n559), .A2(new_n561), .B1(new_n302), .B2(new_n560), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n286), .A2(new_n288), .A3(G244), .A4(G1698), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n286), .A2(new_n288), .A3(G238), .A4(new_n289), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n564), .C1(new_n258), .C2(new_n223), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n562), .B1(new_n565), .B2(new_n298), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n319), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(G169), .B2(new_n566), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n557), .A2(new_n257), .ZN(new_n569));
  INV_X1    g0369(.A(new_n542), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n523), .A2(G87), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n565), .A2(new_n298), .ZN(new_n573));
  INV_X1    g0373(.A(new_n562), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(G190), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n491), .B2(new_n566), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n558), .A2(new_n568), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n541), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n284), .A2(G257), .A3(new_n289), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n340), .A2(G303), .ZN(new_n581));
  INV_X1    g0381(.A(G264), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n581), .C1(new_n336), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n298), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n479), .A2(new_n559), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(G270), .B1(G274), .B2(new_n479), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n350), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n458), .A2(new_n223), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n461), .B2(new_n223), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n235), .B(new_n487), .C1(new_n547), .C2(G33), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT83), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n223), .A2(G20), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n257), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n257), .B2(new_n593), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n591), .B(KEYINPUT20), .C1(new_n594), .C2(new_n595), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n590), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n579), .B1(new_n588), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n600), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(KEYINPUT21), .A3(new_n587), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n538), .A2(new_n319), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n535), .A2(new_n350), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n528), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n584), .A2(new_n586), .A3(G179), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n601), .A2(new_n603), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n584), .A2(new_n586), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G200), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n434), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n602), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n457), .A2(new_n506), .A3(new_n578), .A4(new_n614), .ZN(G372));
  NAND3_X1  g0415(.A1(new_n506), .A2(new_n578), .A3(new_n609), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n501), .A2(new_n505), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT26), .B1(new_n617), .B2(new_n577), .ZN(new_n618));
  INV_X1    g0418(.A(new_n558), .ZN(new_n619));
  INV_X1    g0419(.A(new_n568), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n577), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n476), .A2(new_n502), .A3(new_n504), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n616), .A2(new_n618), .A3(new_n621), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n457), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n352), .B1(new_n315), .B2(new_n317), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n283), .B1(new_n322), .B2(new_n323), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n441), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n431), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n391), .A2(new_n393), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n456), .B(new_n629), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n632), .A2(new_n431), .B1(new_n391), .B2(new_n393), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT75), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n454), .A2(KEYINPUT75), .A3(new_n451), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT86), .B1(new_n636), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n628), .A2(new_n643), .ZN(G369));
  OAI211_X1 g0444(.A(new_n611), .B(new_n600), .C1(new_n434), .C2(new_n610), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n601), .A2(new_n603), .A3(new_n645), .A4(new_n608), .ZN(new_n646));
  INV_X1    g0446(.A(G13), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(G20), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT27), .B1(new_n649), .B2(G1), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n651), .A3(new_n271), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n650), .A2(G213), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G343), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT87), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT88), .B1(new_n655), .B2(new_n602), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n646), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n646), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n657), .A2(KEYINPUT89), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT89), .B1(new_n657), .B2(new_n658), .ZN(new_n660));
  INV_X1    g0460(.A(G330), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT91), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n655), .A2(new_n528), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT90), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n541), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n655), .A2(new_n528), .A3(KEYINPUT90), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(new_n606), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n655), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n606), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n663), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  AOI211_X1 g0473(.A(KEYINPUT91), .B(new_n671), .C1(new_n666), .C2(new_n668), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n662), .A2(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n601), .A2(new_n603), .A3(new_n608), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n655), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n667), .A2(new_n606), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n535), .A2(KEYINPUT85), .A3(new_n491), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT85), .B1(new_n535), .B2(new_n491), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n535), .A2(G190), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT90), .B1(new_n685), .B2(new_n528), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n681), .B1(new_n686), .B2(new_n664), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT91), .B1(new_n687), .B2(new_n671), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n669), .A2(new_n663), .A3(new_n672), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n680), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n606), .A2(new_n655), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n677), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT92), .ZN(G399));
  NAND2_X1  g0494(.A1(new_n554), .A2(new_n223), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n214), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(G1), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n237), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT26), .B1(new_n577), .B2(new_n624), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n622), .A2(new_n501), .A3(new_n623), .A4(new_n505), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n616), .A2(new_n704), .A3(new_n621), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT29), .A3(new_n670), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT29), .B1(new_n627), .B2(new_n670), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n497), .A2(new_n610), .A3(new_n319), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n566), .A2(new_n713), .A3(new_n533), .A4(new_n534), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n573), .A2(new_n574), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n533), .A2(new_n534), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT93), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n712), .A2(KEYINPUT30), .A3(new_n714), .A4(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n607), .A3(new_n490), .A4(new_n714), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n538), .A2(new_n490), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(new_n319), .A3(new_n715), .A4(new_n610), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT31), .B1(new_n724), .B2(new_n655), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n614), .A2(new_n506), .A3(new_n578), .A4(new_n670), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n661), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n711), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n703), .B1(new_n732), .B2(G1), .ZN(G364));
  AOI21_X1  g0533(.A(new_n271), .B1(new_n648), .B2(G45), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n699), .A2(KEYINPUT94), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT94), .ZN(new_n736));
  INV_X1    g0536(.A(new_n734), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n736), .B1(new_n698), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n662), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n661), .B1(new_n659), .B2(new_n660), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n657), .A2(new_n658), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n434), .A2(G20), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT99), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n751), .A2(G179), .A3(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G159), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT32), .Z(new_n754));
  NOR2_X1   g0554(.A1(new_n434), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n319), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n459), .ZN(new_n759));
  NOR4_X1   g0559(.A1(new_n235), .A2(new_n434), .A3(new_n491), .A4(G179), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n284), .B1(new_n761), .B2(new_n512), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n235), .A2(new_n319), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n434), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n759), .B(new_n762), .C1(G68), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT98), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n754), .B(new_n766), .C1(new_n208), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n751), .A2(G179), .A3(new_n491), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n338), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n763), .A2(KEYINPUT97), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT97), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n235), .B2(new_n319), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n777), .A2(new_n779), .A3(new_n755), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n776), .B1(G58), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G190), .A2(G200), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n777), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n261), .B2(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n752), .A2(G329), .B1(new_n781), .B2(G322), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(new_n787), .B2(new_n775), .C1(new_n788), .C2(new_n784), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n340), .B1(new_n761), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G294), .B2(new_n757), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n771), .A2(G326), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT33), .B(G317), .Z(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n793), .C1(new_n764), .C2(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n773), .A2(new_n785), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n234), .B1(G20), .B2(new_n350), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n697), .A2(new_n340), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT95), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G355), .B1(new_n223), .B2(new_n697), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n254), .A2(new_n368), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n340), .A2(new_n214), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT96), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(G45), .B2(new_n701), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n801), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n747), .A2(new_n797), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n739), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n748), .A2(new_n798), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n743), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n627), .A2(new_n670), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n655), .A2(new_n335), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n349), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n352), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n352), .A2(new_n655), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n627), .A2(new_n670), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n729), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT100), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n818), .A2(new_n729), .A3(new_n820), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n823), .A2(new_n739), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n784), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(G159), .B1(G150), .B2(new_n765), .ZN(new_n828));
  INV_X1    g0628(.A(G143), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n829), .B2(new_n780), .C1(new_n772), .C2(new_n830), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT34), .Z(new_n832));
  NAND2_X1  g0632(.A1(new_n774), .A2(G68), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n752), .A2(G132), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n757), .A2(G58), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n340), .B1(new_n760), .B2(G50), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n752), .A2(G311), .B1(new_n827), .B2(G116), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n774), .A2(G87), .ZN(new_n839));
  INV_X1    g0639(.A(G294), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n780), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n340), .B1(new_n761), .B2(new_n338), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n759), .B(new_n842), .C1(G283), .C2(new_n765), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n790), .B2(new_n772), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n832), .A2(new_n837), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n797), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n797), .A2(new_n745), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n739), .B1(new_n261), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n745), .B2(new_n817), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n826), .A2(new_n851), .ZN(G384));
  NAND3_X1  g0652(.A1(new_n237), .A2(G77), .A3(new_n413), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(G50), .B2(new_n203), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(G1), .A3(new_n647), .ZN(new_n855));
  OAI211_X1 g0655(.A(G116), .B(new_n236), .C1(new_n473), .C2(KEYINPUT35), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(KEYINPUT35), .B2(new_n473), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(new_n857), .B2(KEYINPUT36), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(KEYINPUT36), .B2(new_n857), .ZN(new_n859));
  INV_X1    g0659(.A(new_n726), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n728), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n457), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT104), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT40), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n420), .B(new_n653), .C1(new_n444), .C2(new_n445), .ZN(new_n866));
  INV_X1    g0666(.A(new_n653), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n427), .B(new_n867), .C1(new_n350), .C2(new_n426), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n420), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n869), .A2(new_n870), .A3(new_n437), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n869), .B2(new_n437), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n203), .B1(new_n406), .B2(new_n407), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n395), .B1(new_n403), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n416), .A3(new_n257), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n419), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n653), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n444), .B2(new_n445), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n868), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n870), .B1(new_n883), .B2(new_n437), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT102), .B1(new_n871), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n426), .A2(G179), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n426), .A2(new_n350), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n888), .A2(new_n867), .B1(new_n878), .B2(new_n419), .ZN(new_n889));
  INV_X1    g0689(.A(new_n437), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT102), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n869), .A2(new_n870), .A3(new_n437), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n882), .A2(new_n885), .A3(KEYINPUT38), .A4(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT103), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n875), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n670), .A2(new_n283), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n315), .A2(new_n317), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n900), .B1(new_n901), .B2(new_n631), .ZN(new_n902));
  INV_X1    g0702(.A(new_n900), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n326), .A2(new_n318), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n817), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n862), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n865), .B1(new_n899), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n885), .A2(new_n894), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n880), .B1(new_n431), .B2(new_n441), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n895), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n907), .A2(new_n865), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n661), .B1(new_n864), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n864), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n902), .A2(new_n904), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n816), .B(KEYINPUT101), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(new_n820), .B2(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n921), .A2(new_n913), .B1(new_n444), .B2(new_n867), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n912), .B2(new_n895), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n871), .A2(new_n884), .A3(KEYINPUT102), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n927), .A2(KEYINPUT103), .A3(KEYINPUT38), .A4(new_n882), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n895), .A2(new_n896), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n874), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n924), .B1(new_n930), .B2(new_n923), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n326), .A2(new_n655), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n922), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT29), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n812), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n448), .A2(new_n936), .A3(new_n456), .A4(new_n707), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n643), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n934), .B(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n917), .A2(new_n939), .B1(new_n271), .B2(new_n648), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n940), .A2(KEYINPUT105), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n917), .A2(new_n939), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n940), .B2(KEYINPUT105), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n859), .B1(new_n941), .B2(new_n943), .ZN(G367));
  NAND2_X1  g0744(.A1(new_n655), .A2(new_n476), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n506), .A2(new_n945), .B1(new_n625), .B2(new_n655), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n677), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n679), .B1(new_n673), .B2(new_n674), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT42), .B1(new_n948), .B2(new_n946), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT42), .ZN(new_n950));
  INV_X1    g0750(.A(new_n946), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n690), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n617), .A2(new_n655), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n951), .B2(new_n691), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n949), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n655), .A2(new_n572), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n577), .B(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n960));
  INV_X1    g0760(.A(new_n957), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n949), .A2(new_n952), .A3(new_n954), .A4(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT106), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n955), .A2(new_n965), .A3(new_n958), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n947), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n960), .A2(new_n963), .A3(new_n947), .A4(new_n966), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n968), .A2(KEYINPUT107), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(KEYINPUT107), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n698), .B(KEYINPUT41), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n692), .A2(new_n974), .A3(new_n951), .ZN(new_n975));
  INV_X1    g0775(.A(new_n691), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n948), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT44), .B1(new_n977), .B2(new_n946), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT45), .B1(new_n692), .B2(new_n951), .ZN(new_n979));
  AND4_X1   g0779(.A1(KEYINPUT45), .A2(new_n948), .A3(new_n976), .A4(new_n951), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n975), .A2(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n677), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n974), .B1(new_n692), .B2(new_n951), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n977), .A2(KEYINPUT44), .A3(new_n946), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(new_n677), .C1(new_n980), .C2(new_n979), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n675), .A2(new_n680), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n988), .A2(new_n662), .A3(new_n948), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n662), .B1(new_n988), .B2(new_n948), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n731), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n983), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n973), .B1(new_n992), .B2(new_n732), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT108), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n734), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI211_X1 g0795(.A(KEYINPUT108), .B(new_n973), .C1(new_n992), .C2(new_n732), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n971), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n804), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n247), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n807), .B1(new_n214), .B2(new_n331), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n740), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n760), .A2(G116), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT46), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n340), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1002), .A2(new_n1003), .B1(new_n765), .B2(G294), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n338), .B2(new_n758), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G283), .C2(new_n827), .ZN(new_n1007));
  INV_X1    g0807(.A(G317), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n752), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1008), .A2(new_n1009), .B1(new_n775), .B2(new_n547), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G303), .B2(new_n781), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1007), .B(new_n1011), .C1(new_n788), .C2(new_n772), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n284), .B1(new_n761), .B2(new_n202), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n775), .A2(new_n261), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G159), .C2(new_n765), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n757), .A2(G68), .ZN(new_n1016));
  INV_X1    g0816(.A(G150), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n1017), .B2(new_n780), .C1(new_n772), .C2(new_n829), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT109), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n752), .A2(G137), .B1(new_n827), .B2(G50), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1015), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1012), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT47), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n797), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1001), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n747), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n961), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n997), .A2(new_n1031), .ZN(G387));
  OAI21_X1  g0832(.A(new_n804), .B1(new_n243), .B2(new_n368), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n800), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n696), .B2(new_n1034), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n328), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT50), .B1(new_n328), .B2(G50), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1036), .A2(new_n696), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1035), .A2(new_n1039), .B1(new_n338), .B2(new_n697), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n807), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n740), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n780), .A2(new_n208), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n284), .B1(new_n761), .B2(new_n261), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(new_n330), .C2(new_n757), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n784), .A2(new_n203), .B1(new_n328), .B2(new_n764), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT110), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n771), .A2(G159), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G97), .A2(new_n774), .B1(new_n752), .B2(G150), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n284), .B1(new_n752), .B2(G326), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n771), .A2(G322), .B1(G311), .B2(new_n765), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n790), .A2(new_n784), .B1(new_n780), .B2(new_n1008), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1053), .A2(KEYINPUT111), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(KEYINPUT111), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT48), .Z(new_n1057));
  OAI22_X1  g0857(.A1(new_n758), .A2(new_n787), .B1(new_n761), .B2(new_n840), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1051), .B1(new_n223), .B2(new_n775), .C1(new_n1059), .C2(KEYINPUT49), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1059), .A2(KEYINPUT49), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1050), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT112), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1027), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1042), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n676), .B2(new_n1030), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT113), .Z(new_n1068));
  NOR2_X1   g0868(.A1(new_n991), .A2(new_n699), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n989), .A2(new_n990), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n732), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n737), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1068), .A2(new_n1071), .A3(new_n1072), .ZN(G393));
  AND2_X1   g0873(.A1(new_n983), .A2(new_n987), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n946), .A2(new_n747), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n807), .B1(new_n214), .B2(new_n547), .C1(new_n998), .C2(new_n251), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n740), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n284), .B1(new_n761), .B2(new_n404), .C1(new_n758), .C2(new_n261), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n839), .B1(new_n328), .B2(new_n784), .C1(new_n1009), .C2(new_n829), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G50), .C2(new_n765), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n771), .A2(G150), .B1(new_n781), .B2(G159), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT51), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n784), .A2(new_n840), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1084), .B(new_n776), .C1(G322), .C2(new_n752), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n772), .A2(new_n1008), .B1(new_n788), .B2(new_n780), .ZN(new_n1086));
  XOR2_X1   g0886(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n340), .B1(new_n761), .B2(new_n787), .C1(new_n758), .C2(new_n223), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G303), .B2(new_n765), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1085), .A2(new_n1088), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT115), .B1(new_n1083), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n1027), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1083), .A2(KEYINPUT115), .A3(new_n1092), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1077), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1074), .A2(new_n737), .B1(new_n1075), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1074), .A2(new_n991), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n992), .A2(new_n698), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G390));
  AOI211_X1 g0900(.A(KEYINPUT39), .B(new_n874), .C1(new_n928), .C2(new_n929), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n820), .A2(new_n920), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n932), .B1(new_n1102), .B2(new_n918), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1101), .A2(new_n1103), .A3(new_n924), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n706), .A2(new_n670), .A3(new_n815), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n816), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n918), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n899), .A2(new_n933), .A3(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n905), .A2(G330), .A3(new_n862), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1104), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n729), .A2(new_n905), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n923), .B(new_n875), .C1(new_n897), .C2(new_n898), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n924), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(new_n932), .C2(new_n921), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n899), .A2(new_n933), .A3(new_n1107), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1111), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT116), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n918), .B1(new_n729), .B2(new_n819), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1102), .B1(new_n1118), .B2(new_n1109), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n862), .A2(G330), .A3(new_n819), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n919), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1121), .A2(new_n816), .A3(new_n1111), .A4(new_n1105), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n448), .A2(G330), .A3(new_n456), .A4(new_n862), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n643), .A2(new_n937), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT117), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1125), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT117), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1109), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT116), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1114), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1117), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1125), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1132), .A2(new_n1137), .A3(new_n1134), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1138), .A2(new_n698), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1110), .A2(new_n1116), .A3(new_n734), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n931), .A2(new_n745), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n340), .B1(new_n761), .B2(new_n512), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G77), .B2(new_n757), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n338), .B2(new_n764), .C1(new_n787), .C2(new_n772), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n833), .B1(new_n1009), .B2(new_n840), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n223), .A2(new_n780), .B1(new_n784), .B2(new_n547), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n781), .A2(G132), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT118), .Z(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1149), .B1(new_n1152), .B2(new_n784), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n760), .A2(G150), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT53), .Z(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n830), .B2(new_n764), .C1(new_n398), .C2(new_n758), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1153), .B(new_n1156), .C1(G128), .C2(new_n771), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n340), .B1(new_n752), .B2(G125), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n208), .B2(new_n775), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT119), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1148), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n1027), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n739), .B(new_n1163), .C1(new_n328), .C2(new_n847), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1141), .B1(new_n1142), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1140), .A2(new_n1165), .ZN(G378));
  NAND2_X1  g0966(.A1(new_n394), .A2(new_n637), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n452), .A2(new_n653), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(G330), .B1(new_n908), .B2(new_n914), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n913), .A2(new_n1102), .A3(new_n918), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n444), .A2(new_n867), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n932), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT40), .B1(new_n930), .B2(new_n906), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n907), .A2(new_n865), .A3(new_n913), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n661), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n934), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1171), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1171), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n934), .A2(new_n1181), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n847), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n740), .B1(G50), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n340), .B2(new_n367), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1009), .A2(new_n787), .B1(new_n331), .B2(new_n784), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n774), .A2(G58), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n338), .B2(new_n780), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n772), .A2(new_n223), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G41), .B(new_n284), .C1(new_n760), .C2(G77), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(new_n1016), .C1(new_n459), .C2(new_n764), .ZN(new_n1198));
  OR4_X1    g0998(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1192), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT120), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1151), .A2(new_n760), .B1(new_n781), .B2(G128), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n765), .A2(G132), .B1(new_n757), .B2(G150), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n830), .C2(new_n784), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G125), .B2(new_n771), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n774), .A2(G159), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n752), .C2(G124), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1202), .B1(new_n1200), .B2(new_n1199), .C1(new_n1208), .C2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1190), .B1(new_n1213), .B2(new_n797), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1171), .B2(new_n746), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1215), .A2(KEYINPUT121), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(KEYINPUT121), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1188), .A2(new_n737), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1138), .A2(new_n1127), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1185), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1219), .B(KEYINPUT57), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n698), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT57), .B1(new_n1188), .B2(new_n1219), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1218), .B1(new_n1223), .B2(new_n1224), .ZN(G375));
  OAI211_X1 g1025(.A(new_n1131), .B(new_n972), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G128), .A2(new_n752), .B1(new_n1151), .B2(new_n765), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n830), .B2(new_n780), .C1(new_n1017), .C2(new_n784), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n340), .B1(new_n760), .B2(G159), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1194), .B(new_n1229), .C1(new_n208), .C2(new_n758), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n771), .A2(G132), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT122), .Z(new_n1233));
  OAI22_X1  g1033(.A1(new_n1009), .A2(new_n790), .B1(new_n338), .B2(new_n784), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1014), .B(new_n1234), .C1(G283), .C2(new_n781), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n284), .B1(new_n760), .B2(G97), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n223), .B2(new_n764), .C1(new_n331), .C2(new_n758), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G294), .B2(new_n771), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1231), .A2(new_n1233), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n740), .B1(G68), .B2(new_n1189), .C1(new_n1239), .C2(new_n1027), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n919), .B2(new_n745), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1128), .B2(new_n737), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1226), .A2(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT123), .ZN(G381));
  OR4_X1    g1044(.A1(G396), .A2(G390), .A3(G393), .A4(G384), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT57), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n698), .A3(new_n1222), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1140), .A2(new_n1165), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1218), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G387), .A2(new_n1245), .A3(new_n1251), .A4(G381), .ZN(G407));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(G343), .C2(new_n1251), .ZN(G409));
  INV_X1    g1053(.A(G213), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(G343), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1137), .A2(new_n699), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1123), .A2(KEYINPUT60), .A3(new_n1125), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT60), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1260), .A2(G384), .A3(new_n1242), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G384), .B1(new_n1260), .B2(new_n1242), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G2897), .B(new_n1255), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1262), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1260), .A2(G384), .A3(new_n1242), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1255), .A2(G2897), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1250), .B1(new_n1249), .B2(new_n1218), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1219), .B(new_n972), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n737), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n1273), .A2(G378), .B1(new_n1254), .B2(G343), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1268), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT127), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(new_n1279), .A3(new_n1276), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G375), .A2(G378), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1255), .B1(new_n1282), .B2(new_n1250), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1281), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT62), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1285), .A2(KEYINPUT62), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1278), .A2(new_n1280), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(G393), .B(new_n810), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n997), .A2(new_n1031), .A3(G390), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G390), .B1(new_n997), .B2(new_n1031), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT124), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT124), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1294), .B(new_n1289), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1291), .A2(new_n1289), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n997), .A2(new_n1297), .A3(new_n1031), .A4(G390), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n997), .A2(new_n1031), .A3(G390), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT125), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1296), .A2(new_n1298), .A3(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1293), .A2(new_n1295), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1288), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1285), .A2(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1281), .A2(new_n1283), .A3(KEYINPUT63), .A4(new_n1284), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1305), .A2(new_n1276), .A3(new_n1275), .A4(new_n1306), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1302), .A2(new_n1307), .A3(KEYINPUT126), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT126), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1306), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1274), .B1(G378), .B2(G375), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT63), .B1(new_n1311), .B2(new_n1284), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1293), .A2(new_n1295), .A3(new_n1301), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1309), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1303), .B1(new_n1308), .B2(new_n1315), .ZN(G405));
  NAND2_X1  g1116(.A1(new_n1281), .A2(new_n1251), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1317), .B(new_n1284), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1318), .B(new_n1314), .ZN(G402));
endmodule


