//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1149, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G68), .B2(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT67), .B(G77), .Z(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT68), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G20), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n207), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT0), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n228), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n225), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n218), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  INV_X1    g0043(.A(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n253), .A2(new_n255), .B1(G20), .B2(new_n203), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n219), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n260), .A2(new_n262), .B1(new_n202), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n262), .ZN(new_n268));
  INV_X1    g0068(.A(G20), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(G1), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n202), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT9), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(G222), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(new_n278), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n282));
  INV_X1    g0082(.A(new_n213), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n274), .A2(new_n276), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  INV_X1    g0090(.A(new_n282), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n287), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n285), .B(new_n289), .C1(new_n290), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(G200), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n271), .A2(new_n272), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n273), .A2(new_n295), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n271), .C1(G179), .C2(new_n293), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n266), .A2(new_n253), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n270), .B2(new_n253), .ZN(new_n305));
  INV_X1    g0105(.A(G58), .ZN(new_n306));
  INV_X1    g0106(.A(G68), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n308), .A2(new_n201), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(G20), .B1(G159), .B2(new_n258), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n269), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT73), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n274), .A2(new_n276), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n274), .B2(new_n276), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n269), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT7), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(KEYINPUT16), .B(new_n310), .C1(new_n318), .C2(new_n307), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT16), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n317), .B1(new_n284), .B2(G20), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n307), .B1(new_n321), .B2(new_n311), .ZN(new_n322));
  INV_X1    g0122(.A(new_n310), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(new_n262), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT74), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n319), .A2(KEYINPUT74), .A3(new_n262), .A4(new_n324), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n305), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G232), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n289), .B1(new_n292), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT75), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n277), .B1(new_n280), .B2(new_n278), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G226), .B2(new_n278), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G87), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n291), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n294), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(new_n331), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(G200), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n329), .A2(KEYINPUT17), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT17), .B1(new_n329), .B2(new_n340), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n327), .A2(new_n328), .ZN(new_n344));
  INV_X1    g0144(.A(new_n305), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G179), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n332), .A2(new_n347), .A3(new_n337), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G169), .B2(new_n339), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(KEYINPUT18), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT76), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT76), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n346), .A2(new_n353), .A3(KEYINPUT18), .A4(new_n350), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT18), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n329), .B2(new_n349), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n303), .A2(new_n343), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n289), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT71), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n284), .A2(G226), .A3(new_n278), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n284), .A2(G232), .A3(G1698), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n365), .A2(KEYINPUT70), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(KEYINPUT70), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n363), .B(new_n364), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n359), .B1(new_n368), .B2(new_n282), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT13), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n291), .A2(G238), .A3(new_n287), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n370), .B1(new_n369), .B2(new_n371), .ZN(new_n374));
  OAI21_X1  g0174(.A(G169), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT14), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n368), .A2(new_n282), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n371), .A3(new_n289), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT13), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(G179), .A3(new_n372), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(G169), .C1(new_n373), .C2(new_n374), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n255), .A2(G77), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n202), .B2(new_n259), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n269), .A2(G68), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n262), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT11), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n387), .A2(new_n388), .B1(new_n307), .B2(new_n270), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n387), .A2(new_n388), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n264), .A2(new_n386), .ZN(new_n391));
  XOR2_X1   g0191(.A(new_n391), .B(KEYINPUT12), .Z(new_n392));
  NOR3_X1   g0192(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n383), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT72), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n379), .A2(G190), .A3(new_n372), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n393), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n379), .B2(new_n372), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n400), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n402), .A2(KEYINPUT72), .A3(new_n397), .A4(new_n393), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G238), .A2(G1698), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n284), .B(new_n406), .C1(new_n330), .C2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n282), .C1(G107), .C2(new_n284), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n408), .B(new_n289), .C1(new_n212), .C2(new_n292), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n300), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n268), .B(G77), .C1(G1), .C2(new_n269), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n213), .A2(new_n269), .B1(new_n252), .B2(new_n259), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT15), .B(G87), .Z(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n255), .B2(new_n413), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n411), .B1(new_n283), .B2(new_n265), .C1(new_n414), .C2(new_n268), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n410), .B(new_n415), .C1(G179), .C2(new_n409), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n409), .A2(G200), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n294), .B2(new_n409), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n418), .B2(new_n415), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n358), .A2(new_n405), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n266), .A2(new_n246), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n268), .B(new_n265), .C1(G1), .C2(new_n254), .ZN(new_n422));
  AOI21_X1  g0222(.A(G20), .B1(G33), .B2(G283), .ZN(new_n423));
  INV_X1    g0223(.A(G97), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(G33), .B2(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n425), .B(new_n262), .C1(new_n269), .C2(G116), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT20), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n426), .A2(new_n427), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n421), .B1(new_n246), .B2(new_n422), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n278), .A2(G257), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G264), .A2(G1698), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n284), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(new_n282), .C1(G303), .C2(new_n284), .ZN(new_n434));
  INV_X1    g0234(.A(G45), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(G1), .ZN(new_n436));
  AND2_X1   g0236(.A1(KEYINPUT5), .A2(G41), .ZN(new_n437));
  NOR2_X1   g0237(.A1(KEYINPUT5), .A2(G41), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n291), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G270), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n439), .A2(new_n288), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n434), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n430), .A2(G169), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT21), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT21), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n430), .A2(new_n446), .A3(new_n443), .A4(G169), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n430), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n449), .A2(new_n347), .A3(new_n443), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n443), .A2(G200), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n449), .B(new_n452), .C1(new_n294), .C2(new_n443), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n448), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n413), .A2(new_n265), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT19), .ZN(new_n456));
  INV_X1    g0256(.A(new_n255), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(new_n424), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n284), .A2(new_n269), .ZN(new_n459));
  AOI21_X1  g0259(.A(G20), .B1(new_n362), .B2(KEYINPUT19), .ZN(new_n460));
  NOR3_X1   g0260(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n461));
  OAI221_X1 g0261(.A(new_n458), .B1(new_n307), .B2(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n455), .B1(new_n462), .B2(new_n262), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n463), .A2(KEYINPUT77), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(KEYINPUT77), .ZN(new_n465));
  INV_X1    g0265(.A(new_n413), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n464), .A2(new_n465), .B1(new_n466), .B2(new_n422), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n212), .A2(G1698), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(G238), .B2(G1698), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n469), .A2(new_n277), .B1(new_n254), .B2(new_n246), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n470), .A2(new_n282), .B1(G274), .B2(new_n436), .ZN(new_n471));
  INV_X1    g0271(.A(new_n436), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n291), .A2(G250), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n300), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n471), .A2(new_n347), .A3(new_n473), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n467), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G87), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n422), .A2(new_n478), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n463), .A2(KEYINPUT77), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n463), .A2(KEYINPUT77), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n474), .A2(new_n294), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(G200), .B2(new_n474), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n454), .A2(new_n477), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n284), .A2(G244), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT4), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n487), .A2(new_n488), .B1(G33), .B2(G283), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n278), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n284), .B2(G250), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n278), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n282), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n440), .A2(G257), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(G190), .A3(new_n495), .A4(new_n442), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n258), .A2(G77), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n424), .A2(new_n244), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n244), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n321), .A2(new_n311), .ZN(new_n504));
  OAI221_X1 g0304(.A(new_n497), .B1(new_n269), .B2(new_n503), .C1(new_n504), .C2(new_n244), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n262), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n266), .A2(new_n424), .ZN(new_n507));
  INV_X1    g0307(.A(new_n422), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G97), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n496), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n489), .B(new_n490), .C1(new_n278), .C2(new_n492), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(new_n282), .B1(G257), .B2(new_n440), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n399), .B1(new_n512), .B2(new_n442), .ZN(new_n513));
  OR2_X1    g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n244), .A2(G20), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n515), .B(KEYINPUT23), .ZN(new_n516));
  NAND2_X1  g0316(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n459), .B2(new_n478), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n284), .A2(new_n269), .A3(G87), .A4(new_n517), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT24), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n255), .A2(G116), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n262), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n515), .A2(G1), .A3(new_n263), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT25), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n508), .A2(G107), .B1(new_n528), .B2(new_n527), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n442), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n284), .B1(G250), .B2(G1698), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n278), .A2(G257), .ZN(new_n534));
  INV_X1    g0334(.A(G294), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n533), .A2(new_n534), .B1(new_n254), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n536), .B2(new_n282), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n440), .A2(G264), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT79), .B1(new_n440), .B2(G264), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n440), .A2(KEYINPUT79), .A3(G264), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n539), .A2(new_n300), .B1(new_n542), .B2(new_n347), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n531), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n294), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n399), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n547), .A2(new_n529), .A3(new_n526), .A4(new_n530), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n494), .A2(new_n495), .A3(new_n442), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n347), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n512), .A2(new_n442), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n300), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n514), .A2(new_n544), .A3(new_n548), .A4(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n486), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n420), .A2(new_n556), .ZN(G372));
  INV_X1    g0357(.A(new_n302), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n351), .A2(new_n356), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n416), .B(KEYINPUT82), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n404), .A2(new_n560), .B1(new_n394), .B2(new_n383), .ZN(new_n561));
  INV_X1    g0361(.A(new_n343), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n558), .B1(new_n563), .B2(new_n299), .ZN(new_n564));
  INV_X1    g0364(.A(new_n420), .ZN(new_n565));
  XOR2_X1   g0365(.A(new_n475), .B(KEYINPUT80), .Z(new_n566));
  NAND3_X1  g0366(.A1(new_n467), .A2(new_n476), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n477), .A2(new_n569), .A3(new_n485), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n568), .B1(new_n570), .B2(KEYINPUT26), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n510), .A2(new_n513), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n450), .B1(new_n445), .B2(new_n447), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n544), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n569), .B1(new_n574), .B2(new_n548), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT81), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n480), .A2(new_n481), .ZN(new_n577));
  INV_X1    g0377(.A(new_n479), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI211_X1 g0379(.A(KEYINPUT81), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n484), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT26), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n571), .B1(new_n575), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n564), .B1(new_n565), .B2(new_n585), .ZN(G369));
  NOR2_X1   g0386(.A1(new_n263), .A2(G20), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n286), .ZN(new_n588));
  XOR2_X1   g0388(.A(new_n588), .B(KEYINPUT83), .Z(new_n589));
  OR2_X1    g0389(.A1(new_n589), .A2(KEYINPUT27), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(KEYINPUT27), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n591), .A3(G213), .ZN(new_n592));
  INV_X1    g0392(.A(G343), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n454), .B1(new_n449), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n573), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n430), .A3(new_n594), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g0400(.A(KEYINPUT84), .B(G330), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n531), .A2(new_n594), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT85), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT85), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n531), .A2(new_n607), .A3(new_n594), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n606), .A2(new_n544), .A3(new_n548), .A4(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n531), .A2(new_n543), .A3(new_n594), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n597), .A2(new_n595), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n544), .A2(new_n594), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(G399));
  INV_X1    g0418(.A(G41), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n226), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n461), .A2(new_n246), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n621), .A2(new_n622), .A3(new_n286), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n224), .B2(new_n621), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT86), .ZN(new_n625));
  XOR2_X1   g0425(.A(new_n625), .B(KEYINPUT28), .Z(new_n626));
  NOR3_X1   g0426(.A1(new_n585), .A2(KEYINPUT29), .A3(new_n594), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT29), .ZN(new_n628));
  INV_X1    g0428(.A(new_n484), .ZN(new_n629));
  INV_X1    g0429(.A(new_n579), .ZN(new_n630));
  INV_X1    g0430(.A(new_n580), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT26), .B1(new_n632), .B2(new_n554), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n477), .A2(new_n485), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n582), .A3(new_n569), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n581), .A2(new_n574), .A3(new_n554), .A4(new_n548), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n633), .A2(new_n635), .A3(new_n567), .A4(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n628), .B1(new_n637), .B2(new_n595), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n627), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n542), .A2(new_n347), .A3(new_n474), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n434), .A2(new_n441), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n549), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT30), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n443), .A2(new_n347), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n551), .A2(new_n542), .A3(new_n474), .A4(new_n645), .ZN(new_n646));
  AOI211_X1 g0446(.A(KEYINPUT31), .B(new_n595), .C1(new_n644), .C2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT31), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n556), .B2(new_n595), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n644), .A2(new_n646), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n594), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n647), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n601), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n639), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n626), .B1(new_n655), .B2(G1), .ZN(G364));
  NAND2_X1  g0456(.A1(new_n587), .A2(G45), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n620), .A2(G1), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n600), .A2(new_n602), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n604), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n314), .A2(new_n315), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n226), .ZN(new_n663));
  XOR2_X1   g0463(.A(new_n663), .B(KEYINPUT88), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n250), .A2(G45), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n664), .B(new_n665), .C1(G45), .C2(new_n223), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n284), .A2(G355), .A3(new_n226), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n666), .B(new_n667), .C1(G116), .C2(new_n226), .ZN(new_n668));
  NOR2_X1   g0468(.A1(G13), .A2(G33), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G20), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n219), .B1(G20), .B2(new_n300), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n658), .B(KEYINPUT87), .Z(new_n675));
  NOR2_X1   g0475(.A1(new_n269), .A2(new_n294), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n347), .A2(new_n399), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(KEYINPUT91), .B(G326), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n347), .A2(G200), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n269), .A2(G190), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G311), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n682), .ZN(new_n685));
  XOR2_X1   g0485(.A(KEYINPUT33), .B(G317), .Z(new_n686));
  OAI221_X1 g0486(.A(new_n277), .B1(new_n683), .B2(new_n684), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(G179), .A2(G200), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n269), .B1(new_n688), .B2(G190), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI211_X1 g0490(.A(new_n680), .B(new_n687), .C1(G294), .C2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n676), .A2(new_n347), .A3(G200), .ZN(new_n692));
  INV_X1    g0492(.A(G303), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n682), .A2(new_n688), .ZN(new_n694));
  INV_X1    g0494(.A(G329), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n692), .A2(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR4_X1   g0496(.A1(new_n269), .A2(new_n399), .A3(G179), .A4(G190), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT90), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT90), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n696), .B1(new_n701), .B2(G283), .ZN(new_n702));
  INV_X1    g0502(.A(G322), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n676), .A2(new_n681), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n691), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n689), .A2(new_n424), .ZN(new_n706));
  OAI221_X1 g0506(.A(new_n284), .B1(new_n685), .B2(new_n307), .C1(new_n478), .C2(new_n692), .ZN(new_n707));
  INV_X1    g0507(.A(new_n678), .ZN(new_n708));
  AOI211_X1 g0508(.A(new_n706), .B(new_n707), .C1(G50), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n701), .A2(G107), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n213), .A2(new_n683), .B1(new_n704), .B2(new_n306), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT89), .Z(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n694), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G159), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT32), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n705), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n675), .B1(new_n717), .B2(new_n672), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n671), .B(KEYINPUT92), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n674), .B(new_n718), .C1(new_n599), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n660), .A2(new_n721), .ZN(G396));
  NAND2_X1  g0522(.A1(new_n594), .A2(new_n415), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n560), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n419), .A2(new_n723), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n584), .A2(new_n595), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n585), .A2(new_n594), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n726), .B(KEYINPUT94), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(new_n653), .Z(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n658), .ZN(new_n733));
  INV_X1    g0533(.A(new_n704), .ZN(new_n734));
  INV_X1    g0534(.A(new_n685), .ZN(new_n735));
  AOI22_X1  g0535(.A1(G143), .A2(new_n734), .B1(new_n735), .B2(G150), .ZN(new_n736));
  INV_X1    g0536(.A(G137), .ZN(new_n737));
  INV_X1    g0537(.A(G159), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n736), .B1(new_n737), .B2(new_n678), .C1(new_n738), .C2(new_n683), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT34), .ZN(new_n740));
  INV_X1    g0540(.A(G132), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n661), .B1(new_n306), .B2(new_n689), .C1(new_n741), .C2(new_n694), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n701), .B2(G68), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n740), .B(new_n743), .C1(new_n202), .C2(new_n692), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n277), .B1(new_n683), .B2(new_n246), .C1(new_n693), .C2(new_n678), .ZN(new_n745));
  INV_X1    g0545(.A(new_n692), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n706), .B(new_n745), .C1(G107), .C2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT93), .B(G283), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n685), .A2(new_n748), .B1(new_n694), .B2(new_n684), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n701), .B2(G87), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n747), .B(new_n750), .C1(new_n535), .C2(new_n704), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n744), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n675), .B1(new_n752), .B2(new_n672), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n672), .A2(new_n669), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n753), .B1(G77), .B2(new_n755), .C1(new_n727), .C2(new_n670), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n733), .A2(new_n756), .ZN(G384));
  INV_X1    g0557(.A(new_n503), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n246), .B1(new_n758), .B2(KEYINPUT35), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n759), .B(new_n222), .C1(KEYINPUT35), .C2(new_n758), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT36), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n213), .A2(new_n308), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n762), .A2(new_n223), .B1(G50), .B2(new_n307), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G1), .A3(new_n263), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT95), .Z(new_n766));
  INV_X1    g0566(.A(KEYINPUT98), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT38), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n344), .A2(new_n340), .A3(new_n345), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n329), .B2(new_n592), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n329), .A2(new_n349), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n770), .A2(KEYINPUT37), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n277), .A2(KEYINPUT73), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n274), .A2(new_n276), .A3(new_n313), .ZN(new_n774));
  AOI21_X1  g0574(.A(G20), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n311), .B1(new_n775), .B2(KEYINPUT7), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n323), .B1(new_n776), .B2(G68), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n262), .B1(new_n777), .B2(KEYINPUT16), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT96), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n310), .B1(new_n318), .B2(new_n307), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n268), .B1(new_n780), .B2(new_n320), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT96), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n779), .A2(new_n783), .A3(new_n319), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n349), .B1(new_n784), .B2(new_n345), .ZN(new_n785));
  AND3_X1   g0585(.A1(new_n344), .A2(new_n340), .A3(new_n345), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT97), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT97), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n781), .A2(new_n782), .B1(KEYINPUT16), .B2(new_n777), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n305), .B1(new_n789), .B2(new_n779), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n769), .B(new_n788), .C1(new_n790), .C2(new_n349), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n592), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n787), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n772), .B1(new_n794), .B2(KEYINPUT37), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n793), .B1(new_n357), .B2(new_n343), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n768), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n354), .A2(new_n356), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n353), .B1(new_n771), .B2(KEYINPUT18), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n343), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n792), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT37), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n769), .B1(new_n790), .B2(new_n349), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n792), .B1(new_n803), .B2(KEYINPUT97), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n802), .B1(new_n804), .B2(new_n791), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n801), .B(KEYINPUT38), .C1(new_n772), .C2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n767), .B1(new_n797), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n797), .A2(new_n806), .A3(new_n767), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n595), .A2(new_n393), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n405), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n395), .B(new_n404), .C1(new_n393), .C2(new_n595), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n555), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n815), .A2(new_n634), .A3(new_n454), .A4(new_n595), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n816), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n817));
  INV_X1    g0617(.A(new_n647), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n817), .A2(new_n818), .A3(new_n727), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n808), .A2(new_n809), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT40), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT100), .ZN(new_n824));
  INV_X1    g0624(.A(new_n592), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n346), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT17), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n769), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n329), .A2(KEYINPUT17), .A3(new_n340), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT18), .B1(new_n346), .B2(new_n350), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n329), .A2(new_n355), .A3(new_n349), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT37), .B1(new_n770), .B2(new_n771), .ZN(new_n834));
  INV_X1    g0634(.A(new_n771), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n835), .A2(new_n826), .A3(new_n802), .A4(new_n769), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n827), .A2(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n824), .B1(new_n837), .B2(KEYINPUT38), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n834), .A2(new_n836), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n826), .B1(new_n343), .B2(new_n559), .ZN(new_n840));
  OAI211_X1 g0640(.A(KEYINPUT100), .B(new_n768), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n838), .A2(new_n806), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT101), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n814), .A2(new_n819), .A3(new_n822), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n838), .A2(new_n806), .A3(KEYINPUT101), .A4(new_n841), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n823), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n420), .A2(new_n652), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n601), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n797), .A2(new_n806), .A3(new_n767), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n416), .A2(new_n594), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n728), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n813), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n852), .A2(new_n807), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n559), .A2(new_n825), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT99), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT39), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n842), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n797), .A2(new_n806), .A3(KEYINPUT39), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n395), .A2(new_n594), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n856), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n808), .A2(new_n866), .A3(new_n809), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT99), .ZN(new_n868));
  INV_X1    g0668(.A(new_n858), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n859), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n420), .B1(new_n627), .B2(new_n638), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n564), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n871), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n851), .B(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n587), .A2(new_n286), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n766), .B1(new_n875), .B2(new_n876), .ZN(G367));
  NAND3_X1  g0677(.A1(new_n630), .A2(new_n631), .A3(new_n594), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n632), .B2(new_n568), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n568), .B2(new_n878), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT102), .Z(new_n881));
  INV_X1    g0681(.A(KEYINPUT43), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n615), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n553), .A2(new_n594), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n514), .A2(new_n554), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n886), .B1(new_n554), .B2(new_n595), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT103), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n554), .B1(new_n890), .B2(new_n544), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n595), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n883), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT104), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n881), .A2(new_n882), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n883), .A2(new_n893), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n896), .A2(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT105), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n613), .A2(new_n890), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n901), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n620), .B(KEYINPUT41), .Z(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT106), .B1(new_n611), .B2(new_n614), .ZN(new_n909));
  MUX2_X1   g0709(.A(KEYINPUT106), .B(new_n909), .S(new_n884), .Z(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(new_n603), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n654), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n617), .A2(new_n889), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT45), .Z(new_n915));
  NOR2_X1   g0715(.A1(new_n617), .A2(new_n889), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT44), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(new_n613), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n913), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n908), .B1(new_n921), .B2(new_n655), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n657), .A2(G1), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n905), .B(new_n906), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n881), .A2(new_n719), .ZN(new_n925));
  INV_X1    g0725(.A(new_n664), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n673), .B1(new_n226), .B2(new_n466), .C1(new_n926), .C2(new_n240), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n661), .B1(G311), .B2(new_n708), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n928), .B1(new_n244), .B2(new_n689), .C1(new_n535), .C2(new_n685), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT108), .B1(new_n692), .B2(new_n246), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT46), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n701), .A2(G97), .ZN(new_n932));
  INV_X1    g0732(.A(G317), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n683), .A2(new_n748), .B1(new_n694), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n929), .B(new_n936), .C1(G303), .C2(new_n734), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n689), .A2(new_n307), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n284), .B1(new_n694), .B2(new_n737), .C1(new_n692), .C2(new_n306), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n938), .B(new_n939), .C1(G150), .C2(new_n734), .ZN(new_n940));
  INV_X1    g0740(.A(new_n683), .ZN(new_n941));
  AOI22_X1  g0741(.A1(G159), .A2(new_n735), .B1(new_n941), .B2(G50), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n940), .B(new_n942), .C1(new_n213), .C2(new_n700), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G143), .B2(new_n708), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT109), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT47), .Z(new_n947));
  AOI21_X1  g0747(.A(new_n675), .B1(new_n947), .B2(new_n672), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n925), .A2(new_n927), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n924), .A2(new_n949), .ZN(G387));
  INV_X1    g0750(.A(new_n911), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n923), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT110), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n951), .A2(new_n655), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n954), .A2(new_n620), .A3(new_n912), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n746), .A2(new_n283), .ZN(new_n956));
  XNOR2_X1  g0756(.A(KEYINPUT112), .B(G150), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n956), .B1(new_n694), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT113), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n941), .A2(G68), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G159), .A2(new_n708), .B1(new_n735), .B2(new_n253), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n202), .B2(new_n704), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n466), .A2(new_n689), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n963), .A2(new_n662), .A3(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n960), .A2(new_n932), .A3(new_n961), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G311), .A2(new_n735), .B1(new_n734), .B2(G317), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n693), .B2(new_n683), .C1(new_n703), .C2(new_n678), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT48), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n535), .B2(new_n692), .C1(new_n689), .C2(new_n748), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT49), .Z(new_n971));
  OAI221_X1 g0771(.A(new_n662), .B1(new_n679), .B2(new_n694), .C1(new_n700), .C2(new_n246), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT114), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n966), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n675), .B1(new_n974), .B2(new_n672), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n253), .A2(new_n202), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n622), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n978));
  NAND2_X1  g0778(.A1(G68), .A2(G77), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n977), .A2(new_n978), .A3(new_n435), .A4(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n664), .B(new_n980), .C1(new_n435), .C2(new_n237), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n284), .A2(new_n622), .A3(new_n226), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(G107), .B2(new_n226), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT111), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n673), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n611), .A2(new_n719), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n975), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n953), .A2(new_n955), .A3(new_n988), .ZN(G393));
  OAI211_X1 g0789(.A(new_n921), .B(new_n621), .C1(new_n919), .C2(new_n912), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n890), .A2(new_n671), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n673), .B1(new_n424), .B2(new_n226), .C1(new_n926), .C2(new_n247), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n678), .A2(new_n933), .B1(new_n704), .B2(new_n684), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT52), .Z(new_n994));
  OAI22_X1  g0794(.A1(new_n685), .A2(new_n693), .B1(new_n689), .B2(new_n246), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n284), .B1(new_n714), .B2(G322), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n710), .B(new_n996), .C1(new_n692), .C2(new_n748), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n994), .B(new_n995), .C1(new_n997), .C2(KEYINPUT116), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(KEYINPUT116), .B2(new_n997), .C1(new_n535), .C2(new_n683), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n701), .A2(G87), .B1(G143), .B2(new_n714), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n678), .A2(new_n257), .B1(new_n704), .B2(new_n738), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT51), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n662), .B1(G68), .B2(new_n746), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n690), .A2(G77), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n202), .B2(new_n685), .C1(new_n252), .C2(new_n683), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT115), .Z(new_n1007));
  OAI21_X1  g0807(.A(new_n999), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n675), .B1(new_n1008), .B2(new_n672), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n991), .A2(new_n992), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n919), .B2(new_n923), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n990), .A2(new_n1011), .ZN(G390));
  NAND2_X1  g0812(.A1(new_n861), .A2(new_n862), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n864), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n856), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n652), .A2(new_n601), .A3(new_n727), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(new_n814), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n637), .A2(new_n595), .A3(new_n727), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n854), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n813), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1022), .A2(new_n844), .A3(new_n1014), .A4(new_n846), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(KEYINPUT117), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(KEYINPUT117), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1016), .B(new_n1019), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1023), .A2(KEYINPUT117), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1023), .A2(KEYINPUT117), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1027), .A2(new_n1028), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n820), .A2(G330), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1026), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n849), .A2(G330), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n564), .A3(new_n872), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1017), .A2(new_n814), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n855), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n652), .A2(new_n730), .A3(G330), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n814), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1018), .A2(new_n854), .A3(new_n1020), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1034), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1032), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1016), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n1030), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1040), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n1026), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1041), .A2(new_n621), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(G283), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n678), .A2(new_n1047), .B1(new_n683), .B2(new_n424), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G107), .B2(new_n735), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT118), .Z(new_n1050));
  NAND2_X1  g0850(.A1(new_n701), .A2(G68), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n277), .B1(new_n694), .B2(new_n535), .C1(new_n692), .C2(new_n478), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G116), .B2(new_n734), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1005), .A4(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(KEYINPUT54), .B(G143), .Z(new_n1055));
  AOI22_X1  g0855(.A1(new_n735), .A2(G137), .B1(new_n941), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n714), .A2(G125), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n741), .C2(new_n704), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n277), .B(new_n1058), .C1(G159), .C2(new_n690), .ZN(new_n1059));
  INV_X1    g0859(.A(G128), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1059), .B1(new_n202), .B2(new_n700), .C1(new_n1060), .C2(new_n678), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n746), .A2(new_n957), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT53), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1054), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n675), .B1(new_n1064), .B2(new_n672), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n863), .B2(new_n670), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n252), .B2(new_n754), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n1032), .B2(new_n923), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1046), .A2(new_n1068), .ZN(G378));
  NAND3_X1  g0869(.A1(new_n652), .A2(new_n813), .A3(new_n727), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n852), .A2(new_n807), .A3(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n847), .B(G330), .C1(new_n1071), .C2(KEYINPUT40), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n303), .B(KEYINPUT55), .Z(new_n1073));
  NAND2_X1  g0873(.A1(new_n825), .A2(new_n271), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT56), .Z(new_n1075));
  XNOR2_X1  g0875(.A(new_n1073), .B(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1072), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n823), .A2(G330), .A3(new_n847), .A4(new_n1076), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n871), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n871), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(KEYINPUT119), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n871), .B1(new_n1079), .B2(new_n1078), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT119), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1034), .B(KEYINPUT120), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1041), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT57), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1044), .B1(new_n1043), .B2(new_n1026), .ZN(new_n1094));
  OAI211_X1 g0894(.A(KEYINPUT57), .B(new_n1093), .C1(new_n1094), .C2(new_n1089), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n621), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1076), .A2(new_n669), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n754), .A2(new_n202), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n704), .A2(new_n1060), .B1(new_n689), .B2(new_n257), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n746), .A2(new_n1055), .B1(new_n941), .B2(G137), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n741), .B2(new_n685), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G125), .C2(new_n708), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT59), .ZN(new_n1104));
  AOI21_X1  g0904(.A(G41), .B1(new_n701), .B2(G159), .ZN(new_n1105));
  AOI21_X1  g0905(.A(G33), .B1(new_n714), .B2(G124), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n956), .B(new_n619), .C1(new_n466), .C2(new_n683), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n685), .A2(new_n424), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1108), .A2(new_n661), .A3(new_n938), .A4(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n704), .A2(new_n244), .B1(new_n694), .B2(new_n1047), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n701), .B2(G58), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(new_n246), .C2(new_n678), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT58), .ZN(new_n1114));
  AOI21_X1  g0914(.A(G41), .B1(new_n661), .B2(G33), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1107), .B(new_n1114), .C1(G50), .C2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n658), .B1(new_n1116), .B2(new_n672), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1098), .A2(new_n1099), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1088), .B2(new_n923), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1097), .A2(new_n1120), .ZN(G375));
  OAI221_X1 g0921(.A(new_n277), .B1(new_n685), .B2(new_n246), .C1(new_n424), .C2(new_n692), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n964), .B(new_n1122), .C1(G303), .C2(new_n714), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n704), .A2(new_n1047), .B1(new_n683), .B2(new_n244), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n701), .B2(G77), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(new_n535), .C2(new_n678), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT121), .Z(new_n1127));
  OAI221_X1 g0927(.A(new_n661), .B1(new_n202), .B2(new_n689), .C1(new_n257), .C2(new_n683), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G132), .B2(new_n708), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n692), .A2(new_n738), .B1(new_n694), .B2(new_n1060), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n735), .B2(new_n1055), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1129), .B(new_n1131), .C1(new_n306), .C2(new_n700), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G137), .B2(new_n734), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n672), .B1(new_n1127), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n675), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(G68), .C2(new_n755), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT122), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n814), .B2(new_n669), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n923), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1036), .A2(new_n1034), .A3(new_n1039), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n907), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1142), .B2(new_n1040), .ZN(G381));
  NOR2_X1   g0943(.A1(G375), .A2(G378), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n924), .A2(new_n949), .A3(new_n1011), .A4(new_n990), .ZN(new_n1145));
  OR2_X1    g0945(.A1(G393), .A2(G396), .ZN(new_n1146));
  NOR4_X1   g0946(.A1(new_n1145), .A2(G384), .A3(G381), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(G407));
  OAI21_X1  g0948(.A(new_n1144), .B1(new_n593), .B2(new_n1147), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(G213), .ZN(G409));
  NAND2_X1  g0950(.A1(new_n593), .A2(G213), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT125), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1141), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n620), .B1(new_n1153), .B2(KEYINPUT60), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT60), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1141), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1044), .A3(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1157), .A2(G384), .A3(new_n1140), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G384), .B1(new_n1157), .B2(new_n1140), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(G378), .B(new_n1120), .C1(new_n1092), .C2(new_n1096), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n923), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1163), .A2(KEYINPUT123), .A3(new_n1119), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT123), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n871), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n923), .B1(new_n1166), .B2(new_n1085), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n1167), .B2(new_n1118), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1088), .A2(new_n907), .A3(new_n1091), .ZN(new_n1170));
  AOI21_X1  g0970(.A(G378), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1161), .B1(new_n1171), .B2(KEYINPUT124), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT123), .B1(new_n1163), .B2(new_n1119), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1167), .A2(new_n1165), .A3(new_n1118), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1084), .B(new_n1087), .C1(new_n1094), .C2(new_n1089), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1174), .C1(new_n1175), .C2(new_n908), .ZN(new_n1176));
  INV_X1    g0976(.A(G378), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(new_n1177), .A3(KEYINPUT124), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1151), .B(new_n1160), .C1(new_n1172), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT62), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT124), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1184), .A2(new_n1178), .A3(new_n1161), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1151), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n593), .A2(G213), .A3(G2897), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n1160), .B2(KEYINPUT126), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT126), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1158), .A2(new_n1159), .A3(new_n1190), .A4(new_n1187), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1189), .A2(new_n1191), .B1(KEYINPUT126), .B2(new_n1160), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1186), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT61), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT62), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1185), .A2(new_n1196), .A3(new_n1151), .A4(new_n1160), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1181), .A2(new_n1194), .A3(new_n1195), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(G387), .A2(G390), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1145), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(G393), .B(G396), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1145), .A3(new_n1201), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1198), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1192), .B1(new_n1185), .B2(new_n1151), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT63), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1180), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1185), .A2(KEYINPUT63), .A3(new_n1151), .A4(new_n1160), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1205), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1209), .A2(new_n1212), .A3(new_n1195), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1206), .A2(new_n1213), .ZN(G405));
  NAND2_X1  g1014(.A1(G375), .A2(new_n1177), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(new_n1161), .A3(new_n1160), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G378), .B1(new_n1097), .B2(new_n1120), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1161), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1217), .A2(new_n1218), .B1(new_n1159), .B2(new_n1158), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT127), .B1(new_n1220), .B2(new_n1205), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1205), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT127), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1211), .A2(new_n1216), .A3(new_n1219), .A4(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .ZN(G402));
endmodule


