//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n207), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n213), .B(new_n224), .C1(new_n226), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND2_X1  g0045(.A1(new_n203), .A2(G20), .ZN(new_n246));
  INV_X1    g0046(.A(G150), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n207), .A2(G33), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n246), .B1(new_n247), .B2(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n225), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n252), .A2(new_n254), .B1(new_n202), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT66), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(new_n207), .B2(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n206), .A2(KEYINPUT66), .A3(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT67), .B1(new_n262), .B2(new_n202), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n256), .A2(new_n254), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT67), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n261), .A2(new_n265), .A3(G50), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n257), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n257), .A2(KEYINPUT9), .A3(new_n267), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(KEYINPUT65), .A2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT65), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  AND2_X1   g0077(.A1(G1), .A2(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n276), .A2(new_n280), .A3(new_n206), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(G226), .B2(new_n285), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G222), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(G223), .A3(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n289), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n286), .A2(new_n296), .A3(G190), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n286), .A2(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G200), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT68), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n300), .A2(KEYINPUT68), .A3(G200), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n272), .A2(new_n299), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n270), .A2(new_n301), .A3(new_n297), .A4(new_n271), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n286), .A2(new_n296), .A3(new_n311), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n310), .A2(new_n268), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n253), .A2(new_n225), .ZN(new_n317));
  INV_X1    g0117(.A(G58), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT8), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT8), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G58), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n261), .A2(new_n317), .A3(new_n255), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n251), .A2(new_n256), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(KEYINPUT72), .A3(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT16), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n287), .A2(new_n207), .A3(new_n288), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n288), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n215), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(G58), .A2(G68), .ZN(new_n336));
  OAI21_X1  g0136(.A(G20), .B1(new_n336), .B2(new_n201), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n248), .A2(KEYINPUT71), .A3(G159), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT71), .B1(new_n248), .B2(G159), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n330), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT7), .B1(new_n344), .B2(new_n207), .ZN(new_n345));
  NOR4_X1   g0145(.A1(new_n342), .A2(new_n343), .A3(new_n332), .A4(G20), .ZN(new_n346));
  OAI21_X1  g0146(.A(G68), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(KEYINPUT16), .B(new_n337), .C1(new_n338), .C2(new_n339), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n317), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n329), .B1(new_n341), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n283), .A2(G232), .A3(new_n284), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n281), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G223), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n290), .ZN(new_n356));
  INV_X1    g0156(.A(G226), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G1698), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n356), .B(new_n358), .C1(new_n342), .C2(new_n343), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G87), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n283), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n352), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n360), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n295), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n281), .A4(new_n353), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n316), .B1(new_n351), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n350), .A2(new_n341), .ZN(new_n369));
  INV_X1    g0169(.A(new_n328), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT72), .B1(new_n323), .B2(new_n324), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n369), .A2(new_n367), .A3(new_n316), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT17), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  INV_X1    g0176(.A(new_n340), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT16), .B1(new_n347), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n254), .B1(new_n335), .B2(new_n348), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n376), .B1(new_n380), .B2(new_n329), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n369), .A2(new_n372), .A3(KEYINPUT73), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n364), .A2(new_n281), .A3(new_n353), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G169), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n383), .B2(new_n311), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT18), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n369), .A2(new_n372), .A3(new_n367), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT17), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n381), .A2(new_n391), .A3(new_n382), .A4(new_n385), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n375), .A2(new_n387), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n264), .A2(G77), .A3(new_n261), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(G77), .B2(new_n255), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n322), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT15), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G87), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(new_n207), .A3(G33), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n317), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n285), .A2(G244), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n281), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n289), .A2(G232), .A3(new_n290), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n289), .A2(G238), .A3(G1698), .ZN(new_n407));
  INV_X1    g0207(.A(G107), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n406), .B(new_n407), .C1(new_n408), .C2(new_n289), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n405), .B1(new_n409), .B2(new_n295), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n403), .B1(new_n411), .B2(new_n309), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n311), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(G190), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(new_n403), .C1(new_n352), .C2(new_n410), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n315), .A2(new_n393), .A3(new_n417), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n249), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n250), .A2(new_n293), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n254), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT11), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT70), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT11), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n421), .B(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT70), .ZN(new_n427));
  INV_X1    g0227(.A(new_n264), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n428), .A2(new_n262), .A3(new_n215), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT12), .B1(new_n255), .B2(G68), .ZN(new_n430));
  OR3_X1    g0230(.A1(new_n255), .A2(KEYINPUT12), .A3(G68), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n424), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n289), .A2(G232), .A3(G1698), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT69), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n289), .A2(KEYINPUT69), .A3(G232), .A4(G1698), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G97), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n289), .A2(G226), .A3(new_n290), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n437), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n295), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n282), .B1(G238), .B2(new_n285), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT13), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n444), .B1(new_n442), .B2(new_n443), .ZN(new_n446));
  OAI21_X1  g0246(.A(G200), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(new_n443), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT13), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(G190), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n434), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(G169), .B1(new_n445), .B2(new_n446), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT14), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n449), .A2(G179), .A3(new_n450), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT14), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(G169), .C1(new_n445), .C2(new_n446), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n452), .B1(new_n458), .B2(new_n433), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n418), .A2(KEYINPUT75), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT75), .B1(new_n418), .B2(new_n459), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(G244), .B(new_n290), .C1(new_n342), .C2(new_n343), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT4), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n289), .A2(KEYINPUT4), .A3(G244), .A4(new_n290), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n289), .A2(G250), .A3(G1698), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n465), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n295), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT5), .B1(new_n273), .B2(new_n275), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n206), .B(G45), .C1(new_n472), .C2(G41), .ZN(new_n473));
  OAI211_X1 g0273(.A(G257), .B(new_n283), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n473), .ZN(new_n475));
  AND2_X1   g0275(.A1(KEYINPUT65), .A2(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT65), .A2(G41), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n478), .A3(new_n280), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n470), .A2(new_n481), .A3(new_n311), .ZN(new_n482));
  AOI21_X1  g0282(.A(G169), .B1(new_n470), .B2(new_n481), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n256), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n206), .A2(G33), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n264), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n487), .B2(new_n484), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT6), .ZN(new_n489));
  AND2_X1   g0289(.A1(G97), .A2(G107), .ZN(new_n490));
  NOR2_X1   g0290(.A1(G97), .A2(G107), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT76), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT6), .A2(G97), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(G107), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n408), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(G97), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G20), .B1(G77), .B2(new_n248), .ZN(new_n498));
  OAI21_X1  g0298(.A(G107), .B1(new_n345), .B2(new_n346), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n488), .B1(new_n500), .B2(new_n254), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n482), .A2(new_n483), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT77), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n470), .A2(new_n481), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(G200), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n470), .A2(new_n481), .A3(G190), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n504), .A2(new_n503), .A3(G200), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT19), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n207), .B1(new_n439), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n491), .A2(new_n217), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n207), .B(G68), .C1(new_n342), .C2(new_n343), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n511), .B1(new_n250), .B2(new_n484), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n254), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n264), .A2(G87), .A3(new_n486), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT15), .B(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n256), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n216), .A2(new_n290), .ZN(new_n523));
  INV_X1    g0323(.A(G244), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G1698), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n525), .C1(new_n342), .C2(new_n343), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n295), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n218), .B1(new_n274), .B2(G1), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n206), .A2(new_n277), .A3(G45), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n283), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n352), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT79), .B1(new_n522), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n283), .B1(new_n526), .B2(new_n527), .ZN(new_n536));
  OAI21_X1  g0336(.A(G200), .B1(new_n536), .B2(new_n532), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n517), .A2(new_n254), .B1(new_n256), .B2(new_n520), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT79), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n519), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n529), .A2(G190), .A3(new_n533), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n535), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT78), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n400), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n520), .A2(KEYINPUT78), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n264), .A2(new_n544), .A3(new_n545), .A4(new_n486), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n518), .A2(new_n521), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n532), .B1(new_n528), .B2(new_n295), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n311), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n309), .B1(new_n536), .B2(new_n532), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n542), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G264), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n553));
  OAI211_X1 g0353(.A(G257), .B(new_n290), .C1(new_n342), .C2(new_n343), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n287), .A2(G303), .A3(new_n288), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n295), .ZN(new_n557));
  OAI211_X1 g0357(.A(G270), .B(new_n283), .C1(new_n471), .C2(new_n473), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n479), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n264), .A2(G116), .A3(new_n486), .ZN(new_n560));
  INV_X1    g0360(.A(G116), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n256), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n253), .A2(new_n225), .B1(G20), .B2(new_n561), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n467), .B(new_n207), .C1(G33), .C2(new_n484), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n563), .A2(KEYINPUT20), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT20), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n560), .B(new_n562), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n559), .A2(new_n567), .A3(G169), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n556), .A2(new_n295), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n558), .A2(new_n479), .ZN(new_n572));
  OAI21_X1  g0372(.A(G200), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n295), .B1(new_n475), .B2(new_n478), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n273), .A2(new_n275), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n473), .B1(new_n575), .B2(new_n472), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n574), .A2(G270), .B1(new_n576), .B2(new_n280), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(G190), .A3(new_n557), .ZN(new_n578));
  INV_X1    g0378(.A(new_n567), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n567), .A2(new_n577), .A3(G179), .A4(new_n557), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n559), .A2(new_n567), .A3(KEYINPUT21), .A4(G169), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n570), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n552), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT23), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(new_n408), .A3(G20), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n585), .A2(new_n587), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n207), .B(G87), .C1(new_n342), .C2(new_n343), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT22), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT22), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n289), .A2(new_n594), .A3(new_n207), .A4(G87), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n591), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n597), .ZN(new_n599));
  AOI211_X1 g0399(.A(new_n599), .B(new_n591), .C1(new_n593), .C2(new_n595), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n254), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(G257), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n602));
  OAI211_X1 g0402(.A(G250), .B(new_n290), .C1(new_n342), .C2(new_n343), .ZN(new_n603));
  NAND2_X1  g0403(.A1(G33), .A2(G294), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n295), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n574), .A2(G264), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n479), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT82), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n352), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n487), .A2(new_n408), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n408), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT81), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT25), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n255), .B2(G107), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n615), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n601), .A2(new_n610), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n609), .B1(new_n608), .B2(new_n352), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(G190), .B2(new_n608), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n608), .A2(G179), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n309), .B2(new_n608), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n601), .A2(new_n618), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n619), .A2(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n510), .A2(new_n584), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n462), .A2(new_n626), .ZN(G372));
  NAND2_X1  g0427(.A1(new_n619), .A2(new_n621), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n541), .A2(new_n537), .A3(new_n538), .A4(new_n519), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n551), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT83), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT83), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n551), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n501), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n504), .A2(new_n309), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n480), .B1(new_n295), .B2(new_n469), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n311), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT77), .B1(new_n637), .B2(new_n352), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(new_n509), .A3(new_n501), .A4(new_n506), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n628), .A2(new_n634), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n623), .A2(new_n624), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n582), .A2(new_n581), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n570), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n551), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n639), .B1(new_n633), .B2(new_n631), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT26), .B1(new_n552), .B2(new_n639), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n462), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT84), .Z(new_n655));
  OAI21_X1  g0455(.A(new_n385), .B1(new_n380), .B2(new_n329), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(new_n391), .ZN(new_n657));
  INV_X1    g0457(.A(new_n452), .ZN(new_n658));
  INV_X1    g0458(.A(new_n414), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n658), .A2(new_n659), .B1(new_n458), .B2(new_n433), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n375), .A2(new_n390), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n313), .B1(new_n662), .B2(new_n308), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n655), .A2(new_n663), .ZN(G369));
  NAND3_X1  g0464(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  INV_X1    g0467(.A(G213), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(KEYINPUT85), .B(G343), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n579), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n645), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n583), .B2(new_n672), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n671), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n624), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n625), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n643), .A2(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n676), .B1(new_n644), .B2(new_n570), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n625), .A2(new_n682), .B1(new_n643), .B2(new_n671), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n210), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n575), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n513), .A2(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT86), .ZN(new_n690));
  OAI22_X1  g0490(.A1(new_n689), .A2(new_n690), .B1(new_n228), .B2(new_n687), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n690), .B2(new_n689), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT28), .Z(new_n693));
  NAND4_X1  g0493(.A1(new_n510), .A2(new_n584), .A3(new_n625), .A4(new_n671), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n557), .A2(G179), .A3(new_n479), .A4(new_n558), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT87), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n577), .A2(KEYINPUT87), .A3(G179), .A4(new_n557), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n548), .A2(new_n607), .A3(new_n606), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n697), .A2(new_n637), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n548), .A2(G179), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n504), .A2(new_n608), .A3(new_n559), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n637), .A2(KEYINPUT30), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n676), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(KEYINPUT31), .B(new_n676), .C1(new_n702), .C2(new_n707), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n694), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT88), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(KEYINPUT88), .A3(G330), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n653), .B2(new_n676), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n634), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n502), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n649), .B1(new_n552), .B2(new_n639), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT89), .B1(new_n648), .B2(KEYINPUT26), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT29), .B(new_n671), .C1(new_n724), .C2(new_n647), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n693), .B1(new_n728), .B2(G1), .ZN(G364));
  INV_X1    g0529(.A(G13), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n206), .B1(new_n731), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n686), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n225), .B1(G20), .B2(new_n309), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n207), .A2(G179), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G190), .A2(G200), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G159), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT32), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n207), .A2(new_n311), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n739), .ZN(new_n748));
  INV_X1    g0548(.A(new_n747), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n749), .A2(new_n365), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n289), .B1(new_n293), .B2(new_n748), .C1(new_n751), .C2(new_n318), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n749), .A2(G190), .A3(new_n352), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n738), .A2(new_n365), .A3(G200), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n215), .B1(new_n755), .B2(new_n408), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n365), .A2(G179), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n207), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n484), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n738), .A2(G190), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n217), .ZN(new_n761));
  NOR4_X1   g0561(.A1(new_n752), .A2(new_n756), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n747), .A2(G190), .A3(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT93), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n763), .A2(KEYINPUT93), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n746), .B(new_n762), .C1(new_n202), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n344), .B1(new_n751), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n748), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(G311), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n767), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G326), .ZN(new_n774));
  INV_X1    g0574(.A(G283), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n755), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G294), .ZN(new_n777));
  INV_X1    g0577(.A(G303), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n758), .A2(new_n777), .B1(new_n760), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n776), .B(new_n779), .C1(new_n753), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n743), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G329), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n772), .A2(new_n774), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n737), .B1(new_n768), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT92), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n736), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n685), .A2(new_n289), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G45), .B2(new_n228), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G45), .B2(new_n244), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT90), .ZN(new_n793));
  NAND2_X1  g0593(.A1(G355), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(G355), .A2(new_n793), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n210), .A2(new_n289), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G116), .B2(new_n210), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n797), .A2(KEYINPUT91), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(KEYINPUT91), .B2(new_n797), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n735), .B(new_n785), .C1(new_n789), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n788), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n674), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT95), .Z(new_n804));
  NOR2_X1   g0604(.A1(new_n674), .A2(G330), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n675), .A2(new_n805), .A3(new_n734), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  OAI21_X1  g0608(.A(new_n416), .B1(new_n403), .B2(new_n671), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n414), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n659), .A2(new_n671), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n653), .B2(new_n676), .ZN(new_n813));
  INV_X1    g0613(.A(new_n812), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n671), .B(new_n814), .C1(new_n647), .C2(new_n652), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n734), .B1(new_n717), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n717), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n736), .A2(new_n786), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n735), .B1(new_n293), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n755), .A2(new_n217), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n759), .A2(new_n821), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n822), .B1(new_n408), .B2(new_n760), .C1(new_n775), .C2(new_n754), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n289), .B1(new_n750), .B2(G294), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n561), .B2(new_n748), .C1(new_n743), .C2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n823), .B(new_n826), .C1(G303), .C2(new_n773), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n750), .A2(G143), .B1(G159), .B2(new_n771), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n247), .B2(new_n754), .C1(new_n767), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT34), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n755), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n344), .B1(new_n833), .B2(G68), .ZN(new_n834));
  INV_X1    g0634(.A(new_n758), .ZN(new_n835));
  INV_X1    g0635(.A(new_n760), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n835), .A2(G58), .B1(new_n836), .B2(G50), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n834), .B(new_n837), .C1(new_n743), .C2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n830), .B2(new_n831), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n827), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n820), .B1(new_n841), .B2(new_n737), .C1(new_n814), .C2(new_n787), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n818), .A2(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n731), .A2(new_n206), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n369), .A2(new_n324), .A3(new_n323), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n669), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n393), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n368), .A2(new_n374), .A3(KEYINPUT37), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n381), .B(new_n382), .C1(new_n385), .C2(new_n669), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n845), .B1(new_n385), .B2(new_n669), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n388), .A2(KEYINPUT74), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(new_n853), .A3(new_n373), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT38), .B1(new_n848), .B2(new_n856), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n856), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n381), .A2(new_n382), .A3(new_n669), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n388), .A3(new_n656), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n849), .A2(new_n850), .B1(new_n863), .B2(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT96), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n375), .A2(new_n865), .A3(new_n390), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n389), .B1(new_n853), .B2(new_n373), .ZN(new_n867));
  INV_X1    g0667(.A(new_n390), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT96), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n869), .A3(new_n657), .ZN(new_n870));
  INV_X1    g0670(.A(new_n862), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n864), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n861), .B1(new_n872), .B2(KEYINPUT38), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n860), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n458), .A2(new_n433), .A3(new_n671), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n815), .A2(new_n811), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n457), .A2(new_n455), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n449), .A2(new_n450), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n456), .B1(new_n881), .B2(G169), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n433), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n433), .A2(new_n676), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(new_n658), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n433), .B(new_n676), .C1(new_n458), .C2(new_n452), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n879), .A2(new_n888), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n889), .A2(new_n859), .B1(new_n657), .B2(new_n669), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n878), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n719), .B(new_n725), .C1(new_n460), .C2(new_n461), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n663), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n891), .B(new_n893), .Z(new_n894));
  INV_X1    g0694(.A(G330), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n812), .B1(new_n885), .B2(new_n886), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n708), .A2(KEYINPUT97), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n709), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n708), .A2(KEYINPUT97), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n711), .B(new_n694), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n896), .B(new_n900), .C1(new_n857), .C2(new_n858), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n901), .A2(KEYINPUT98), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT98), .B1(new_n901), .B2(new_n902), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n900), .A2(new_n896), .A3(KEYINPUT40), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n904), .A2(new_n906), .B1(new_n873), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n694), .A2(new_n711), .ZN(new_n909));
  INV_X1    g0709(.A(new_n899), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n709), .A3(new_n897), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n462), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n895), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n908), .B2(new_n912), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n844), .B1(new_n894), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n894), .B2(new_n914), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n917), .A2(G116), .A3(new_n226), .A4(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n228), .A2(new_n293), .A3(new_n336), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n215), .A2(G50), .ZN(new_n922));
  OAI211_X1 g0722(.A(G1), .B(new_n730), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n916), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT99), .ZN(G367));
  OAI21_X1  g0725(.A(new_n289), .B1(new_n751), .B2(new_n247), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(G50), .B2(new_n771), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n773), .A2(G143), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n833), .A2(G77), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n754), .B2(new_n744), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n758), .A2(new_n215), .B1(new_n760), .B2(new_n318), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n782), .A2(G137), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n927), .A2(new_n928), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n344), .B1(new_n775), .B2(new_n748), .C1(new_n751), .C2(new_n778), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n760), .A2(new_n561), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(KEYINPUT46), .B2(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n754), .A2(new_n777), .B1(new_n408), .B2(new_n758), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(G97), .B2(new_n833), .ZN(new_n939));
  XOR2_X1   g0739(.A(KEYINPUT106), .B(G317), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n782), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n773), .A2(G311), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n937), .A2(new_n939), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n936), .A2(KEYINPUT46), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT105), .Z(new_n945));
  OAI21_X1  g0745(.A(new_n934), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT47), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n737), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n947), .B2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n789), .B1(new_n210), .B2(new_n520), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n237), .A2(new_n685), .A3(new_n289), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n734), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT104), .Z(new_n953));
  AND2_X1   g0753(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n676), .A2(new_n522), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT100), .Z(new_n956));
  INV_X1    g0756(.A(new_n551), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT101), .ZN(new_n959));
  INV_X1    g0759(.A(new_n634), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(KEYINPUT101), .C1(new_n960), .C2(new_n956), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n954), .B1(new_n963), .B2(new_n802), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT103), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n623), .A2(new_n624), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n682), .A2(new_n628), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n680), .B2(new_n682), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(new_n675), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n717), .A2(new_n726), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n641), .B(new_n639), .C1(new_n501), .C2(new_n671), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n502), .A2(new_n676), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n643), .A2(new_n671), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n967), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n971), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n972), .A2(new_n973), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n683), .A2(new_n978), .A3(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n974), .A2(KEYINPUT44), .A3(new_n976), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n683), .B2(new_n978), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n681), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n980), .A2(new_n984), .A3(new_n681), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n965), .B1(new_n970), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n717), .A2(new_n726), .A3(new_n969), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n992), .A2(new_n989), .A3(KEYINPUT103), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n728), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n686), .B(new_n995), .Z(new_n996));
  AOI21_X1  g0796(.A(new_n733), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n978), .A2(new_n625), .A3(new_n682), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n639), .B1(new_n972), .B2(new_n966), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n998), .A2(KEYINPUT42), .B1(new_n671), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT42), .B2(new_n998), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n1001), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n962), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n681), .A2(new_n974), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n964), .B1(new_n997), .B2(new_n1010), .ZN(G387));
  AOI22_X1  g0811(.A1(new_n750), .A2(new_n940), .B1(G303), .B2(new_n771), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n825), .B2(new_n754), .C1(new_n767), .C2(new_n769), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT48), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n835), .A2(G283), .B1(new_n836), .B2(G294), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT49), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n782), .A2(G326), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n289), .B1(new_n833), .B2(G116), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n760), .A2(new_n293), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n754), .A2(new_n251), .B1(new_n755), .B2(new_n484), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(G159), .C2(new_n773), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n289), .B1(new_n215), .B2(new_n748), .C1(new_n751), .C2(new_n202), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n544), .A2(new_n545), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1028), .B1(new_n1030), .B2(new_n835), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1027), .B(new_n1031), .C1(new_n247), .C2(new_n743), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n737), .B1(new_n1024), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n234), .A2(new_n274), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT107), .ZN(new_n1035));
  XOR2_X1   g0835(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n1036));
  OR3_X1    g0836(.A1(new_n1036), .A2(G50), .A3(new_n251), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(G50), .B2(new_n251), .ZN(new_n1038));
  AOI21_X1  g0838(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1037), .A2(new_n688), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1035), .A2(new_n790), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n210), .A2(new_n289), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1041), .B1(G107), .B2(new_n210), .C1(new_n688), .C2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n735), .B(new_n1033), .C1(new_n789), .C2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n678), .A2(new_n679), .A3(new_n788), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1044), .A2(new_n1045), .B1(new_n733), .B2(new_n969), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n969), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n727), .A2(KEYINPUT109), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n686), .A3(new_n992), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT109), .B1(new_n727), .B2(new_n1047), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(G393));
  INV_X1    g0851(.A(KEYINPUT110), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n988), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n681), .B1(new_n980), .B2(new_n984), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n686), .B1(new_n1055), .B2(new_n970), .C1(new_n991), .C2(new_n993), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n974), .A2(new_n788), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n773), .A2(G317), .B1(G311), .B2(new_n750), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT52), .Z(new_n1059));
  OAI22_X1  g0859(.A1(new_n754), .A2(new_n778), .B1(new_n760), .B2(new_n775), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G116), .B2(new_n835), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n344), .B1(new_n748), .B2(new_n777), .C1(new_n408), .C2(new_n755), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n782), .B2(G322), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n773), .A2(G150), .B1(G159), .B2(new_n750), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n754), .A2(new_n202), .B1(new_n760), .B2(new_n215), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G77), .B2(new_n835), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n289), .B1(new_n748), .B2(new_n251), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n821), .B(new_n1071), .C1(new_n782), .C2(G143), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n737), .B1(new_n1064), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n790), .A2(new_n241), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n736), .B(new_n788), .C1(G97), .C2(new_n685), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n735), .B(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT112), .Z(new_n1078));
  AOI22_X1  g0878(.A1(new_n1055), .A2(new_n733), .B1(new_n1057), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1056), .A2(new_n1079), .ZN(G390));
  NAND2_X1  g0880(.A1(new_n889), .A2(new_n877), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT38), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n656), .B(KEYINPUT18), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n661), .B2(KEYINPUT96), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n862), .B1(new_n1084), .B2(new_n866), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1082), .B1(new_n1085), .B2(new_n864), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT39), .B1(new_n1086), .B2(new_n861), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n857), .A2(new_n858), .A3(new_n874), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1081), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n715), .A2(new_n716), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n814), .A3(new_n888), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n877), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1086), .B2(new_n861), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n671), .B(new_n810), .C1(new_n724), .C2(new_n647), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n887), .B1(new_n1094), .B2(new_n811), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT113), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n873), .A2(new_n877), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT113), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n1095), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1089), .B(new_n1091), .C1(new_n1097), .C2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1093), .A2(new_n1096), .A3(KEYINPUT113), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1099), .B1(new_n1098), .B2(new_n1095), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1102), .A2(new_n1103), .B1(new_n876), .B2(new_n1081), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n895), .B1(new_n911), .B2(new_n909), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1105), .A2(new_n896), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1101), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n888), .B1(new_n1090), .B2(new_n814), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n879), .B1(new_n1109), .B2(new_n1106), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1094), .A2(new_n811), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1105), .A2(new_n814), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n887), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1091), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1105), .B1(new_n460), .B2(new_n461), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n892), .A2(new_n663), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n687), .B1(new_n1108), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1117), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n1101), .C1(new_n1104), .C2(new_n1107), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n819), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n734), .B1(new_n322), .B2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT114), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n782), .A2(G125), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n755), .A2(new_n202), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n289), .B1(new_n751), .B2(new_n838), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(G159), .C2(new_n835), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n760), .A2(new_n247), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n773), .A2(G128), .ZN(new_n1133));
  AND4_X1   g0933(.A1(new_n1127), .A2(new_n1130), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n753), .A2(G137), .B1(new_n771), .B2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT115), .Z(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n289), .B(new_n761), .C1(G116), .C2(new_n750), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n835), .A2(G77), .B1(new_n833), .B2(G68), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n777), .C2(new_n743), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n753), .A2(G107), .B1(G97), .B2(new_n771), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT116), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n775), .B2(new_n767), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1144), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(KEYINPUT116), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1134), .A2(new_n1139), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1126), .B1(new_n1151), .B2(new_n736), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n876), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n787), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT117), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1101), .B(new_n733), .C1(new_n1104), .C2(new_n1107), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1123), .A2(new_n1155), .A3(new_n1156), .ZN(G378));
  AOI21_X1  g0957(.A(new_n895), .B1(new_n907), .B2(new_n873), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n903), .B2(new_n905), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n268), .A2(new_n669), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT55), .Z(new_n1161));
  XNOR2_X1  g0961(.A(new_n315), .B(new_n1161), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1158), .B(new_n1166), .C1(new_n903), .C2(new_n905), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1165), .A2(new_n891), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n891), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n733), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n735), .B1(new_n202), .B2(new_n819), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n767), .A2(new_n561), .B1(new_n215), .B2(new_n758), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT118), .Z(new_n1173));
  NAND3_X1  g0973(.A1(new_n344), .A2(new_n273), .A3(new_n275), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1174), .B(new_n1025), .C1(G107), .C2(new_n750), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n318), .B2(new_n755), .C1(new_n484), .C2(new_n754), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n743), .A2(new_n775), .B1(new_n1029), .B2(new_n748), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1173), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1178), .A2(KEYINPUT58), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(KEYINPUT58), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n773), .A2(G125), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n753), .A2(G132), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n750), .A2(G128), .B1(G137), .B2(new_n771), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n835), .A2(G150), .B1(new_n836), .B2(new_n1136), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n782), .A2(G124), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G33), .B(G41), .C1(new_n833), .C2(G159), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1174), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1191));
  AND4_X1   g0991(.A1(new_n1179), .A2(new_n1180), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1171), .B1(new_n737), .B2(new_n1192), .C1(new_n1166), .C2(new_n787), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1170), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT57), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1122), .A2(new_n1118), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n686), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n891), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1165), .A2(new_n891), .A3(new_n1167), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1122), .A2(new_n1118), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1194), .B1(new_n1197), .B2(new_n1204), .ZN(G375));
  AOI21_X1  g1005(.A(new_n732), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT120), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT120), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n289), .B1(new_n748), .B2(new_n247), .C1(new_n318), .C2(new_n755), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n758), .A2(new_n202), .B1(new_n760), .B2(new_n744), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(new_n782), .C2(G128), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT121), .Z(new_n1212));
  AOI22_X1  g1012(.A1(G137), .A2(new_n750), .B1(new_n753), .B2(new_n1136), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n838), .C2(new_n767), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n929), .B1(new_n484), .B2(new_n760), .C1(new_n754), .C2(new_n561), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G294), .B2(new_n773), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1030), .A2(new_n835), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n782), .A2(G303), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n344), .B1(new_n751), .B2(new_n775), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G107), .B2(new_n771), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n737), .B1(new_n1214), .B2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n735), .B(new_n1222), .C1(new_n215), .C2(new_n819), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n786), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n888), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1207), .A2(new_n1208), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1110), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1119), .A2(new_n996), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(G381));
  INV_X1    g1030(.A(G375), .ZN(new_n1231));
  OR2_X1    g1031(.A1(G390), .A2(G384), .ZN(new_n1232));
  OR2_X1    g1032(.A1(G393), .A2(G396), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(G381), .A2(new_n1232), .A3(G387), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1231), .A2(new_n1234), .A3(new_n1236), .ZN(G407));
  NOR2_X1   g1037(.A1(new_n670), .A2(new_n668), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1231), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(G407), .A2(new_n1239), .A3(G213), .ZN(G409));
  INV_X1    g1040(.A(G390), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(G387), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n964), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n970), .A2(new_n990), .A3(new_n965), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT103), .B1(new_n992), .B2(new_n989), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n727), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n996), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n732), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1243), .B1(new_n1248), .B2(new_n1009), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(G390), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(G393), .B(new_n807), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1242), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT125), .B1(new_n1249), .B2(G390), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1255), .A2(new_n1252), .B1(new_n1242), .B2(new_n1250), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G378), .B(new_n1194), .C1(new_n1197), .C2(new_n1204), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1202), .A2(new_n996), .A3(new_n1203), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1170), .A2(new_n1193), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1236), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1238), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  XOR2_X1   g1063(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n1264));
  NAND2_X1  g1064(.A1(new_n1119), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1228), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n686), .B1(new_n1228), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  OR2_X1    g1070(.A1(G384), .A2(KEYINPUT123), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1227), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(G384), .B(KEYINPUT123), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1268), .B1(new_n1265), .B2(new_n1228), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(new_n1274), .B2(new_n1226), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1238), .A2(G2897), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1272), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1257), .B(new_n1258), .C1(new_n1263), .C2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1238), .B(new_n1276), .C1(new_n1259), .C2(new_n1262), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT63), .B1(new_n1284), .B2(KEYINPUT124), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1276), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1263), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT124), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1283), .A2(new_n1285), .A3(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1263), .A2(new_n1286), .A3(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1258), .B1(new_n1263), .B2(new_n1281), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT126), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT62), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1263), .B2(new_n1286), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1293), .A2(new_n1294), .A3(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1291), .B1(new_n1298), .B2(new_n1257), .ZN(G405));
  INV_X1    g1099(.A(new_n1256), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1253), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G375), .A2(new_n1236), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(KEYINPUT127), .A3(new_n1259), .A4(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1259), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1286), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1257), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1303), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1306), .B1(new_n1303), .B2(new_n1307), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(G402));
endmodule


