//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  AND3_X1   g004(.A1(new_n190), .A2(KEYINPUT1), .A3(G146), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n191), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n193), .A3(new_n194), .ZN(new_n199));
  AOI21_X1  g013(.A(G125), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT0), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n196), .A3(KEYINPUT64), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(KEYINPUT0), .B2(G128), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n205), .A2(new_n207), .B1(KEYINPUT0), .B2(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n203), .B1(new_n208), .B2(new_n201), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n200), .B1(G125), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G224), .ZN(new_n211));
  OR3_X1    g025(.A1(new_n211), .A2(KEYINPUT85), .A3(G953), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT85), .B1(new_n211), .B2(G953), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n189), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n197), .A2(new_n199), .ZN(new_n216));
  MUX2_X1   g030(.A(new_n216), .B(new_n209), .S(G125), .Z(new_n217));
  INV_X1    g031(.A(new_n214), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(KEYINPUT86), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n211), .A2(G953), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(KEYINPUT84), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(KEYINPUT84), .B2(new_n221), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n215), .A2(new_n219), .B1(new_n210), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G116), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G119), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n226), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n232), .A2(G116), .A3(new_n225), .A4(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n234), .A3(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n226), .A2(new_n228), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT2), .B(G113), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G107), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT74), .A3(G104), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n240), .A2(G104), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G101), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n246), .A2(new_n240), .A3(KEYINPUT74), .A4(G104), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n242), .A2(new_n244), .A3(new_n245), .A4(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G104), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(G107), .ZN(new_n250));
  OAI21_X1  g064(.A(G101), .B1(new_n250), .B2(new_n243), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n239), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n242), .A2(new_n247), .A3(new_n244), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G101), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT75), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT75), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n254), .A2(new_n258), .A3(new_n255), .A4(G101), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G116), .B(G119), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(new_n237), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n255), .B1(new_n254), .B2(G101), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(new_n248), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n253), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G110), .B(G122), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n238), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n234), .A2(G113), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT82), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n269), .A2(new_n270), .B1(KEYINPUT5), .B2(new_n261), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n234), .A2(KEYINPUT82), .A3(G113), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(new_n252), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n266), .B(KEYINPUT8), .ZN(new_n275));
  INV_X1    g089(.A(new_n252), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(new_n239), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT83), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n277), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT83), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n279), .B(new_n280), .C1(new_n252), .C2(new_n273), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n224), .A2(new_n267), .A3(new_n278), .A4(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n220), .B(KEYINPUT81), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n217), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n266), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n287), .B(new_n253), .C1(new_n260), .C2(new_n264), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(KEYINPUT80), .ZN(new_n290));
  OAI22_X1  g104(.A1(new_n288), .A2(new_n289), .B1(new_n265), .B2(new_n290), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n265), .A2(new_n289), .A3(new_n290), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n286), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n188), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n286), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n260), .A2(new_n264), .ZN(new_n297));
  INV_X1    g111(.A(new_n253), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n290), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n267), .A2(KEYINPUT6), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n296), .B1(new_n301), .B2(new_n292), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n302), .A2(new_n283), .A3(new_n187), .A4(new_n282), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G469), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n205), .A2(new_n207), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n201), .B1(new_n308), .B2(new_n202), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n201), .A2(new_n202), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT67), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n312), .B(new_n203), .C1(new_n208), .C2(new_n201), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n263), .A2(new_n248), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n260), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT65), .A2(G131), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT65), .A2(G131), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT11), .ZN(new_n320));
  INV_X1    g134(.A(G134), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(G137), .ZN(new_n322));
  INV_X1    g136(.A(G137), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT11), .A3(G134), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(G137), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n319), .A2(new_n322), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n322), .A2(new_n324), .A3(new_n328), .A4(new_n325), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n329), .A2(G131), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n327), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n199), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n201), .A2(KEYINPUT76), .A3(new_n198), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n197), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n248), .A3(new_n251), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT10), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(new_n197), .B2(new_n199), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n338), .A2(new_n339), .B1(new_n276), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n316), .A2(new_n333), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n332), .A2(G131), .A3(new_n329), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT77), .B1(new_n343), .B2(new_n326), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n345));
  OAI22_X1  g159(.A1(new_n201), .A2(G128), .B1(new_n345), .B2(new_n194), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT76), .B1(new_n201), .B2(new_n198), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n252), .B1(new_n348), .B2(new_n336), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n216), .B1(new_n248), .B2(new_n251), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n344), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT12), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT12), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(new_n344), .C1(new_n349), .C2(new_n350), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n342), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G110), .B(G140), .ZN(new_n356));
  INV_X1    g170(.A(G953), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n357), .A2(G227), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n356), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n316), .A2(new_n341), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n343), .A2(new_n326), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n359), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n342), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n307), .B1(new_n366), .B2(new_n283), .ZN(new_n367));
  XOR2_X1   g181(.A(KEYINPUT72), .B(G902), .Z(new_n368));
  AOI21_X1  g182(.A(new_n364), .B1(new_n363), .B2(new_n342), .ZN(new_n369));
  AND4_X1   g183(.A1(new_n342), .A2(new_n352), .A3(new_n354), .A4(new_n364), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n307), .B(new_n368), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT78), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n316), .A2(new_n333), .A3(new_n341), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n333), .B1(new_n316), .B2(new_n341), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n359), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n342), .A2(new_n352), .A3(new_n354), .A4(new_n364), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n378), .A2(KEYINPUT78), .A3(new_n307), .A4(new_n368), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n367), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT9), .B(G234), .ZN(new_n381));
  OAI21_X1  g195(.A(G221), .B1(new_n381), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n306), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n357), .A3(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n190), .ZN(new_n388));
  NOR2_X1   g202(.A1(G237), .A2(G953), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(G143), .A3(G214), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT18), .A2(G131), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(KEYINPUT18), .A3(G131), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n192), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G113), .B(G122), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n249), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n317), .A2(new_n318), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n391), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT17), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n388), .A2(new_n319), .A3(new_n390), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n401), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT16), .ZN(new_n407));
  INV_X1    g221(.A(G140), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(G125), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(G125), .ZN(new_n410));
  INV_X1    g224(.A(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n409), .B1(new_n413), .B2(new_n407), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n192), .ZN(new_n415));
  OAI211_X1 g229(.A(G146), .B(new_n409), .C1(new_n413), .C2(new_n407), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n406), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n398), .B(new_n400), .C1(new_n405), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT87), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n420), .A2(new_n415), .A3(new_n416), .A4(new_n406), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n400), .A4(new_n398), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n396), .B(KEYINPUT19), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n192), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n402), .A2(new_n404), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n416), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n398), .ZN(new_n429));
  INV_X1    g243(.A(new_n400), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n434), .B(KEYINPUT88), .Z(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT20), .A4(new_n436), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n433), .A2(KEYINPUT20), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(KEYINPUT20), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n419), .A2(new_n423), .B1(new_n430), .B2(new_n429), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n438), .B(new_n439), .C1(new_n440), .C2(new_n435), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n400), .B1(new_n421), .B2(new_n398), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(new_n419), .B2(new_n423), .ZN(new_n443));
  OAI21_X1  g257(.A(G475), .B1(new_n443), .B2(G902), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n437), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(G128), .A3(new_n190), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n190), .A2(G128), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n196), .A2(G143), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n448), .B(G134), .C1(new_n451), .C2(new_n447), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT91), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT91), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n321), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n227), .A2(G122), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G116), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n460), .A2(new_n240), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n240), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n452), .B(new_n456), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT93), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT91), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT91), .B1(new_n449), .B2(new_n450), .ZN(new_n466));
  OAI21_X1  g280(.A(G134), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n456), .ZN(new_n468));
  OAI211_X1 g282(.A(KEYINPUT92), .B(KEYINPUT14), .C1(new_n458), .C2(G116), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT92), .B1(new_n457), .B2(KEYINPUT14), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n459), .B1(new_n457), .B2(KEYINPUT14), .ZN(new_n473));
  OAI21_X1  g287(.A(G107), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n461), .ZN(new_n475));
  AND4_X1   g289(.A1(new_n464), .A2(new_n468), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n461), .B1(new_n467), .B2(new_n456), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n464), .B1(new_n477), .B2(new_n474), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n463), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G217), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n381), .A2(new_n480), .A3(G953), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT94), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n482), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n484), .B(new_n463), .C1(new_n476), .C2(new_n478), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(KEYINPUT95), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n479), .A2(new_n487), .A3(new_n482), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n368), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(G478), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(G478), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n486), .A2(new_n368), .A3(new_n488), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n446), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G952), .ZN(new_n496));
  AOI211_X1 g310(.A(G953), .B(new_n496), .C1(G234), .C2(G237), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n357), .B(new_n368), .C1(G234), .C2(G237), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT21), .B(G898), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n384), .A2(new_n385), .A3(new_n495), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n373), .A2(new_n379), .ZN(new_n503));
  INV_X1    g317(.A(new_n367), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n305), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n295), .B2(new_n303), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n505), .A2(new_n382), .A3(new_n507), .A4(new_n501), .ZN(new_n508));
  INV_X1    g322(.A(new_n495), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT96), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n321), .A2(G137), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n323), .A2(G134), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n331), .B2(new_n401), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n514), .A2(new_n515), .B1(new_n197), .B2(new_n199), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n326), .A2(KEYINPUT68), .A3(new_n513), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n314), .A2(new_n362), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT28), .B1(new_n518), .B2(new_n262), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n520));
  INV_X1    g334(.A(new_n262), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n515), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n522), .A2(new_n517), .A3(new_n216), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n311), .A2(new_n313), .B1(new_n343), .B2(new_n326), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n206), .A2(KEYINPUT0), .A3(G128), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT64), .B1(new_n204), .B2(new_n196), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n202), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n195), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n312), .B1(new_n529), .B2(new_n203), .ZN(new_n530));
  INV_X1    g344(.A(new_n313), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n362), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n516), .A2(new_n517), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n262), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n520), .B1(new_n525), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT71), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n519), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n523), .A2(new_n524), .A3(new_n521), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n262), .B1(new_n532), .B2(new_n533), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT28), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT71), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n389), .A2(G210), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT27), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n537), .A2(new_n541), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n534), .A2(new_n520), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n518), .A2(KEYINPUT28), .A3(new_n262), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n216), .A2(new_n326), .A3(new_n513), .ZN(new_n552));
  INV_X1    g366(.A(new_n209), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n552), .B1(new_n333), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n521), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n550), .A2(new_n545), .A3(new_n551), .A4(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n557), .B(new_n552), .C1(new_n333), .C2(new_n553), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n518), .B2(new_n557), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n538), .B1(new_n559), .B2(new_n521), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n547), .B(new_n556), .C1(new_n560), .C2(new_n545), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n549), .A2(new_n368), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G472), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n521), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n534), .A2(new_n545), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT31), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT30), .B1(new_n523), .B2(new_n524), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n262), .B1(new_n569), .B2(new_n558), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n570), .B2(new_n565), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n546), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(KEYINPUT69), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n567), .A2(new_n571), .B1(new_n546), .B2(new_n573), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n577), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n563), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n480), .B1(new_n368), .B2(G234), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n415), .A2(new_n416), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n225), .A2(G128), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n225), .A2(G128), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(KEYINPUT23), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT24), .B(G110), .Z(new_n591));
  XNOR2_X1  g405(.A(G119), .B(G128), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n590), .A2(G110), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT73), .B(G110), .Z(new_n595));
  OAI22_X1  g409(.A1(new_n590), .A2(new_n595), .B1(new_n591), .B2(new_n592), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(new_n416), .C1(G146), .C2(new_n413), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT22), .B(G137), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n357), .A2(G221), .A3(G234), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n594), .B2(new_n597), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT25), .B1(new_n605), .B2(new_n368), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT25), .ZN(new_n607));
  INV_X1    g421(.A(new_n368), .ZN(new_n608));
  NOR4_X1   g422(.A1(new_n603), .A2(new_n604), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n585), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n585), .A2(G902), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n584), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n502), .A2(new_n510), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  OAI21_X1  g432(.A(G472), .B1(new_n582), .B2(new_n608), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n575), .A2(new_n578), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n384), .A2(new_n615), .A3(new_n501), .A4(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n486), .A2(new_n623), .A3(new_n488), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n483), .A2(KEYINPUT33), .A3(new_n485), .ZN(new_n625));
  INV_X1    g439(.A(G478), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n608), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n489), .A2(new_n626), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n629), .B1(new_n628), .B2(new_n630), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n446), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n622), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND2_X1  g450(.A1(new_n437), .A2(new_n441), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT98), .ZN(new_n638));
  INV_X1    g452(.A(new_n444), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n491), .B2(new_n493), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n622), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G107), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR2_X1   g459(.A1(new_n602), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n598), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n611), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n610), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n502), .A2(new_n510), .A3(new_n621), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  AND2_X1   g466(.A1(new_n584), .A2(new_n649), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n497), .B1(new_n498), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n638), .A2(new_n640), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n653), .A2(new_n657), .A3(new_n384), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  XNOR2_X1  g473(.A(new_n304), .B(KEYINPUT38), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n560), .A2(new_n546), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n525), .A2(new_n534), .A3(new_n546), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n283), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n579), .A2(new_n583), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n445), .B1(new_n491), .B2(new_n493), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n649), .A2(new_n506), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n660), .A2(new_n665), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT100), .Z(new_n669));
  NOR2_X1   g483(.A1(new_n380), .A2(new_n383), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n655), .B(KEYINPUT39), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT40), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT101), .B(G143), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G45));
  OAI211_X1 g490(.A(new_n446), .B(new_n656), .C1(new_n631), .C2(new_n632), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n653), .A3(new_n384), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  AOI21_X1  g494(.A(new_n307), .B1(new_n378), .B2(new_n368), .ZN(new_n681));
  AOI211_X1 g495(.A(new_n383), .B(new_n681), .C1(new_n373), .C2(new_n379), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n682), .A2(new_n584), .A3(new_n615), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n507), .A2(new_n501), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n633), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT41), .B(G113), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT102), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n686), .B(new_n688), .ZN(G15));
  NAND3_X1  g503(.A1(new_n682), .A2(new_n584), .A3(new_n615), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n638), .A2(new_n507), .A3(new_n501), .A4(new_n640), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n227), .ZN(G18));
  AND4_X1   g507(.A1(new_n445), .A2(new_n491), .A3(new_n493), .A4(new_n501), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n584), .A2(new_n694), .A3(new_n649), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n682), .A2(new_n507), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n225), .ZN(G21));
  NAND3_X1  g512(.A1(new_n507), .A2(new_n446), .A3(new_n494), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT103), .B(G472), .Z(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n582), .B2(new_n608), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n567), .A2(new_n571), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n545), .B1(new_n537), .B2(new_n541), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n578), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n701), .A2(new_n704), .A3(new_n615), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n681), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n503), .A2(new_n382), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n500), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NOR2_X1   g525(.A1(new_n708), .A2(new_n306), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n628), .A2(new_n630), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT97), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n445), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n701), .A2(new_n704), .A3(new_n649), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n712), .A2(new_n716), .A3(new_n717), .A4(new_n656), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n720));
  AOI21_X1  g534(.A(G902), .B1(new_n360), .B2(new_n365), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n720), .B1(new_n721), .B2(new_n307), .ZN(new_n722));
  INV_X1    g536(.A(new_n366), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n720), .A2(new_n307), .A3(G902), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n722), .A2(new_n725), .B1(new_n373), .B2(new_n379), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n295), .A2(new_n303), .A3(new_n305), .ZN(new_n728));
  NOR4_X1   g542(.A1(new_n726), .A2(new_n727), .A3(new_n383), .A4(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT32), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n582), .B2(new_n577), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n563), .A2(new_n579), .A3(new_n731), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n732), .A2(KEYINPUT105), .A3(new_n615), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT105), .B1(new_n732), .B2(new_n615), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n729), .B(new_n678), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n722), .A2(new_n725), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n383), .B1(new_n736), .B2(new_n503), .ZN(new_n737));
  INV_X1    g551(.A(new_n728), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n584), .A3(new_n615), .A4(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n727), .B1(new_n739), .B2(new_n677), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n735), .A2(KEYINPUT106), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT106), .B1(new_n735), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  NOR3_X1   g558(.A1(new_n726), .A2(new_n383), .A3(new_n728), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n616), .A2(new_n745), .A3(new_n657), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n631), .A2(new_n632), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n446), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n749), .C2(new_n446), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n621), .B1(new_n610), .B2(new_n648), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n756), .A2(KEYINPUT44), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(KEYINPUT44), .A3(new_n755), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n723), .A2(KEYINPUT45), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n307), .B1(new_n366), .B2(new_n760), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n759), .A2(new_n761), .B1(G469), .B2(G902), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT46), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(KEYINPUT46), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n503), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n382), .A3(new_n671), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n728), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n757), .A2(new_n758), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  AND3_X1   g583(.A1(new_n765), .A2(KEYINPUT47), .A3(new_n382), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT47), .B1(new_n765), .B2(new_n382), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n677), .A2(new_n584), .A3(new_n615), .A4(new_n728), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT108), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  INV_X1    g591(.A(new_n705), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n752), .A2(new_n497), .A3(new_n778), .A4(new_n753), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n660), .A2(new_n305), .A3(new_n708), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT50), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n708), .A2(new_n728), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n752), .A2(new_n497), .A3(new_n753), .A4(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(KEYINPUT114), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(KEYINPUT114), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n717), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n497), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n665), .A2(new_n614), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(new_n445), .A3(new_n783), .A4(new_n749), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n782), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n681), .B1(new_n373), .B2(new_n379), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n383), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n728), .B1(new_n772), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n779), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT51), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n791), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n785), .A2(new_n786), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n733), .A2(new_n734), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT48), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT48), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n789), .A2(new_n716), .A3(new_n783), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(G952), .A3(new_n357), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n795), .B2(new_n712), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n798), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n791), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n796), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n791), .A2(new_n811), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n735), .A2(new_n740), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT106), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n735), .A2(new_n740), .A3(KEYINPUT106), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n678), .A2(new_n745), .A3(new_n717), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n649), .A2(new_n444), .A3(new_n656), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n494), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(new_n638), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(new_n584), .A3(new_n670), .A4(new_n738), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n824), .A3(new_n746), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n818), .A2(new_n819), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n699), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n610), .A2(new_n648), .A3(new_n656), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT112), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n828), .A2(new_n665), .A3(new_n737), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n679), .A2(new_n658), .A3(new_n718), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n384), .B(new_n653), .C1(new_n678), .C2(new_n657), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n718), .A4(new_n831), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n827), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n691), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n584), .A2(new_n694), .A3(new_n649), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n683), .A2(new_n839), .B1(new_n840), .B2(new_n712), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n683), .A2(new_n685), .B1(new_n709), .B2(new_n706), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n306), .A2(new_n500), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n716), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n701), .A2(new_n704), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n615), .A3(new_n507), .A4(new_n666), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n682), .A2(new_n501), .ZN(new_n849));
  OAI22_X1  g663(.A1(new_n846), .A2(new_n690), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n690), .A2(new_n691), .B1(new_n695), .B2(new_n696), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT110), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n844), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n633), .A2(KEYINPUT111), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT111), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n855), .B(new_n446), .C1(new_n631), .C2(new_n632), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n640), .A2(new_n437), .A3(new_n441), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n622), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n617), .A3(new_n650), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT53), .B1(new_n838), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n861), .A2(new_n617), .A3(new_n650), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n850), .A2(new_n851), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n866), .A2(KEYINPUT113), .A3(new_n816), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT113), .B1(new_n866), .B2(new_n816), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n825), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n833), .A3(new_n836), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n864), .A2(new_n873), .A3(KEYINPUT54), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n502), .A2(new_n510), .A3(new_n616), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n622), .B1(new_n857), .B2(new_n858), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n650), .A3(new_n852), .A4(new_n844), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n878), .A2(new_n837), .A3(new_n827), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT53), .ZN(new_n880));
  INV_X1    g694(.A(new_n837), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n741), .A2(new_n742), .A3(new_n825), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n863), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n870), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n874), .B1(KEYINPUT54), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n809), .A2(new_n815), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT116), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n496), .A2(new_n357), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(KEYINPUT116), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n750), .A2(new_n615), .A3(new_n382), .A4(new_n305), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n660), .A2(new_n665), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n792), .B(KEYINPUT49), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT109), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n895), .B(new_n896), .C1(new_n892), .C2(new_n897), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n890), .A2(new_n891), .B1(new_n894), .B2(new_n898), .ZN(G75));
  NOR2_X1   g713(.A1(new_n357), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n871), .A2(new_n833), .A3(new_n836), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n902), .B(new_n865), .C1(new_n868), .C2(new_n867), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n368), .B1(new_n884), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT56), .B1(new_n904), .B2(new_n188), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n291), .A2(new_n286), .A3(new_n293), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n906), .A2(new_n302), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n901), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n905), .B2(new_n908), .ZN(G51));
  NAND2_X1  g724(.A1(G469), .A2(G902), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT57), .Z(new_n912));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n884), .B2(new_n903), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n874), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n378), .ZN(new_n917));
  INV_X1    g731(.A(new_n912), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT54), .B1(new_n864), .B2(new_n873), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n913), .B(new_n903), .C1(new_n879), .C2(KEYINPUT53), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n378), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT117), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n904), .A2(new_n759), .A3(new_n761), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n917), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n901), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT118), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(KEYINPUT118), .A3(new_n901), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(G54));
  AND3_X1   g744(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n901), .B1(new_n931), .B2(new_n432), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n432), .B2(new_n931), .ZN(G60));
  NAND2_X1  g747(.A1(new_n624), .A2(new_n625), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT119), .Z(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT59), .Z(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n874), .B2(new_n914), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n901), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n940), .A2(KEYINPUT120), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n935), .B1(new_n886), .B2(new_n937), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(KEYINPUT120), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n864), .B2(new_n873), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n603), .B2(new_n604), .ZN(new_n948));
  INV_X1    g762(.A(new_n647), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n948), .B(new_n901), .C1(new_n949), .C2(new_n947), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT121), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT61), .ZN(G66));
  NOR2_X1   g766(.A1(new_n863), .A2(G953), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT122), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n499), .B2(new_n211), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n291), .B(new_n293), .C1(G898), .C2(new_n357), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  XNOR2_X1  g772(.A(new_n559), .B(new_n425), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT123), .Z(new_n960));
  AND2_X1   g774(.A1(new_n776), .A2(new_n768), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n674), .A2(new_n718), .A3(new_n834), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n672), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n859), .A2(new_n616), .A3(new_n965), .A4(new_n738), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n961), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(G953), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n357), .A2(G900), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n800), .A2(new_n828), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(new_n766), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n834), .A2(new_n718), .A3(new_n746), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n776), .A2(new_n768), .A3(new_n743), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n969), .B1(new_n974), .B2(new_n357), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n959), .B1(new_n975), .B2(KEYINPUT124), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n968), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT125), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n960), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n357), .B1(G227), .B2(G900), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n968), .B(new_n983), .C1(new_n976), .C2(new_n977), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n974), .B2(new_n878), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n546), .A3(new_n560), .ZN(new_n989));
  INV_X1    g803(.A(new_n661), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n560), .A2(new_n546), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT127), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n900), .B1(new_n885), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n961), .A2(new_n863), .A3(new_n964), .A4(new_n966), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n990), .B1(new_n996), .B2(new_n987), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(KEYINPUT126), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(G57));
endmodule


