//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT71), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT64), .A2(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(G143), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n193), .A2(new_n196), .A3(G143), .A4(new_n194), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n190), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n194), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT64), .A2(G146), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n204), .A2(new_n205), .A3(new_n197), .ZN(new_n206));
  OAI21_X1  g020(.A(G128), .B1(new_n206), .B2(new_n202), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n197), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n197), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT68), .B1(new_n207), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n190), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n210), .B1(new_n208), .B2(new_n197), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n203), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G134), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G134), .ZN(new_n223));
  INV_X1    g037(.A(G134), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n221), .B1(new_n226), .B2(KEYINPUT67), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(G134), .ZN(new_n229));
  AOI21_X1  g043(.A(G137), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n219), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(new_n229), .A3(G137), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n224), .A2(G137), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n228), .A2(new_n229), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT11), .B1(new_n239), .B2(new_n220), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n238), .A2(new_n240), .A3(G131), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(G131), .B1(new_n238), .B2(new_n240), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT66), .B(G134), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n234), .B1(new_n244), .B2(G137), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n236), .B1(new_n244), .B2(G137), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n219), .B(new_n245), .C1(new_n246), .C2(new_n234), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n209), .B2(new_n211), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n201), .B2(KEYINPUT0), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n218), .A2(new_n242), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g066(.A(G116), .B(G119), .Z(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT2), .B(G113), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT28), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n248), .A2(new_n251), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n207), .A2(KEYINPUT68), .A3(new_n212), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n216), .B1(new_n214), .B2(new_n215), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n259), .A2(new_n260), .B1(new_n202), .B2(new_n201), .ZN(new_n261));
  OAI22_X1  g075(.A1(new_n230), .A2(new_n231), .B1(G134), .B2(new_n220), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n263));
  OAI21_X1  g077(.A(G131), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n247), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n258), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n255), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n258), .B(new_n256), .C1(new_n261), .C2(new_n265), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n257), .B1(new_n269), .B2(KEYINPUT28), .ZN(new_n270));
  INV_X1    g084(.A(G237), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G210), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n273), .B(KEYINPUT27), .Z(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n274), .B(new_n275), .Z(new_n276));
  OAI21_X1  g090(.A(new_n189), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n276), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n267), .B2(new_n268), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT71), .B(new_n278), .C1(new_n280), .C2(new_n257), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  INV_X1    g096(.A(new_n268), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n266), .A2(KEYINPUT30), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n258), .B(new_n285), .C1(new_n261), .C2(new_n265), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n283), .B1(new_n287), .B2(new_n255), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n282), .B1(new_n288), .B2(new_n276), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n277), .A2(new_n281), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n256), .B1(new_n284), .B2(new_n286), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n293));
  NOR4_X1   g107(.A1(new_n292), .A2(new_n283), .A3(new_n278), .A4(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n286), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n218), .A2(new_n242), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n285), .B1(new_n296), .B2(new_n258), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n255), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n268), .A3(new_n276), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT31), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n294), .B1(new_n300), .B2(KEYINPUT69), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n188), .B1(new_n291), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT72), .B1(new_n302), .B2(KEYINPUT32), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(KEYINPUT32), .ZN(new_n304));
  INV_X1    g118(.A(new_n257), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n278), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n307), .B(new_n309), .C1(new_n270), .C2(new_n306), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(KEYINPUT74), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n270), .A2(new_n276), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n316), .B(new_n308), .C1(new_n288), .C2(new_n276), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G472), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n299), .A2(new_n290), .A3(KEYINPUT31), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n256), .B1(new_n296), .B2(new_n258), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT28), .B1(new_n283), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n305), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT71), .B1(new_n323), .B2(new_n278), .ZN(new_n324));
  INV_X1    g138(.A(new_n281), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n320), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n292), .A2(new_n283), .A3(new_n278), .ZN(new_n327));
  INV_X1    g141(.A(new_n293), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n289), .B2(new_n290), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n187), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT72), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT32), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n303), .A2(new_n304), .A3(new_n319), .A4(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G234), .ZN(new_n336));
  OAI21_X1  g150(.A(G217), .B1(new_n336), .B2(G902), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT75), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n340), .A2(G140), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT16), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT79), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n340), .A3(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(KEYINPUT77), .A2(G140), .ZN(new_n349));
  NOR2_X1   g163(.A1(KEYINPUT77), .A2(G140), .ZN(new_n350));
  OAI21_X1  g164(.A(G125), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT78), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(G125), .C1(new_n349), .C2(new_n350), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n348), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n343), .B1(new_n355), .B2(new_n342), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G146), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n192), .B(new_n343), .C1(new_n355), .C2(new_n342), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT23), .B1(new_n190), .B2(G119), .ZN(new_n360));
  INV_X1    g174(.A(G119), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n360), .B(KEYINPUT76), .C1(new_n361), .C2(G128), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(G128), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(KEYINPUT23), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G110), .ZN(new_n368));
  XOR2_X1   g182(.A(G119), .B(G128), .Z(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT24), .B(G110), .ZN(new_n370));
  OAI22_X1  g184(.A1(new_n367), .A2(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n359), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n341), .A2(new_n344), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(new_n208), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n367), .A2(new_n368), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n369), .A2(new_n370), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n357), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT22), .B(G137), .ZN(new_n380));
  INV_X1    g194(.A(G221), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n381), .A2(new_n336), .A3(G953), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n380), .B(new_n382), .Z(new_n383));
  NAND3_X1  g197(.A1(new_n373), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n383), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n378), .A2(new_n357), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n371), .B1(new_n357), .B2(new_n358), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n388), .A3(new_n311), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT25), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n384), .A2(new_n388), .A3(KEYINPUT25), .A4(new_n311), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n339), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n384), .A2(new_n388), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n338), .A2(G902), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G214), .B1(G237), .B2(G902), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n201), .A2(KEYINPUT0), .ZN(new_n399));
  INV_X1    g213(.A(new_n250), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G125), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n272), .A2(G224), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT85), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT84), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT86), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n251), .A2(new_n340), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n340), .B2(new_n261), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n404), .B(new_n408), .C1(new_n410), .C2(new_n403), .ZN(new_n411));
  INV_X1    g225(.A(new_n408), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n203), .B(new_n340), .C1(new_n213), .C2(new_n217), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n403), .B1(new_n402), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n409), .A2(KEYINPUT83), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G104), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT3), .B1(new_n418), .B2(G107), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT3), .ZN(new_n420));
  INV_X1    g234(.A(G107), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n421), .A3(G104), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(G107), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G101), .ZN(new_n425));
  INV_X1    g239(.A(G101), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n419), .A2(new_n422), .A3(new_n426), .A4(new_n423), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(KEYINPUT4), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n424), .A2(new_n429), .A3(G101), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n255), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n418), .A2(G107), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n421), .A2(G104), .ZN(new_n433));
  OAI21_X1  g247(.A(G101), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n253), .A2(new_n254), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n361), .A3(G116), .ZN(new_n439));
  OAI211_X1 g253(.A(G113), .B(new_n439), .C1(new_n253), .C2(new_n438), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n431), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT81), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n431), .A2(new_n445), .A3(new_n441), .ZN(new_n446));
  XNOR2_X1  g260(.A(G110), .B(G122), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n443), .A2(new_n444), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT82), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n442), .B2(KEYINPUT81), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT82), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n444), .A4(new_n446), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n446), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n431), .A2(new_n441), .A3(new_n447), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n417), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G210), .B1(G237), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n406), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n404), .B(new_n461), .C1(new_n410), .C2(new_n403), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n440), .A2(new_n437), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n436), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n447), .B(KEYINPUT8), .Z(new_n465));
  OAI21_X1  g279(.A(new_n456), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n461), .B1(new_n402), .B2(new_n413), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(G902), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n458), .A2(new_n459), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n459), .B1(new_n458), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n398), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n473));
  INV_X1    g287(.A(G116), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT90), .B1(new_n474), .B2(G122), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n476));
  INV_X1    g290(.A(G122), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(G116), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n474), .A2(G122), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n421), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(KEYINPUT14), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n479), .B(new_n480), .C1(KEYINPUT14), .C2(new_n421), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n197), .A2(G128), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n190), .A2(G143), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G128), .B(G143), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n485), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n239), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n486), .A2(new_n487), .A3(new_n485), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n493), .A2(new_n488), .A3(new_n244), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n483), .B(new_n484), .C1(new_n492), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(KEYINPUT13), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(G134), .C1(KEYINPUT13), .C2(new_n486), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n244), .B1(new_n493), .B2(new_n488), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n479), .A2(new_n421), .A3(new_n480), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n497), .B(new_n498), .C1(new_n499), .C2(new_n481), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT9), .B(G234), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n502), .A2(G217), .A3(new_n272), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n495), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT92), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n495), .A2(new_n500), .A3(new_n506), .A4(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n495), .A2(new_n500), .ZN(new_n508));
  INV_X1    g322(.A(new_n503), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n311), .ZN(new_n512));
  INV_X1    g326(.A(G478), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n511), .B(new_n311), .C1(KEYINPUT15), .C2(new_n513), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT87), .B(G143), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n271), .A2(new_n272), .A3(G214), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n271), .A2(new_n272), .A3(G214), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT87), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n522), .B1(new_n523), .B2(new_n197), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n521), .A2(new_n219), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n219), .B1(new_n521), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n518), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n521), .A2(new_n524), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT17), .B1(new_n528), .B2(new_n219), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n357), .A2(new_n530), .A3(new_n358), .ZN(new_n531));
  AND2_X1   g345(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G131), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n528), .A2(new_n533), .B1(new_n526), .B2(new_n532), .ZN(new_n534));
  OAI22_X1  g348(.A1(new_n355), .A2(new_n192), .B1(new_n208), .B2(new_n374), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n418), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT89), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n531), .A2(KEYINPUT89), .A3(new_n536), .A4(new_n540), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n311), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G475), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT20), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n525), .A2(new_n526), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n341), .A2(new_n548), .A3(new_n344), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n355), .B2(new_n548), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n357), .B(new_n547), .C1(new_n208), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n539), .B1(new_n534), .B2(new_n535), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n537), .A2(new_n539), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(G475), .A2(G902), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n546), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n553), .A2(new_n546), .A3(new_n554), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n517), .B(new_n545), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(G234), .A2(G237), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(G952), .A3(new_n272), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(G902), .A3(G953), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT21), .B(G898), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n473), .B1(new_n557), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n537), .A2(new_n539), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n551), .A2(new_n552), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n554), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT20), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n553), .A2(new_n546), .A3(new_n554), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n569), .A2(new_n570), .B1(G475), .B2(new_n544), .ZN(new_n571));
  INV_X1    g385(.A(new_n564), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n571), .A2(KEYINPUT93), .A3(new_n517), .A4(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n472), .B1(new_n565), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G140), .ZN(new_n575));
  INV_X1    g389(.A(G227), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(G953), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n575), .B(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n428), .A2(new_n430), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n251), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n436), .A2(KEYINPUT10), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n261), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(G128), .B1(new_n210), .B2(new_n202), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n199), .A2(new_n200), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n203), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n584), .B1(new_n587), .B2(new_n436), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n582), .A2(new_n248), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n248), .ZN(new_n590));
  INV_X1    g404(.A(new_n581), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n218), .A2(new_n591), .B1(new_n579), .B2(new_n251), .ZN(new_n592));
  AOI211_X1 g406(.A(KEYINPUT1), .B(new_n190), .C1(new_n199), .C2(new_n200), .ZN(new_n593));
  INV_X1    g407(.A(new_n586), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n436), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n583), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n590), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n578), .B1(new_n589), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n578), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n592), .A2(new_n590), .A3(new_n596), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n203), .B(new_n435), .C1(new_n213), .C2(new_n217), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n601), .B(new_n590), .C1(new_n602), .C2(new_n595), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n595), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT12), .B1(new_n604), .B2(new_n248), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n599), .B(new_n600), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G469), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n311), .ZN(new_n609));
  INV_X1    g423(.A(new_n597), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n599), .A3(new_n600), .ZN(new_n611));
  INV_X1    g425(.A(new_n603), .ZN(new_n612));
  INV_X1    g426(.A(new_n605), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n589), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n611), .B(G469), .C1(new_n614), .C2(new_n599), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n608), .A2(new_n311), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n609), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n381), .B1(new_n502), .B2(new_n311), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n574), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n335), .A2(new_n397), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  NAND2_X1  g439(.A1(new_n277), .A2(new_n281), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT69), .B1(new_n327), .B2(new_n282), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n329), .A4(new_n320), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n311), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(G472), .ZN(new_n630));
  INV_X1    g444(.A(new_n397), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n621), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n331), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n458), .A2(new_n469), .ZN(new_n635));
  INV_X1    g449(.A(new_n459), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n458), .A2(new_n459), .A3(new_n469), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(KEYINPUT94), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT94), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n458), .A2(new_n469), .A3(new_n640), .A4(new_n459), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n641), .A2(new_n398), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n571), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n311), .A2(G478), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n503), .B1(new_n495), .B2(new_n500), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI221_X4 g462(.A(new_n645), .B1(new_n648), .B2(new_n504), .C1(new_n511), .C2(new_n647), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(KEYINPUT92), .B2(new_n504), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n650), .B2(new_n507), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT95), .B1(new_n651), .B2(G478), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT95), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n512), .A2(new_n653), .A3(new_n513), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n644), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n643), .A2(new_n564), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n634), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G104), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  NAND2_X1  g476(.A1(new_n515), .A2(new_n516), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n663), .B(new_n545), .C1(new_n556), .C2(new_n555), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n643), .A2(new_n564), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n634), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n391), .A2(new_n392), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n373), .A2(new_n379), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n385), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n669), .A2(new_n338), .B1(new_n395), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n621), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n574), .A2(new_n630), .A3(new_n331), .A4(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  AND2_X1   g491(.A1(new_n639), .A2(new_n642), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n272), .A2(G900), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(G902), .A3(new_n558), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n559), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT98), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n664), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n674), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n335), .A2(new_n678), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  NOR2_X1   g502(.A1(new_n571), .A2(new_n517), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n398), .A3(new_n673), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT99), .Z(new_n691));
  NAND2_X1  g505(.A1(new_n637), .A2(new_n638), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT38), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n637), .A2(KEYINPUT38), .A3(new_n638), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n684), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n622), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT40), .ZN(new_n701));
  INV_X1    g515(.A(G472), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n269), .A2(new_n278), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n299), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n704), .B2(new_n311), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n302), .B2(KEYINPUT32), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n303), .A2(new_n706), .A3(new_n334), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n698), .A2(new_n701), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT100), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  INV_X1    g526(.A(new_n684), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n644), .A2(new_n656), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n621), .A3(new_n673), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n335), .A2(new_n678), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT101), .B(G146), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G48));
  INV_X1    g532(.A(new_n607), .ZN(new_n719));
  OAI21_X1  g533(.A(G469), .B1(new_n719), .B2(G902), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n620), .A3(new_n609), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n720), .A2(KEYINPUT102), .A3(new_n620), .A4(new_n609), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n335), .A2(new_n397), .A3(new_n658), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n335), .A2(new_n665), .A3(new_n397), .A4(new_n725), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  AOI211_X1 g544(.A(new_n673), .B(new_n721), .C1(new_n565), .C2(new_n573), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n335), .A2(new_n678), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  NOR2_X1   g547(.A1(new_n289), .A2(new_n294), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n307), .B1(new_n270), .B2(new_n306), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n278), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n188), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  OR3_X1    g552(.A1(new_n393), .A2(KEYINPUT103), .A3(new_n396), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT103), .B1(new_n393), .B2(new_n396), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n630), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n639), .A2(new_n642), .A3(new_n689), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n723), .A2(new_n572), .A3(new_n724), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n477), .ZN(G24));
  AOI21_X1  g561(.A(new_n702), .B1(new_n628), .B2(new_n311), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n748), .A2(new_n673), .A3(new_n714), .A4(new_n737), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n643), .A2(new_n721), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  NAND3_X1  g566(.A1(new_n637), .A2(new_n398), .A3(new_n638), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n621), .A2(new_n714), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n304), .A2(new_n319), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n302), .A2(KEYINPUT32), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n741), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT42), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n621), .A2(new_n753), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n335), .A2(new_n397), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n219), .ZN(G33));
  NAND4_X1  g577(.A1(new_n335), .A2(new_n397), .A3(new_n685), .A4(new_n759), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  OAI21_X1  g579(.A(new_n611), .B1(new_n614), .B2(new_n599), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n608), .B1(new_n766), .B2(new_n767), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n616), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n609), .B1(new_n770), .B2(KEYINPUT46), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n620), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n699), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT104), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n656), .A2(new_n571), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT43), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n656), .A2(new_n779), .A3(new_n571), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT105), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n630), .A2(new_n331), .ZN(new_n783));
  INV_X1    g597(.A(new_n673), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(KEYINPUT44), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n753), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT106), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n776), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(KEYINPUT106), .A3(new_n786), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  XNOR2_X1  g608(.A(new_n773), .B(KEYINPUT47), .ZN(new_n795));
  OR4_X1    g609(.A1(new_n335), .A2(new_n397), .A3(new_n714), .A4(new_n753), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  INV_X1    g612(.A(G952), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n778), .A2(new_n560), .A3(new_n780), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT111), .ZN(new_n801));
  INV_X1    g615(.A(new_n741), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n748), .A3(new_n737), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n799), .B(G953), .C1(new_n804), .C2(new_n750), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n755), .A2(new_n756), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n802), .ZN(new_n807));
  INV_X1    g621(.A(new_n721), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n786), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(new_n801), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g627(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n809), .A2(new_n631), .A3(new_n559), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n708), .A2(new_n644), .A3(new_n656), .A4(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n805), .A2(new_n813), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n708), .A2(new_n571), .A3(new_n655), .A4(new_n816), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n748), .A2(new_n673), .A3(new_n737), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n801), .A2(new_n820), .A3(new_n810), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n697), .A2(new_n398), .A3(new_n721), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n804), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n801), .A2(new_n803), .A3(new_n826), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n824), .A2(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n823), .B1(new_n832), .B2(KEYINPUT114), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT47), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n773), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n773), .A2(new_n834), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n720), .A2(new_n619), .A3(new_n609), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n801), .A2(new_n803), .A3(new_n786), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT112), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n827), .A2(new_n831), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n833), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n827), .A2(new_n831), .A3(new_n821), .A4(new_n819), .ZN(new_n848));
  INV_X1    g662(.A(new_n840), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT51), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n818), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n557), .A2(new_n684), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n674), .A2(new_n786), .A3(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n335), .A2(new_n856), .B1(new_n749), .B2(new_n759), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n664), .B1(new_n571), .B2(new_n655), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n572), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n472), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(new_n630), .A3(new_n331), .A4(new_n632), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(new_n675), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(new_n764), .A3(new_n624), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n762), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT107), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n729), .A2(new_n732), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n803), .A2(new_n572), .A3(new_n725), .A4(new_n743), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n726), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n865), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n723), .A2(new_n397), .A3(new_n724), .ZN(new_n870));
  AOI211_X1 g684(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n628), .C2(new_n187), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n332), .B1(new_n331), .B2(new_n333), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g687(.A1(KEYINPUT32), .A2(new_n302), .B1(new_n318), .B2(G472), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n746), .B1(new_n875), .B2(new_n658), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(KEYINPUT107), .A3(new_n729), .A4(new_n732), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n864), .A2(new_n869), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n687), .A2(new_n751), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT52), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT108), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n673), .A2(new_n713), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n621), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n672), .A2(new_n395), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n884), .A2(new_n393), .A3(new_n684), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(KEYINPUT108), .A3(new_n620), .A4(new_n618), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n743), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n707), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n879), .A2(new_n880), .A3(new_n716), .A4(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n687), .A2(new_n716), .A3(new_n751), .A4(new_n888), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n854), .B1(new_n878), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n890), .B(new_n880), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT109), .B1(new_n866), .B2(new_n868), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT109), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n876), .A2(new_n896), .A3(new_n729), .A4(new_n732), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n687), .A2(new_n751), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n854), .B1(new_n899), .B2(KEYINPUT52), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n894), .A2(new_n898), .A3(new_n864), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n893), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n903), .A2(KEYINPUT110), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(KEYINPUT110), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n869), .A2(new_n877), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n854), .B1(new_n879), .B2(new_n880), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n894), .A3(new_n864), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n893), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n853), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(G952), .A2(G953), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n620), .A2(new_n398), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n720), .A2(new_n609), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n914), .B(new_n777), .C1(KEYINPUT49), .C2(new_n915), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n915), .A2(KEYINPUT49), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n696), .A3(new_n741), .A4(new_n917), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n912), .A2(new_n913), .B1(new_n707), .B2(new_n918), .ZN(G75));
  NAND2_X1  g733(.A1(new_n799), .A2(G953), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT118), .Z(new_n921));
  AOI21_X1  g735(.A(new_n311), .B1(new_n893), .B2(new_n901), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT56), .B1(new_n922), .B2(G210), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n454), .A2(new_n457), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n417), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT55), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n921), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n922), .A2(G210), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(KEYINPUT117), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n928), .B2(KEYINPUT117), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n927), .B1(new_n929), .B2(new_n932), .ZN(G51));
  INV_X1    g747(.A(new_n921), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n922), .A2(new_n768), .A3(new_n769), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n893), .A2(new_n901), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT54), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n903), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n616), .B(KEYINPUT119), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT57), .Z(new_n940));
  AOI21_X1  g754(.A(new_n719), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n935), .B1(new_n941), .B2(KEYINPUT120), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n943));
  INV_X1    g757(.A(new_n940), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n937), .B2(new_n903), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n719), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n934), .B1(new_n942), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  INV_X1    g762(.A(new_n553), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n934), .ZN(G60));
  INV_X1    g766(.A(new_n938), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n511), .A2(new_n647), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n648), .A2(new_n504), .ZN(new_n955));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT59), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n921), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n911), .A2(new_n958), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n954), .A2(new_n955), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G63));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT60), .Z(new_n965));
  NAND3_X1  g779(.A1(new_n936), .A2(new_n672), .A3(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n936), .A2(new_n965), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n394), .B(KEYINPUT121), .Z(new_n968));
  OAI211_X1 g782(.A(new_n921), .B(new_n966), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G66));
  INV_X1    g785(.A(G224), .ZN(new_n972));
  OAI21_X1  g786(.A(G953), .B1(new_n563), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n862), .A2(new_n624), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n906), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n973), .B1(new_n976), .B2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n924), .B1(G898), .B2(new_n272), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT122), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n977), .B(new_n979), .ZN(G69));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n709), .B(KEYINPUT100), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n879), .A2(new_n716), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT62), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n711), .A2(new_n985), .A3(new_n716), .A4(new_n879), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n795), .A2(new_n796), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n335), .A2(new_n397), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI211_X1 g803(.A(new_n753), .B(new_n700), .C1(new_n657), .C2(new_n664), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n984), .A2(new_n986), .A3(new_n793), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n272), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n287), .B(new_n550), .Z(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT123), .Z(new_n995));
  AOI21_X1  g809(.A(new_n981), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n807), .A2(new_n743), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n776), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(new_n983), .ZN(new_n999));
  INV_X1    g813(.A(new_n764), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n987), .A2(new_n762), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n793), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n679), .B1(new_n1002), .B2(new_n272), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n994), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n996), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n679), .B1(new_n576), .B2(G953), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT124), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1009), .B(new_n996), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(G72));
  XNOR2_X1  g827(.A(new_n288), .B(KEYINPUT127), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n992), .A2(new_n975), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  AOI211_X1 g831(.A(new_n278), .B(new_n1014), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1002), .A2(new_n975), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1017), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1014), .A2(new_n278), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n921), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n288), .A2(new_n276), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1017), .B1(new_n1024), .B2(new_n327), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(new_n908), .B2(new_n893), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n1018), .A2(new_n1023), .A3(new_n1026), .ZN(G57));
endmodule


