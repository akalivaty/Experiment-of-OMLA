//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI211_X1 g003(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n189), .C2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(G104), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT77), .B1(new_n196), .B2(KEYINPUT3), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n193), .A2(new_n194), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT77), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n200), .A3(new_n203), .A4(new_n190), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(new_n204), .A3(KEYINPUT4), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n206), .B(G101), .C1(new_n195), .C2(new_n197), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT68), .A2(G119), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(G116), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G119), .ZN(new_n216));
  INV_X1    g030(.A(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT2), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G113), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n214), .A2(new_n221), .A3(KEYINPUT69), .A4(new_n216), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n221), .B1(new_n214), .B2(new_n216), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n209), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  AOI211_X1 g043(.A(KEYINPUT70), .B(new_n227), .C1(new_n224), .C2(new_n225), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n208), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n196), .A2(new_n194), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n204), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n214), .A2(KEYINPUT5), .A3(new_n216), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(G113), .C1(KEYINPUT5), .C2(new_n214), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n226), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(G110), .B(G122), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT6), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n231), .A2(new_n237), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n238), .B(KEYINPUT80), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT6), .ZN(new_n245));
  INV_X1    g059(.A(new_n242), .ZN(new_n246));
  AOI211_X1 g060(.A(new_n245), .B(new_n246), .C1(new_n231), .C2(new_n237), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G143), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT64), .B(G146), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G143), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n249), .A2(G143), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(new_n251), .B2(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n253), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G125), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT81), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT81), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n263), .A3(G125), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT64), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n268), .A3(G143), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n270));
  INV_X1    g084(.A(new_n257), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n269), .A2(new_n270), .A3(G128), .A4(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G128), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n269), .B2(KEYINPUT1), .ZN(new_n274));
  INV_X1    g088(.A(new_n250), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n266), .A2(new_n268), .ZN(new_n276));
  INV_X1    g090(.A(G143), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n265), .B(new_n272), .C1(new_n274), .C2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n262), .A2(new_n264), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G224), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G953), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n282), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n262), .A2(new_n284), .A3(new_n264), .A4(new_n279), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n244), .A2(new_n248), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n238), .B(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n237), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n234), .B1(new_n226), .B2(new_n236), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n279), .A2(KEYINPUT83), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n261), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n279), .A2(KEYINPUT83), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n295));
  OAI22_X1  g109(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n282), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT84), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n282), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(new_n297), .B2(new_n282), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n262), .A2(new_n264), .A3(new_n279), .A4(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n291), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n239), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n188), .B1(new_n286), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n283), .A2(new_n285), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n239), .A2(KEYINPUT6), .B1(new_n241), .B2(new_n242), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(new_n247), .ZN(new_n309));
  AOI21_X1  g123(.A(G902), .B1(new_n302), .B2(new_n239), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(new_n187), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(G234), .A2(G237), .ZN(new_n313));
  INV_X1    g127(.A(G953), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n313), .A2(G952), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(G902), .A3(G953), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n316), .B(KEYINPUT95), .Z(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT21), .B(G898), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G214), .B1(G237), .B2(G902), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n312), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT9), .B(G234), .ZN(new_n323));
  OAI21_X1  g137(.A(G221), .B1(new_n323), .B2(G902), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT76), .Z(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AND4_X1   g140(.A1(new_n270), .A2(new_n269), .A3(G128), .A4(new_n271), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n273), .B1(new_n250), .B2(KEYINPUT1), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(new_n269), .B2(new_n271), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n204), .B(new_n233), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT10), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n272), .B1(new_n274), .B2(new_n278), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n234), .A2(KEYINPUT10), .A3(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n252), .A2(new_n255), .B1(new_n258), .B2(new_n253), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n205), .A2(new_n335), .A3(new_n207), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT11), .ZN(new_n337));
  INV_X1    g151(.A(G134), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(G137), .ZN(new_n339));
  INV_X1    g153(.A(G137), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT11), .A3(G134), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(G137), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G131), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT65), .B(G131), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n345), .A2(new_n339), .A3(new_n341), .A4(new_n342), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n332), .A2(new_n334), .A3(new_n336), .A4(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G110), .B(G140), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n314), .A2(G227), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT79), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n330), .B1(new_n234), .B2(new_n333), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n347), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT12), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(KEYINPUT12), .A3(new_n347), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n274), .A2(new_n278), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n204), .A2(new_n233), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(new_n272), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n358), .B(new_n348), .C1(new_n365), .C2(new_n330), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT12), .B1(new_n356), .B2(new_n347), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT78), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n349), .A2(new_n369), .A3(new_n353), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n355), .A2(new_n362), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n332), .A2(new_n334), .A3(new_n336), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n347), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n349), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n352), .ZN(new_n375));
  AOI211_X1 g189(.A(G469), .B(G902), .C1(new_n371), .C2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n349), .A3(new_n353), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n332), .A2(new_n334), .A3(new_n336), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n359), .A2(new_n361), .B1(new_n378), .B2(new_n348), .ZN(new_n379));
  OAI211_X1 g193(.A(G469), .B(new_n377), .C1(new_n379), .C2(new_n353), .ZN(new_n380));
  INV_X1    g194(.A(G469), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n304), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n326), .B1(new_n376), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT93), .ZN(new_n386));
  INV_X1    g200(.A(new_n345), .ZN(new_n387));
  INV_X1    g201(.A(G237), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n314), .A3(G214), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT85), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT86), .B1(new_n390), .B2(G143), .ZN(new_n391));
  NOR2_X1   g205(.A1(KEYINPUT86), .A2(G143), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n389), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n391), .A2(new_n389), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n389), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n277), .A2(KEYINPUT85), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n392), .B1(new_n399), .B2(KEYINPUT86), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n345), .B(new_n398), .C1(new_n400), .C2(new_n389), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G140), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G125), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n265), .A2(G140), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT74), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(KEYINPUT74), .A3(G125), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n249), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n249), .A3(new_n411), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT17), .B(new_n387), .C1(new_n394), .C2(new_n395), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n402), .A2(new_n413), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(G113), .B(G122), .Z(new_n417));
  XOR2_X1   g231(.A(KEYINPUT90), .B(G104), .Z(new_n418));
  XOR2_X1   g232(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n422));
  INV_X1    g236(.A(G131), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT87), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n394), .B2(new_n395), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n424), .B(new_n398), .C1(new_n400), .C2(new_n389), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n407), .A2(new_n408), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT88), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n407), .A2(new_n430), .A3(new_n408), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(G146), .A3(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n404), .A2(new_n405), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n251), .ZN(new_n434));
  AOI221_X4 g248(.A(KEYINPUT89), .B1(new_n426), .B2(new_n427), .C1(new_n432), .C2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n434), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n426), .A2(new_n427), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n416), .B(new_n421), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT92), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n407), .A2(new_n430), .A3(new_n408), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n430), .B1(new_n407), .B2(new_n408), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n442), .A2(new_n443), .A3(new_n249), .ZN(new_n444));
  INV_X1    g258(.A(new_n434), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n438), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT89), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n437), .A2(new_n436), .A3(new_n438), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n419), .B1(new_n449), .B2(new_n416), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n441), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n416), .B1(new_n435), .B2(new_n439), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n453));
  INV_X1    g267(.A(new_n419), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n304), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n386), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  AND4_X1   g271(.A1(new_n414), .A2(new_n402), .A3(new_n413), .A4(new_n415), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n447), .B2(new_n448), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n440), .B(KEYINPUT92), .C1(new_n459), .C2(new_n419), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n460), .A2(KEYINPUT93), .A3(new_n304), .A4(new_n455), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(G475), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT19), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n433), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n429), .A2(new_n431), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n251), .B(new_n464), .C1(new_n465), .C2(new_n463), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n412), .B1(new_n396), .B2(new_n401), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n447), .A2(new_n448), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n440), .B1(new_n468), .B2(new_n419), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G475), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n304), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT20), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT20), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n469), .A2(new_n474), .A3(new_n471), .A4(new_n304), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT13), .B1(new_n273), .B2(G143), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(new_n338), .ZN(new_n478));
  XNOR2_X1  g292(.A(G128), .B(G143), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G116), .B(G122), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n483), .A2(G107), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(G107), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n215), .A2(KEYINPUT14), .A3(G122), .ZN(new_n487));
  INV_X1    g301(.A(new_n481), .ZN(new_n488));
  OAI211_X1 g302(.A(G107), .B(new_n487), .C1(new_n488), .C2(KEYINPUT14), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n479), .B(new_n338), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n489), .B(new_n490), .C1(new_n483), .C2(G107), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G217), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n323), .A2(new_n493), .A3(G953), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n492), .B(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n304), .ZN(new_n497));
  INV_X1    g311(.A(G478), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(KEYINPUT15), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n497), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n462), .A2(new_n476), .A3(new_n501), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n322), .A2(new_n385), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT25), .ZN(new_n504));
  NOR2_X1   g318(.A1(G119), .A2(G128), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(KEYINPUT68), .A2(G119), .ZN(new_n507));
  NOR2_X1   g321(.A1(KEYINPUT68), .A2(G119), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(KEYINPUT23), .B(new_n506), .C1(new_n509), .C2(new_n273), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n509), .B2(G128), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G110), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n212), .A2(new_n213), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n505), .B1(new_n515), .B2(G128), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT24), .B(G110), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n414), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n514), .B(new_n518), .C1(new_n519), .C2(new_n412), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n412), .A2(new_n445), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n517), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n513), .B2(G110), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT22), .B(G137), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n314), .A2(G221), .A3(G234), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n520), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n520), .B2(new_n524), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n528), .A2(new_n529), .A3(G902), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n504), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n520), .A2(new_n524), .A3(new_n527), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n304), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n493), .B1(G234), .B2(new_n304), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(G902), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(G472), .A2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n226), .A2(new_n228), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT70), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n226), .A2(new_n209), .A3(new_n228), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n343), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT66), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n338), .B2(G137), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n340), .A2(KEYINPUT66), .A3(G134), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n342), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n548), .A2(new_n345), .B1(new_n552), .B2(G131), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n347), .A2(new_n335), .B1(new_n333), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT30), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT67), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n333), .A2(new_n556), .A3(new_n553), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n260), .A2(new_n348), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n333), .B2(new_n553), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n547), .B(new_n555), .C1(new_n560), .C2(KEYINPUT30), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n545), .A2(new_n554), .A3(new_n546), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n388), .A2(new_n314), .A3(G210), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT27), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT26), .B(G101), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n562), .A2(KEYINPUT71), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT71), .B1(new_n562), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n561), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT31), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n561), .B(KEYINPUT31), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OR3_X1    g387(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n333), .A2(new_n553), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n348), .B2(new_n260), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n576), .A2(new_n229), .A3(new_n230), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n574), .A2(new_n547), .B1(new_n577), .B2(KEYINPUT28), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT28), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n562), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n566), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n543), .B1(new_n573), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n576), .B1(new_n230), .B2(new_n229), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n562), .A3(KEYINPUT73), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n547), .A2(new_n586), .A3(new_n576), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(KEYINPUT28), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n588), .A2(KEYINPUT29), .A3(new_n566), .A4(new_n580), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n574), .A2(new_n547), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n577), .A2(KEYINPUT28), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n580), .ZN(new_n593));
  INV_X1    g407(.A(new_n566), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n566), .B1(new_n561), .B2(new_n562), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n589), .B(new_n304), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n583), .A2(KEYINPUT32), .B1(G472), .B2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n599));
  AOI21_X1  g413(.A(new_n581), .B1(new_n571), .B2(new_n572), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n543), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n541), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n503), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n462), .A2(new_n476), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n496), .A2(new_n606), .A3(KEYINPUT33), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n492), .A2(new_n495), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n494), .B1(new_n486), .B2(new_n491), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(G478), .A3(new_n304), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n497), .A2(new_n498), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n605), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT98), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n605), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n309), .A2(new_n310), .A3(new_n187), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n187), .B1(new_n309), .B2(new_n310), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n321), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT96), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n312), .A2(new_n626), .A3(new_n321), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n319), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n573), .A2(new_n582), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n304), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n583), .B1(new_n630), .B2(G472), .ZN(new_n631));
  AOI21_X1  g445(.A(G902), .B1(new_n371), .B2(new_n375), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n384), .B1(new_n632), .B2(new_n381), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n633), .A2(new_n541), .A3(new_n325), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n621), .A2(new_n628), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  AOI21_X1  g452(.A(new_n626), .B1(new_n312), .B2(new_n321), .ZN(new_n639));
  INV_X1    g453(.A(new_n321), .ZN(new_n640));
  AOI211_X1 g454(.A(KEYINPUT96), .B(new_n640), .C1(new_n306), .C2(new_n311), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n320), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n461), .A2(G475), .ZN(new_n644));
  AOI21_X1  g458(.A(G902), .B1(new_n450), .B2(new_n453), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT93), .B1(new_n645), .B2(new_n460), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n457), .A2(KEYINPUT99), .A3(G475), .A4(new_n461), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n647), .A2(new_n648), .B1(new_n473), .B2(new_n475), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n497), .B(new_n499), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n642), .A2(KEYINPUT100), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  INV_X1    g467(.A(new_n651), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n653), .B1(new_n654), .B2(new_n628), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n635), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT101), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT35), .B(G107), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR2_X1   g473(.A1(new_n385), .A2(new_n502), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n319), .B(new_n640), .C1(new_n306), .C2(new_n311), .ZN(new_n661));
  INV_X1    g475(.A(new_n527), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(KEYINPUT36), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n520), .A2(new_n524), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n520), .B2(new_n524), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT102), .B1(new_n666), .B2(new_n539), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n668));
  INV_X1    g482(.A(new_n539), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n664), .A2(new_n665), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n538), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n660), .A2(new_n631), .A3(new_n661), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  AOI21_X1  g489(.A(new_n385), .B1(new_n625), .B2(new_n627), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n647), .A2(new_n648), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n315), .B1(new_n317), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n476), .A2(new_n677), .A3(new_n650), .A4(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n672), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n598), .B2(new_n601), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n676), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  NAND3_X1  g499(.A1(new_n585), .A2(new_n594), .A3(new_n587), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n569), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n304), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n583), .A2(KEYINPUT32), .B1(G472), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n689), .A2(new_n601), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n605), .A2(new_n650), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n690), .A2(new_n640), .A3(new_n672), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n312), .B(KEYINPUT38), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n679), .B(KEYINPUT39), .Z(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n385), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT40), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n692), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NAND2_X1  g513(.A1(new_n625), .A2(new_n627), .ZN(new_n700));
  INV_X1    g514(.A(new_n385), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n605), .A2(new_n616), .A3(new_n680), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n683), .A2(new_n700), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  OR2_X1    g518(.A1(new_n632), .A2(new_n381), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n371), .A2(new_n375), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n381), .A3(new_n304), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n326), .A3(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n621), .A2(new_n628), .A3(new_n602), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND2_X1  g526(.A1(new_n602), .A2(new_n709), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT100), .B1(new_n642), .B2(new_n651), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n654), .A2(new_n628), .A3(new_n653), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n215), .ZN(G18));
  NAND3_X1  g531(.A1(new_n629), .A2(KEYINPUT32), .A3(new_n542), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n597), .A2(G472), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n601), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n502), .A2(new_n319), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n720), .A2(new_n721), .A3(new_n672), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n708), .B1(new_n625), .B2(new_n627), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  INV_X1    g539(.A(new_n541), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n588), .A2(new_n580), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n594), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n543), .B1(new_n573), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(G472), .B1(new_n600), .B2(G902), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT103), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n732), .B(G472), .C1(new_n600), .C2(G902), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n729), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n691), .A2(new_n319), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n723), .A2(new_n726), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NAND4_X1  g551(.A1(new_n723), .A2(new_n672), .A3(new_n702), .A4(new_n734), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  OAI21_X1  g553(.A(new_n598), .B1(KEYINPUT32), .B2(new_n583), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n726), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n617), .A2(new_n743), .A3(new_n679), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n306), .A2(new_n321), .A3(new_n311), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n385), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n702), .A2(new_n746), .A3(new_n720), .A4(new_n726), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT104), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n743), .B1(new_n748), .B2(KEYINPUT104), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  NAND3_X1  g567(.A1(new_n681), .A2(new_n602), .A3(new_n746), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  INV_X1    g569(.A(new_n605), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n616), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(KEYINPUT43), .A3(new_n616), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n758), .B1(new_n757), .B2(new_n759), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT108), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n763), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n761), .A3(new_n766), .A4(new_n760), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n631), .A2(new_n682), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n764), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n764), .A2(new_n767), .A3(KEYINPUT44), .A4(new_n768), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n377), .B1(new_n379), .B2(new_n353), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(G469), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n773), .B(new_n774), .C1(new_n780), .C2(new_n382), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n382), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT105), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n376), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n326), .A3(new_n694), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n745), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n771), .A2(new_n772), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT109), .B(G137), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G39));
  INV_X1    g604(.A(new_n720), .ZN(new_n791));
  INV_X1    g605(.A(new_n745), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n541), .A3(new_n702), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n785), .A2(new_n326), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n785), .A2(KEYINPUT47), .A3(new_n326), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n403), .ZN(G42));
  OAI211_X1 g613(.A(new_n602), .B(new_n709), .C1(new_n652), .C2(new_n655), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n462), .A2(new_n476), .A3(new_n650), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n631), .A2(new_n661), .A3(new_n634), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n673), .A2(new_n803), .A3(KEYINPUT110), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT110), .B1(new_n673), .B2(new_n803), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n617), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n635), .A2(new_n661), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n724), .A2(new_n809), .A3(new_n603), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n710), .A2(new_n736), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n800), .A2(new_n807), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n731), .A2(new_n733), .ZN(new_n814));
  INV_X1    g628(.A(new_n729), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n702), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n720), .A2(new_n649), .A3(new_n501), .A4(new_n680), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n385), .A2(new_n745), .A3(new_n682), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n752), .A2(new_n754), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n813), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  INV_X1    g637(.A(new_n384), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n707), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n679), .B(KEYINPUT111), .Z(new_n826));
  AND3_X1   g640(.A1(new_n538), .A2(new_n671), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n326), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n601), .B2(new_n689), .ZN(new_n829));
  INV_X1    g643(.A(new_n691), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n700), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n738), .A2(new_n684), .A3(new_n703), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT53), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n822), .A2(KEYINPUT53), .A3(new_n834), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT112), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n722), .A2(new_n723), .B1(new_n503), .B2(new_n602), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n710), .A3(new_n736), .A4(new_n809), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n673), .A2(new_n803), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n804), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n839), .A2(new_n843), .A3(new_n716), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n820), .A2(new_n754), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n748), .A2(KEYINPUT104), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n749), .A3(new_n743), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n847), .B2(new_n747), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n738), .A2(new_n684), .A3(new_n703), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n738), .A2(new_n684), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n831), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n834), .A2(new_n844), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(KEYINPUT54), .B(new_n835), .C1(new_n837), .C2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(KEYINPUT53), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n822), .A2(new_n853), .A3(new_n834), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n315), .ZN(new_n863));
  INV_X1    g677(.A(new_n762), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n864), .B2(new_n765), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n734), .A2(new_n726), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n693), .A2(new_n321), .A3(new_n708), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n708), .A2(new_n745), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n726), .A2(new_n690), .A3(new_n315), .A4(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n756), .A3(new_n615), .A4(new_n614), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n315), .B(new_n871), .C1(new_n762), .C2(new_n763), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n734), .A2(new_n672), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n865), .A2(new_n866), .A3(new_n792), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n705), .A2(new_n707), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n796), .B(new_n797), .C1(new_n326), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n876), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT51), .B1(new_n870), .B2(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n874), .A2(new_n741), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT116), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n885), .A3(KEYINPUT48), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n882), .B2(KEYINPUT48), .ZN(new_n888));
  OR4_X1    g702(.A1(new_n887), .A2(new_n874), .A3(KEYINPUT48), .A4(new_n741), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n884), .A2(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n865), .A2(new_n723), .A3(new_n866), .ZN(new_n891));
  INV_X1    g705(.A(G952), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n892), .B(G953), .C1(new_n872), .C2(new_n621), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n881), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n870), .A2(KEYINPUT51), .A3(new_n880), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI22_X1  g714(.A1(new_n862), .A2(new_n900), .B1(G952), .B2(G953), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n878), .B(KEYINPUT49), .Z(new_n902));
  NOR4_X1   g716(.A1(new_n757), .A2(new_n541), .A3(new_n640), .A4(new_n325), .ZN(new_n903));
  INV_X1    g717(.A(new_n693), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .A4(new_n690), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n314), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n858), .A2(new_n859), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n304), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT56), .B1(new_n910), .B2(G210), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n308), .A2(new_n247), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n307), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n913), .B(new_n914), .Z(new_n915));
  OAI21_X1  g729(.A(new_n908), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n915), .ZN(new_n917));
  AOI211_X1 g731(.A(KEYINPUT56), .B(new_n917), .C1(new_n910), .C2(G210), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n918), .ZN(G51));
  XOR2_X1   g733(.A(new_n706), .B(KEYINPUT118), .Z(new_n920));
  NOR2_X1   g734(.A1(new_n909), .A2(new_n856), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n860), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n382), .B(KEYINPUT57), .Z(new_n923));
  OAI21_X1  g737(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n910), .A2(new_n780), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n907), .B1(new_n924), .B2(new_n925), .ZN(G54));
  NAND3_X1  g740(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n907), .B1(new_n927), .B2(new_n470), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .A4(new_n469), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G60));
  XNOR2_X1  g744(.A(new_n613), .B(KEYINPUT119), .ZN(new_n931));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT59), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n931), .B1(new_n862), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n931), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n908), .B1(new_n922), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT60), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n858), .A2(new_n859), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n533), .A2(new_n534), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n907), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n666), .B(KEYINPUT120), .Z(new_n943));
  NAND4_X1  g757(.A1(new_n858), .A2(new_n859), .A3(new_n939), .A4(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(KEYINPUT61), .B(new_n942), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(G66));
  OAI21_X1  g765(.A(G953), .B1(new_n318), .B2(new_n281), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n813), .B(KEYINPUT122), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n912), .B1(G898), .B2(new_n314), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  NAND3_X1  g770(.A1(new_n742), .A2(new_n700), .A3(new_n830), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n754), .B1(new_n957), .B2(new_n786), .ZN(new_n958));
  INV_X1    g772(.A(new_n849), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n798), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n788), .A3(new_n752), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n960), .A2(new_n788), .A3(new_n963), .A4(new_n752), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n314), .A3(new_n964), .ZN(new_n965));
  MUX2_X1   g779(.A(new_n560), .B(new_n576), .S(KEYINPUT30), .Z(new_n966));
  OAI21_X1  g780(.A(new_n464), .B1(new_n465), .B2(new_n463), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT123), .Z(new_n968));
  XOR2_X1   g782(.A(new_n966), .B(new_n968), .Z(new_n969));
  OAI211_X1 g783(.A(new_n965), .B(new_n969), .C1(new_n678), .C2(new_n314), .ZN(new_n970));
  INV_X1    g784(.A(new_n969), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n849), .A2(new_n698), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n602), .A2(new_n746), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n695), .B(new_n974), .C1(new_n617), .C2(new_n801), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n798), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n788), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n971), .B1(new_n980), .B2(G953), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n970), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n969), .A2(KEYINPUT125), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n314), .B1(G227), .B2(G900), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n970), .A2(new_n981), .A3(new_n985), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n980), .B2(new_n953), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n561), .A2(new_n562), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n566), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT126), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n997));
  INV_X1    g811(.A(new_n995), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n844), .B(KEYINPUT122), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n999), .A2(new_n978), .A3(new_n979), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n997), .B(new_n998), .C1(new_n1000), .C2(new_n992), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n962), .A2(new_n953), .A3(new_n964), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n991), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n994), .A2(new_n566), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n907), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n596), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n992), .B1(new_n1007), .B2(new_n569), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n835), .B(new_n1008), .C1(new_n837), .C2(new_n854), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1002), .A2(new_n1006), .A3(new_n1009), .ZN(G57));
endmodule


