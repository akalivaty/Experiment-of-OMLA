//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT85), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT81), .B1(new_n205), .B2(G141gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT81), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(G148gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT82), .B(G148gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n209), .C1(new_n210), .C2(new_n208), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n214), .B2(KEYINPUT2), .ZN(new_n215));
  XOR2_X1   g014(.A(G141gat), .B(G148gat), .Z(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(new_n213), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n211), .A2(new_n215), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G127gat), .ZN(new_n222));
  INV_X1    g021(.A(G134gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT72), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT72), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G134gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n223), .A2(G127gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT73), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230));
  INV_X1    g029(.A(G120gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(G113gat), .ZN(new_n232));
  INV_X1    g031(.A(G113gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(G120gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n230), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT73), .ZN(new_n236));
  INV_X1    g035(.A(new_n228), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT72), .B(G134gat), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n236), .B(new_n237), .C1(new_n238), .C2(new_n222), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n229), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G127gat), .B(G134gat), .ZN(new_n241));
  OR2_X1    g040(.A1(KEYINPUT74), .A2(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(KEYINPUT74), .A2(G120gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n233), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT75), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n231), .B2(G113gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n233), .A2(KEYINPUT75), .A3(G120gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n230), .B(new_n241), .C1(new_n244), .C2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n221), .A2(new_n240), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT4), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT83), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n219), .B1(new_n217), .B2(new_n213), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n206), .A2(new_n209), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(G148gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n205), .A2(KEYINPUT82), .ZN(new_n257));
  OAI21_X1  g056(.A(G141gat), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n253), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G141gat), .B(G148gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n220), .B1(new_n260), .B2(KEYINPUT2), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n252), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n205), .A2(KEYINPUT82), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n255), .A2(G148gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n208), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n206), .A2(new_n209), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n215), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT83), .A3(new_n261), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n263), .A2(KEYINPUT3), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n261), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n240), .A2(KEYINPUT84), .A3(new_n249), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT84), .B1(new_n240), .B2(new_n249), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n270), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n204), .B1(new_n251), .B2(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n263), .B(new_n269), .C1(new_n274), .C2(new_n275), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n278), .A2(new_n204), .A3(new_n250), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT39), .ZN(new_n280));
  OR3_X1    g079(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT92), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT87), .B(KEYINPUT0), .Z(new_n283));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  AOI211_X1 g086(.A(new_n282), .B(new_n287), .C1(new_n277), .C2(new_n280), .ZN(new_n288));
  INV_X1    g087(.A(new_n276), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n250), .B(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n280), .B(new_n203), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n287), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT92), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n281), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT93), .A2(KEYINPUT40), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n296), .B(new_n281), .C1(new_n288), .C2(new_n294), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT80), .B(G64gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(G92gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G8gat), .B(G36gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(G183gat), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT68), .B1(new_n307), .B2(KEYINPUT27), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n306), .B(new_n308), .C1(new_n309), .C2(KEYINPUT68), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(KEYINPUT69), .A3(new_n311), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n309), .A2(KEYINPUT28), .A3(new_n306), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(KEYINPUT26), .ZN(new_n320));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(KEYINPUT26), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(KEYINPUT70), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n318), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n317), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n318), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n307), .A2(new_n306), .ZN(new_n334));
  NAND3_X1  g133(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT65), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n338), .A2(G169gat), .A3(G176gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n321), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n326), .A2(KEYINPUT23), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n333), .A2(new_n334), .A3(new_n343), .A4(new_n335), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n337), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(KEYINPUT66), .A3(new_n346), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT67), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n307), .A2(new_n306), .A3(KEYINPUT67), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n352), .A2(new_n333), .A3(new_n335), .A4(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n342), .A3(KEYINPUT25), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n349), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT79), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n331), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n358), .A2(KEYINPUT29), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n362), .B1(new_n331), .B2(new_n356), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  INV_X1    g163(.A(G211gat), .ZN(new_n365));
  INV_X1    g164(.A(G218gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n364), .B1(KEYINPUT22), .B2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(G211gat), .B(G218gat), .Z(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n360), .A2(new_n363), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n331), .A2(new_n356), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n361), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n370), .B1(new_n374), .B2(new_n359), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n305), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n371), .B1(new_n360), .B2(new_n363), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n370), .A3(new_n359), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n304), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(KEYINPUT30), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n381), .B(new_n305), .C1(new_n372), .C2(new_n375), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  AOI211_X1 g182(.A(new_n383), .B(new_n204), .C1(new_n278), .C2(new_n250), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n251), .A2(new_n204), .A3(new_n276), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n383), .A2(KEYINPUT86), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n386), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n251), .A2(new_n204), .A3(new_n276), .A4(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n384), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n287), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n380), .A2(new_n382), .A3(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n300), .A2(KEYINPUT94), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT94), .B1(new_n300), .B2(new_n392), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT3), .B1(new_n370), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n263), .A2(new_n269), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n399));
  OR3_X1    g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G228gat), .ZN(new_n401));
  INV_X1    g200(.A(G233gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n371), .B1(new_n272), .B2(KEYINPUT29), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n397), .B2(new_n398), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n400), .A2(new_n403), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n397), .B2(new_n221), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n401), .B2(new_n402), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G22gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT90), .B(G22gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT91), .ZN(new_n418));
  INV_X1    g217(.A(new_n416), .ZN(new_n419));
  INV_X1    g218(.A(new_n413), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n412), .B1(new_n406), .B2(new_n408), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT91), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n410), .A2(new_n423), .A3(new_n413), .A4(new_n416), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n418), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n391), .A2(KEYINPUT6), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n387), .A2(new_n389), .ZN(new_n427));
  INV_X1    g226(.A(new_n384), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(KEYINPUT88), .A3(new_n293), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT88), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n390), .B2(new_n287), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n426), .B1(new_n434), .B2(new_n391), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT37), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n377), .A2(new_n378), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n377), .B2(new_n378), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n304), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT38), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT38), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n441), .B(new_n304), .C1(new_n437), .C2(new_n438), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n376), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n425), .B1(new_n435), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT95), .B1(new_n395), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n380), .A2(new_n382), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n425), .B1(new_n435), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT36), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT76), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n240), .A2(new_n249), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n449), .B1(new_n373), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n373), .A2(new_n450), .ZN(new_n452));
  INV_X1    g251(.A(new_n450), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n331), .A2(new_n356), .A3(KEYINPUT76), .A4(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT33), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G43gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n451), .A2(new_n456), .A3(new_n452), .A4(new_n454), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT34), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n465), .A2(KEYINPUT34), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n470), .B(new_n466), .C1(new_n458), .C2(new_n463), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n457), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n469), .B2(new_n471), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n448), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n469), .A2(new_n471), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n473), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(KEYINPUT36), .A3(new_n475), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n447), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n300), .A2(new_n392), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n300), .A2(new_n392), .A3(KEYINPUT94), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n425), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n434), .A2(new_n391), .ZN(new_n489));
  INV_X1    g288(.A(new_n426), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n440), .A2(new_n376), .A3(new_n442), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT95), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n487), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n445), .A2(new_n482), .A3(new_n495), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n476), .A2(new_n477), .A3(new_n488), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n446), .A4(new_n435), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n480), .A2(new_n425), .A3(new_n475), .A4(new_n446), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT35), .B1(new_n500), .B2(new_n491), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(G1gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT16), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(G1gat), .B2(new_n504), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(G8gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(G8gat), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT21), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G183gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G127gat), .B(G155gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT20), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n521), .B(new_n523), .Z(new_n524));
  NOR2_X1   g323(.A1(new_n516), .A2(KEYINPUT21), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G211gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n525), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n524), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT100), .B(G134gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT41), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535));
  INV_X1    g334(.A(G85gat), .ZN(new_n536));
  INV_X1    g335(.A(G92gat), .ZN(new_n537));
  AOI22_X1  g336(.A1(KEYINPUT8), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT7), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(new_n536), .B2(new_n537), .ZN(new_n540));
  NAND3_X1  g339(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G99gat), .B(G106gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT101), .Z(new_n545));
  NOR2_X1   g344(.A1(G29gat), .A2(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G43gat), .B(G50gat), .ZN(new_n549));
  INV_X1    g348(.A(G29gat), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT96), .B(G36gat), .Z(new_n551));
  OAI221_X1 g350(.A(new_n548), .B1(KEYINPUT15), .B2(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n553), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n552), .B(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT17), .B1(new_n559), .B2(KEYINPUT97), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n545), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT102), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n559), .A2(new_n544), .B1(KEYINPUT41), .B2(new_n532), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n534), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n563), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT102), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n533), .ZN(new_n570));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G162gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n566), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n566), .B2(new_n570), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n531), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n566), .A2(new_n570), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n572), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n566), .A2(new_n570), .A3(new_n573), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n530), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n529), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n503), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n511), .B1(new_n557), .B2(new_n560), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n554), .A2(new_n511), .ZN(new_n585));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT18), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n554), .A2(new_n511), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n586), .B(KEYINPUT13), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n584), .A2(KEYINPUT18), .A3(new_n585), .A4(new_n586), .ZN(new_n595));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G197gat), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT11), .B(G169gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT12), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n589), .A2(new_n594), .A3(new_n595), .A4(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n601), .A2(KEYINPUT98), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(KEYINPUT98), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n589), .A2(new_n594), .A3(new_n595), .ZN(new_n604));
  INV_X1    g403(.A(new_n600), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n602), .A2(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n516), .B1(KEYINPUT103), .B2(new_n543), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(new_n544), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n516), .A2(new_n544), .A3(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n614), .B(new_n618), .C1(new_n613), .C2(new_n608), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n613), .B(KEYINPUT104), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n610), .B2(new_n611), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n608), .A2(new_n613), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n617), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n606), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n583), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n435), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT106), .B(G1gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1324gat));
  INV_X1    g431(.A(new_n446), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT108), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n627), .A2(KEYINPUT108), .A3(new_n633), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT16), .B(G8gat), .Z(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n637), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(G8gat), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n627), .A2(KEYINPUT42), .A3(new_n633), .A4(new_n638), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(G1325gat));
  NOR2_X1   g444(.A1(new_n476), .A2(new_n477), .ZN(new_n646));
  AOI21_X1  g445(.A(G15gat), .B1(new_n627), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n478), .A2(new_n481), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(G15gat), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n627), .B2(new_n650), .ZN(G1326gat));
  NAND2_X1  g450(.A1(new_n627), .A2(new_n488), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G22gat), .ZN(new_n653));
  INV_X1    g452(.A(G22gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n627), .A2(new_n654), .A3(new_n488), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  INV_X1    g457(.A(new_n581), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n496), .B2(new_n502), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n626), .A2(new_n529), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(new_n550), .A3(new_n629), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(KEYINPUT110), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(KEYINPUT110), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT45), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n503), .B2(new_n581), .ZN(new_n670));
  AOI211_X1 g469(.A(KEYINPUT44), .B(new_n659), .C1(new_n496), .C2(new_n502), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n661), .ZN(new_n673));
  INV_X1    g472(.A(new_n629), .ZN(new_n674));
  OAI21_X1  g473(.A(G29gat), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n664), .A2(KEYINPUT45), .A3(new_n665), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n668), .A2(new_n675), .A3(new_n676), .ZN(G1328gat));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n551), .A3(new_n633), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT111), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(KEYINPUT111), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n551), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n673), .B2(new_n446), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n679), .A2(KEYINPUT46), .A3(new_n680), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(G1329gat));
  AND2_X1   g486(.A1(new_n662), .A2(new_n646), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(G43gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n649), .A2(G43gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n673), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT47), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n689), .B(new_n693), .C1(new_n673), .C2(new_n690), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(G1330gat));
  OAI211_X1 g494(.A(new_n488), .B(new_n661), .C1(new_n670), .C2(new_n671), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n425), .A2(G50gat), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n696), .A2(G50gat), .B1(new_n662), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT112), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n699), .A2(KEYINPUT112), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1331gat));
  NAND2_X1  g502(.A1(new_n606), .A2(new_n625), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n583), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n629), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g508(.A1(new_n706), .A2(new_n446), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n711));
  AND2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n710), .B2(new_n711), .ZN(G1333gat));
  NAND3_X1  g513(.A1(new_n707), .A2(G71gat), .A3(new_n649), .ZN(new_n715));
  INV_X1    g514(.A(new_n646), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n706), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(G71gat), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g518(.A1(new_n707), .A2(new_n488), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g520(.A1(new_n529), .A2(new_n606), .ZN(new_n722));
  INV_X1    g521(.A(new_n625), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT113), .Z(new_n725));
  AND2_X1   g524(.A1(new_n672), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n726), .A2(G85gat), .A3(new_n629), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n503), .A2(new_n581), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT51), .B1(new_n728), .B2(new_n722), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n660), .A2(new_n730), .A3(new_n606), .A4(new_n529), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(new_n625), .A3(new_n629), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n727), .B1(new_n536), .B2(new_n733), .ZN(G1336gat));
  NAND4_X1  g533(.A1(new_n729), .A2(new_n625), .A3(new_n633), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n537), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n672), .A2(G92gat), .A3(new_n633), .A4(new_n725), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1337gat));
  NAND2_X1  g539(.A1(new_n726), .A2(new_n649), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G99gat), .ZN(new_n742));
  INV_X1    g541(.A(G99gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n732), .A2(new_n743), .A3(new_n625), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n744), .B2(new_n716), .ZN(G1338gat));
  OAI211_X1 g544(.A(new_n488), .B(new_n725), .C1(new_n670), .C2(new_n671), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G106gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n425), .A2(G106gat), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n625), .A3(new_n731), .A4(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(KEYINPUT114), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n747), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(new_n754), .A3(KEYINPUT53), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1339gat));
  AND2_X1   g557(.A1(new_n584), .A2(new_n585), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n759), .A2(new_n586), .B1(new_n591), .B2(new_n593), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n599), .ZN(new_n761));
  INV_X1    g560(.A(new_n603), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n601), .A2(KEYINPUT98), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n625), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n614), .B(KEYINPUT54), .C1(new_n620), .C2(new_n612), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n618), .B1(new_n622), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n765), .A2(KEYINPUT55), .A3(new_n767), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n619), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n764), .B1(new_n606), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n659), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n602), .A2(new_n603), .B1(new_n599), .B2(new_n760), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n770), .A2(new_n619), .A3(new_n771), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n581), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n529), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n604), .A2(new_n605), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n762), .B2(new_n763), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n529), .A2(new_n581), .A3(new_n781), .A4(new_n625), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n674), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n500), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n606), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(new_n233), .ZN(G1340gat));
  OAI21_X1  g587(.A(G120gat), .B1(new_n786), .B2(new_n723), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n242), .A2(new_n243), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n625), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT116), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT117), .ZN(G1341gat));
  NOR2_X1   g593(.A1(new_n786), .A2(new_n529), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(new_n222), .ZN(G1342gat));
  NAND3_X1  g595(.A1(new_n784), .A2(new_n581), .A3(new_n785), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n238), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(KEYINPUT56), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(KEYINPUT56), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n797), .B2(G134gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n797), .A2(new_n801), .A3(G134gat), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n799), .A2(new_n800), .B1(new_n802), .B2(new_n804), .ZN(G1343gat));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806));
  INV_X1    g605(.A(new_n529), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n774), .B2(new_n777), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n806), .B(new_n488), .C1(new_n808), .C2(new_n782), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n649), .A2(new_n674), .A3(new_n633), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n768), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT55), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n768), .A2(new_n811), .A3(new_n769), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n781), .A2(new_n619), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n581), .B1(new_n815), .B2(new_n764), .ZN(new_n816));
  INV_X1    g615(.A(new_n777), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n529), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n425), .B1(new_n818), .B2(new_n783), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n809), .B(new_n810), .C1(new_n819), .C2(new_n806), .ZN(new_n820));
  OAI21_X1  g619(.A(G141gat), .B1(new_n820), .B2(new_n606), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n648), .A2(new_n488), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(KEYINPUT121), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(KEYINPUT121), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n784), .A2(new_n446), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(G141gat), .A3(new_n606), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT122), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n828), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n821), .A4(new_n822), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n783), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n488), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT57), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n809), .A2(new_n810), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n820), .A2(KEYINPUT120), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n781), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n828), .B1(new_n840), .B2(G141gat), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n829), .B(new_n832), .C1(new_n841), .C2(new_n822), .ZN(G1344gat));
  NAND2_X1  g641(.A1(new_n779), .A2(new_n783), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n488), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT57), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n819), .A2(new_n806), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n625), .A3(new_n810), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n849));
  OR3_X1    g648(.A1(new_n827), .A2(new_n723), .A3(new_n210), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n836), .A2(new_n837), .A3(new_n833), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n820), .A2(KEYINPUT120), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n723), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n256), .A3(new_n257), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n849), .B(new_n850), .C1(new_n854), .C2(KEYINPUT59), .ZN(G1345gat));
  INV_X1    g654(.A(new_n827), .ZN(new_n856));
  INV_X1    g655(.A(G155gat), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n857), .A3(new_n807), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n529), .B1(new_n851), .B2(new_n852), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n857), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT123), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n858), .B(new_n862), .C1(new_n859), .C2(new_n857), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1346gat));
  AOI21_X1  g663(.A(G162gat), .B1(new_n856), .B2(new_n581), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n659), .B1(new_n851), .B2(new_n852), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(G162gat), .ZN(G1347gat));
  NAND3_X1  g666(.A1(new_n843), .A2(new_n633), .A3(new_n674), .ZN(new_n868));
  INV_X1    g667(.A(new_n497), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n781), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(G169gat), .ZN(G1348gat));
  NOR2_X1   g672(.A1(new_n870), .A2(new_n723), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(KEYINPUT124), .A3(G176gat), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT124), .B1(new_n874), .B2(G176gat), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(G176gat), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1349gat));
  OR3_X1    g677(.A1(new_n870), .A2(new_n529), .A3(new_n309), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n307), .B1(new_n870), .B2(new_n529), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(G1350gat));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G190gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n659), .ZN(new_n887));
  MUX2_X1   g686(.A(new_n885), .B(new_n886), .S(new_n887), .Z(G1351gat));
  NAND3_X1  g687(.A1(new_n674), .A2(new_n633), .A3(new_n648), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n847), .A2(new_n781), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G197gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n843), .A2(new_n488), .A3(new_n890), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(G197gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n892), .B1(new_n606), .B2(new_n894), .ZN(G1352gat));
  AOI21_X1  g694(.A(new_n893), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n896));
  INV_X1    g695(.A(G204gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n625), .ZN(new_n898));
  NOR2_X1   g697(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n898), .B(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n845), .A2(new_n625), .A3(new_n846), .A4(new_n890), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(G204gat), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(G1353gat));
  INV_X1    g705(.A(new_n893), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n365), .A3(new_n807), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n847), .A2(new_n807), .A3(new_n890), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT63), .B1(new_n909), .B2(G211gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1354gat));
  NAND4_X1  g711(.A1(new_n845), .A2(new_n581), .A3(new_n846), .A4(new_n890), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G218gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n907), .A2(new_n366), .A3(new_n581), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


